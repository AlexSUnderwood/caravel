VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 28.980 2924.800 30.180 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2374.980 2924.800 2376.180 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2609.580 2924.800 2610.780 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2844.180 2924.800 2845.380 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3078.780 2924.800 3079.980 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3313.380 2924.800 3314.580 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 263.580 2924.800 264.780 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3482.700 2.400 3483.900 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3195.060 2.400 3196.260 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2908.100 2.400 2909.300 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2620.460 2.400 2621.660 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2333.500 2.400 2334.700 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2045.860 2.400 2047.060 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 498.180 2924.800 499.380 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1758.900 2.400 1760.100 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 732.780 2924.800 733.980 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 967.380 2924.800 968.580 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1201.980 2924.800 1203.180 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1436.580 2924.800 1437.780 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1671.180 2924.800 1672.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1905.780 2924.800 1906.980 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2140.380 2924.800 2141.580 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2380.110 84.560 2380.430 84.620 ;
        RECT 2414.610 84.560 2414.930 84.620 ;
        RECT 2380.110 84.420 2414.930 84.560 ;
        RECT 2380.110 84.360 2380.430 84.420 ;
        RECT 2414.610 84.360 2414.930 84.420 ;
        RECT 2476.710 84.220 2477.030 84.280 ;
        RECT 2511.210 84.220 2511.530 84.280 ;
        RECT 2476.710 84.080 2511.530 84.220 ;
        RECT 2476.710 84.020 2477.030 84.080 ;
        RECT 2511.210 84.020 2511.530 84.080 ;
        RECT 2705.330 83.880 2705.650 83.940 ;
        RECT 2729.250 83.880 2729.570 83.940 ;
        RECT 2705.330 83.740 2729.570 83.880 ;
        RECT 2705.330 83.680 2705.650 83.740 ;
        RECT 2729.250 83.680 2729.570 83.740 ;
        RECT 2235.210 83.540 2235.530 83.600 ;
        RECT 2246.250 83.540 2246.570 83.600 ;
        RECT 2235.210 83.400 2246.570 83.540 ;
        RECT 2235.210 83.340 2235.530 83.400 ;
        RECT 2246.250 83.340 2246.570 83.400 ;
      LAYER via ;
        RECT 2380.140 84.360 2380.400 84.620 ;
        RECT 2414.640 84.360 2414.900 84.620 ;
        RECT 2476.740 84.020 2477.000 84.280 ;
        RECT 2511.240 84.020 2511.500 84.280 ;
        RECT 2705.360 83.680 2705.620 83.940 ;
        RECT 2729.280 83.680 2729.540 83.940 ;
        RECT 2235.240 83.340 2235.500 83.600 ;
        RECT 2246.280 83.340 2246.540 83.600 ;
      LAYER met2 ;
        RECT 802.330 2380.835 802.610 2381.205 ;
        RECT 802.400 2377.880 802.540 2380.835 ;
        RECT 802.380 2373.880 802.660 2377.880 ;
        RECT 2221.430 85.155 2221.710 85.525 ;
        RECT 2607.830 85.155 2608.110 85.525 ;
        RECT 1849.750 84.050 1850.030 84.165 ;
        RECT 2139.550 84.050 2139.830 84.165 ;
        RECT 1848.900 83.910 1850.030 84.050 ;
        RECT 1848.900 83.485 1849.040 83.910 ;
        RECT 1849.750 83.795 1850.030 83.910 ;
        RECT 2138.700 83.910 2139.830 84.050 ;
        RECT 2138.700 83.485 2138.840 83.910 ;
        RECT 2139.550 83.795 2139.830 83.910 ;
        RECT 2221.500 83.485 2221.640 85.155 ;
        RECT 2318.030 84.475 2318.310 84.845 ;
        RECT 2246.270 83.795 2246.550 84.165 ;
        RECT 2246.340 83.630 2246.480 83.795 ;
        RECT 2235.240 83.485 2235.500 83.630 ;
        RECT 1848.830 83.115 1849.110 83.485 ;
        RECT 2138.630 83.115 2138.910 83.485 ;
        RECT 2221.430 83.115 2221.710 83.485 ;
        RECT 2235.230 83.115 2235.510 83.485 ;
        RECT 2246.280 83.310 2246.540 83.630 ;
        RECT 2318.100 82.125 2318.240 84.475 ;
        RECT 2380.140 84.330 2380.400 84.650 ;
        RECT 2414.630 84.475 2414.910 84.845 ;
        RECT 2511.230 84.475 2511.510 84.845 ;
        RECT 2414.640 84.330 2414.900 84.475 ;
        RECT 2380.200 84.165 2380.340 84.330 ;
        RECT 2511.300 84.310 2511.440 84.475 ;
        RECT 2476.740 84.165 2477.000 84.310 ;
        RECT 2380.130 83.795 2380.410 84.165 ;
        RECT 2476.730 83.795 2477.010 84.165 ;
        RECT 2511.240 83.990 2511.500 84.310 ;
        RECT 2607.900 83.485 2608.040 85.155 ;
        RECT 2655.670 84.730 2655.950 84.845 ;
        RECT 2655.280 84.590 2655.950 84.730 ;
        RECT 2655.280 84.165 2655.420 84.590 ;
        RECT 2655.670 84.475 2655.950 84.590 ;
        RECT 2655.210 83.795 2655.490 84.165 ;
        RECT 2705.350 83.795 2705.630 84.165 ;
        RECT 2705.360 83.650 2705.620 83.795 ;
        RECT 2729.280 83.650 2729.540 83.970 ;
        RECT 2729.340 83.485 2729.480 83.650 ;
        RECT 2607.830 83.115 2608.110 83.485 ;
        RECT 2729.270 83.115 2729.550 83.485 ;
        RECT 2318.030 81.755 2318.310 82.125 ;
      LAYER via2 ;
        RECT 802.330 2380.880 802.610 2381.160 ;
        RECT 2221.430 85.200 2221.710 85.480 ;
        RECT 2607.830 85.200 2608.110 85.480 ;
        RECT 1849.750 83.840 1850.030 84.120 ;
        RECT 2139.550 83.840 2139.830 84.120 ;
        RECT 2318.030 84.520 2318.310 84.800 ;
        RECT 2246.270 83.840 2246.550 84.120 ;
        RECT 1848.830 83.160 1849.110 83.440 ;
        RECT 2138.630 83.160 2138.910 83.440 ;
        RECT 2221.430 83.160 2221.710 83.440 ;
        RECT 2235.230 83.160 2235.510 83.440 ;
        RECT 2414.630 84.520 2414.910 84.800 ;
        RECT 2511.230 84.520 2511.510 84.800 ;
        RECT 2380.130 83.840 2380.410 84.120 ;
        RECT 2476.730 83.840 2477.010 84.120 ;
        RECT 2655.670 84.520 2655.950 84.800 ;
        RECT 2655.210 83.840 2655.490 84.120 ;
        RECT 2705.350 83.840 2705.630 84.120 ;
        RECT 2607.830 83.160 2608.110 83.440 ;
        RECT 2729.270 83.160 2729.550 83.440 ;
        RECT 2318.030 81.800 2318.310 82.080 ;
      LAYER met3 ;
        RECT 802.305 2381.170 802.635 2381.185 ;
        RECT 1783.230 2381.170 1783.610 2381.180 ;
        RECT 802.305 2380.870 1783.610 2381.170 ;
        RECT 802.305 2380.855 802.635 2380.870 ;
        RECT 1783.230 2380.860 1783.610 2380.870 ;
        RECT 2917.600 88.210 2924.800 88.660 ;
        RECT 2916.710 87.910 2924.800 88.210 ;
        RECT 1869.710 86.850 1870.090 86.860 ;
        RECT 1917.550 86.850 1917.930 86.860 ;
        RECT 1869.710 86.550 1917.930 86.850 ;
        RECT 1869.710 86.540 1870.090 86.550 ;
        RECT 1917.550 86.540 1917.930 86.550 ;
        RECT 1918.470 85.180 1918.850 85.500 ;
        RECT 2173.310 85.490 2173.690 85.500 ;
        RECT 2221.405 85.490 2221.735 85.505 ;
        RECT 2173.310 85.190 2221.735 85.490 ;
        RECT 2173.310 85.180 2173.690 85.190 ;
        RECT 1917.550 84.810 1917.930 84.820 ;
        RECT 1918.510 84.810 1918.810 85.180 ;
        RECT 2221.405 85.175 2221.735 85.190 ;
        RECT 2559.710 85.490 2560.090 85.500 ;
        RECT 2607.805 85.490 2608.135 85.505 ;
        RECT 2559.710 85.190 2608.135 85.490 ;
        RECT 2559.710 85.180 2560.090 85.190 ;
        RECT 2607.805 85.175 2608.135 85.190 ;
        RECT 1917.550 84.510 1918.810 84.810 ;
        RECT 1919.390 84.810 1919.770 84.820 ;
        RECT 2318.005 84.810 2318.335 84.825 ;
        RECT 2414.605 84.810 2414.935 84.825 ;
        RECT 2511.205 84.810 2511.535 84.825 ;
        RECT 2655.645 84.810 2655.975 84.825 ;
        RECT 2752.910 84.810 2753.290 84.820 ;
        RECT 1919.390 84.510 1994.250 84.810 ;
        RECT 1917.550 84.500 1917.930 84.510 ;
        RECT 1919.390 84.500 1919.770 84.510 ;
        RECT 1849.725 84.130 1850.055 84.145 ;
        RECT 1869.710 84.130 1870.090 84.140 ;
        RECT 1849.725 83.830 1870.090 84.130 ;
        RECT 1993.950 84.130 1994.250 84.510 ;
        RECT 2042.710 84.510 2090.850 84.810 ;
        RECT 1993.950 83.830 2042.090 84.130 ;
        RECT 1849.725 83.815 1850.055 83.830 ;
        RECT 1869.710 83.820 1870.090 83.830 ;
        RECT 1783.230 83.450 1783.610 83.460 ;
        RECT 1848.805 83.450 1849.135 83.465 ;
        RECT 1783.230 83.150 1849.135 83.450 ;
        RECT 2041.790 83.450 2042.090 83.830 ;
        RECT 2042.710 83.450 2043.010 84.510 ;
        RECT 2041.790 83.150 2043.010 83.450 ;
        RECT 2090.550 83.450 2090.850 84.510 ;
        RECT 2318.005 84.510 2332.810 84.810 ;
        RECT 2318.005 84.495 2318.335 84.510 ;
        RECT 2139.525 84.130 2139.855 84.145 ;
        RECT 2173.310 84.130 2173.690 84.140 ;
        RECT 2139.525 83.830 2173.690 84.130 ;
        RECT 2139.525 83.815 2139.855 83.830 ;
        RECT 2173.310 83.820 2173.690 83.830 ;
        RECT 2246.245 84.130 2246.575 84.145 ;
        RECT 2269.910 84.130 2270.290 84.140 ;
        RECT 2246.245 83.830 2270.290 84.130 ;
        RECT 2332.510 84.130 2332.810 84.510 ;
        RECT 2414.605 84.510 2429.410 84.810 ;
        RECT 2414.605 84.495 2414.935 84.510 ;
        RECT 2380.105 84.130 2380.435 84.145 ;
        RECT 2332.510 83.830 2380.435 84.130 ;
        RECT 2429.110 84.130 2429.410 84.510 ;
        RECT 2511.205 84.510 2526.010 84.810 ;
        RECT 2511.205 84.495 2511.535 84.510 ;
        RECT 2476.705 84.130 2477.035 84.145 ;
        RECT 2429.110 83.830 2477.035 84.130 ;
        RECT 2525.710 84.130 2526.010 84.510 ;
        RECT 2655.645 84.510 2669.530 84.810 ;
        RECT 2655.645 84.495 2655.975 84.510 ;
        RECT 2559.710 84.130 2560.090 84.140 ;
        RECT 2525.710 83.830 2560.090 84.130 ;
        RECT 2246.245 83.815 2246.575 83.830 ;
        RECT 2269.910 83.820 2270.290 83.830 ;
        RECT 2380.105 83.815 2380.435 83.830 ;
        RECT 2476.705 83.815 2477.035 83.830 ;
        RECT 2559.710 83.820 2560.090 83.830 ;
        RECT 2608.470 84.130 2608.850 84.140 ;
        RECT 2655.185 84.130 2655.515 84.145 ;
        RECT 2608.470 83.830 2655.515 84.130 ;
        RECT 2608.470 83.820 2608.850 83.830 ;
        RECT 2655.185 83.815 2655.515 83.830 ;
        RECT 2669.230 83.960 2669.530 84.510 ;
        RECT 2752.910 84.510 2836.050 84.810 ;
        RECT 2752.910 84.500 2753.290 84.510 ;
        RECT 2705.325 84.130 2705.655 84.145 ;
        RECT 2671.070 83.960 2705.655 84.130 ;
        RECT 2669.230 83.830 2705.655 83.960 ;
        RECT 2835.750 84.130 2836.050 84.510 ;
        RECT 2916.710 84.130 2917.010 87.910 ;
        RECT 2917.600 87.460 2924.800 87.910 ;
        RECT 2835.750 83.830 2883.890 84.130 ;
        RECT 2669.230 83.660 2671.370 83.830 ;
        RECT 2705.325 83.815 2705.655 83.830 ;
        RECT 2138.605 83.450 2138.935 83.465 ;
        RECT 2090.550 83.150 2138.935 83.450 ;
        RECT 1783.230 83.140 1783.610 83.150 ;
        RECT 1848.805 83.135 1849.135 83.150 ;
        RECT 2138.605 83.135 2138.935 83.150 ;
        RECT 2221.405 83.450 2221.735 83.465 ;
        RECT 2235.205 83.450 2235.535 83.465 ;
        RECT 2221.405 83.150 2235.535 83.450 ;
        RECT 2221.405 83.135 2221.735 83.150 ;
        RECT 2235.205 83.135 2235.535 83.150 ;
        RECT 2607.805 83.450 2608.135 83.465 ;
        RECT 2608.470 83.450 2608.850 83.460 ;
        RECT 2607.805 83.150 2608.850 83.450 ;
        RECT 2607.805 83.135 2608.135 83.150 ;
        RECT 2608.470 83.140 2608.850 83.150 ;
        RECT 2729.245 83.450 2729.575 83.465 ;
        RECT 2752.910 83.450 2753.290 83.460 ;
        RECT 2729.245 83.150 2753.290 83.450 ;
        RECT 2883.590 83.450 2883.890 83.830 ;
        RECT 2884.510 83.830 2917.010 84.130 ;
        RECT 2884.510 83.450 2884.810 83.830 ;
        RECT 2883.590 83.150 2884.810 83.450 ;
        RECT 2729.245 83.135 2729.575 83.150 ;
        RECT 2752.910 83.140 2753.290 83.150 ;
        RECT 2269.910 82.090 2270.290 82.100 ;
        RECT 2318.005 82.090 2318.335 82.105 ;
        RECT 2269.910 81.790 2318.335 82.090 ;
        RECT 2269.910 81.780 2270.290 81.790 ;
        RECT 2318.005 81.775 2318.335 81.790 ;
      LAYER via3 ;
        RECT 1783.260 2380.860 1783.580 2381.180 ;
        RECT 1869.740 86.540 1870.060 86.860 ;
        RECT 1917.580 86.540 1917.900 86.860 ;
        RECT 1918.500 85.180 1918.820 85.500 ;
        RECT 2173.340 85.180 2173.660 85.500 ;
        RECT 1917.580 84.500 1917.900 84.820 ;
        RECT 2559.740 85.180 2560.060 85.500 ;
        RECT 1919.420 84.500 1919.740 84.820 ;
        RECT 1869.740 83.820 1870.060 84.140 ;
        RECT 1783.260 83.140 1783.580 83.460 ;
        RECT 2173.340 83.820 2173.660 84.140 ;
        RECT 2269.940 83.820 2270.260 84.140 ;
        RECT 2559.740 83.820 2560.060 84.140 ;
        RECT 2608.500 83.820 2608.820 84.140 ;
        RECT 2752.940 84.500 2753.260 84.820 ;
        RECT 2608.500 83.140 2608.820 83.460 ;
        RECT 2752.940 83.140 2753.260 83.460 ;
        RECT 2269.940 81.780 2270.260 82.100 ;
      LAYER met4 ;
        RECT 1783.255 2380.855 1783.585 2381.185 ;
        RECT 1783.270 83.465 1783.570 2380.855 ;
        RECT 1869.735 86.535 1870.065 86.865 ;
        RECT 1917.575 86.535 1917.905 86.865 ;
        RECT 1918.510 86.550 1919.730 86.850 ;
        RECT 1869.750 84.145 1870.050 86.535 ;
        RECT 1917.590 84.825 1917.890 86.535 ;
        RECT 1918.510 85.505 1918.810 86.550 ;
        RECT 1918.495 85.175 1918.825 85.505 ;
        RECT 1919.430 84.825 1919.730 86.550 ;
        RECT 2173.335 85.175 2173.665 85.505 ;
        RECT 2559.735 85.175 2560.065 85.505 ;
        RECT 1917.575 84.495 1917.905 84.825 ;
        RECT 1919.415 84.495 1919.745 84.825 ;
        RECT 2173.350 84.145 2173.650 85.175 ;
        RECT 2559.750 84.145 2560.050 85.175 ;
        RECT 2752.935 84.495 2753.265 84.825 ;
        RECT 1869.735 83.815 1870.065 84.145 ;
        RECT 2173.335 83.815 2173.665 84.145 ;
        RECT 2269.935 83.815 2270.265 84.145 ;
        RECT 2559.735 83.815 2560.065 84.145 ;
        RECT 2608.495 83.815 2608.825 84.145 ;
        RECT 1783.255 83.135 1783.585 83.465 ;
        RECT 2269.950 82.105 2270.250 83.815 ;
        RECT 2608.510 83.465 2608.810 83.815 ;
        RECT 2752.950 83.465 2753.250 84.495 ;
        RECT 2608.495 83.135 2608.825 83.465 ;
        RECT 2752.935 83.135 2753.265 83.465 ;
        RECT 2269.935 81.775 2270.265 82.105 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1778.430 2429.200 1778.750 2429.260 ;
        RECT 2900.830 2429.200 2901.150 2429.260 ;
        RECT 1778.430 2429.060 2901.150 2429.200 ;
        RECT 1778.430 2429.000 1778.750 2429.060 ;
        RECT 2900.830 2429.000 2901.150 2429.060 ;
        RECT 1767.390 1715.540 1767.710 1715.600 ;
        RECT 1778.430 1715.540 1778.750 1715.600 ;
        RECT 1767.390 1715.400 1778.750 1715.540 ;
        RECT 1767.390 1715.340 1767.710 1715.400 ;
        RECT 1778.430 1715.340 1778.750 1715.400 ;
      LAYER via ;
        RECT 1778.460 2429.000 1778.720 2429.260 ;
        RECT 2900.860 2429.000 2901.120 2429.260 ;
        RECT 1767.420 1715.340 1767.680 1715.600 ;
        RECT 1778.460 1715.340 1778.720 1715.600 ;
      LAYER met2 ;
        RECT 2900.850 2433.875 2901.130 2434.245 ;
        RECT 2900.920 2429.290 2901.060 2433.875 ;
        RECT 1778.460 2428.970 1778.720 2429.290 ;
        RECT 2900.860 2428.970 2901.120 2429.290 ;
        RECT 1778.520 1715.630 1778.660 2428.970 ;
        RECT 1767.420 1715.485 1767.680 1715.630 ;
        RECT 1767.410 1715.115 1767.690 1715.485 ;
        RECT 1778.460 1715.310 1778.720 1715.630 ;
      LAYER via2 ;
        RECT 2900.850 2433.920 2901.130 2434.200 ;
        RECT 1767.410 1715.160 1767.690 1715.440 ;
      LAYER met3 ;
        RECT 2900.825 2434.210 2901.155 2434.225 ;
        RECT 2917.600 2434.210 2924.800 2434.660 ;
        RECT 2900.825 2433.910 2924.800 2434.210 ;
        RECT 2900.825 2433.895 2901.155 2433.910 ;
        RECT 2917.600 2433.460 2924.800 2433.910 ;
        RECT 1755.835 1715.450 1759.835 1715.455 ;
        RECT 1767.385 1715.450 1767.715 1715.465 ;
        RECT 1755.835 1715.150 1767.715 1715.450 ;
        RECT 1755.835 1714.855 1759.835 1715.150 ;
        RECT 1767.385 1715.135 1767.715 1715.150 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1517.610 2663.800 1517.930 2663.860 ;
        RECT 2900.830 2663.800 2901.150 2663.860 ;
        RECT 1517.610 2663.660 2901.150 2663.800 ;
        RECT 1517.610 2663.600 1517.930 2663.660 ;
        RECT 2900.830 2663.600 2901.150 2663.660 ;
        RECT 1513.470 2388.060 1513.790 2388.120 ;
        RECT 1517.610 2388.060 1517.930 2388.120 ;
        RECT 1513.470 2387.920 1517.930 2388.060 ;
        RECT 1513.470 2387.860 1513.790 2387.920 ;
        RECT 1517.610 2387.860 1517.930 2387.920 ;
      LAYER via ;
        RECT 1517.640 2663.600 1517.900 2663.860 ;
        RECT 2900.860 2663.600 2901.120 2663.860 ;
        RECT 1513.500 2387.860 1513.760 2388.120 ;
        RECT 1517.640 2387.860 1517.900 2388.120 ;
      LAYER met2 ;
        RECT 2900.850 2669.155 2901.130 2669.525 ;
        RECT 2900.920 2663.890 2901.060 2669.155 ;
        RECT 1517.640 2663.570 1517.900 2663.890 ;
        RECT 2900.860 2663.570 2901.120 2663.890 ;
        RECT 1517.700 2388.150 1517.840 2663.570 ;
        RECT 1513.500 2387.830 1513.760 2388.150 ;
        RECT 1517.640 2387.830 1517.900 2388.150 ;
        RECT 1513.560 2377.880 1513.700 2387.830 ;
        RECT 1513.540 2373.880 1513.820 2377.880 ;
      LAYER via2 ;
        RECT 2900.850 2669.200 2901.130 2669.480 ;
      LAYER met3 ;
        RECT 2900.825 2669.490 2901.155 2669.505 ;
        RECT 2917.600 2669.490 2924.800 2669.940 ;
        RECT 2900.825 2669.190 2924.800 2669.490 ;
        RECT 2900.825 2669.175 2901.155 2669.190 ;
        RECT 2917.600 2668.740 2924.800 2669.190 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1777.050 2898.400 1777.370 2898.460 ;
        RECT 2900.830 2898.400 2901.150 2898.460 ;
        RECT 1777.050 2898.260 2901.150 2898.400 ;
        RECT 1777.050 2898.200 1777.370 2898.260 ;
        RECT 2900.830 2898.200 2901.150 2898.260 ;
        RECT 1487.710 1322.840 1488.030 1322.900 ;
        RECT 1777.050 1322.840 1777.370 1322.900 ;
        RECT 1487.710 1322.700 1777.370 1322.840 ;
        RECT 1487.710 1322.640 1488.030 1322.700 ;
        RECT 1777.050 1322.640 1777.370 1322.700 ;
      LAYER via ;
        RECT 1777.080 2898.200 1777.340 2898.460 ;
        RECT 2900.860 2898.200 2901.120 2898.460 ;
        RECT 1487.740 1322.640 1488.000 1322.900 ;
        RECT 1777.080 1322.640 1777.340 1322.900 ;
      LAYER met2 ;
        RECT 2900.850 2903.755 2901.130 2904.125 ;
        RECT 2900.920 2898.490 2901.060 2903.755 ;
        RECT 1777.080 2898.170 1777.340 2898.490 ;
        RECT 2900.860 2898.170 2901.120 2898.490 ;
        RECT 1487.780 1323.135 1488.060 1327.135 ;
        RECT 1487.800 1322.930 1487.940 1323.135 ;
        RECT 1777.140 1322.930 1777.280 2898.170 ;
        RECT 1487.740 1322.610 1488.000 1322.930 ;
        RECT 1777.080 1322.610 1777.340 1322.930 ;
      LAYER via2 ;
        RECT 2900.850 2903.800 2901.130 2904.080 ;
      LAYER met3 ;
        RECT 2900.825 2904.090 2901.155 2904.105 ;
        RECT 2917.600 2904.090 2924.800 2904.540 ;
        RECT 2900.825 2903.790 2924.800 2904.090 ;
        RECT 2900.825 2903.775 2901.155 2903.790 ;
        RECT 2917.600 2903.340 2924.800 2903.790 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 708.930 3133.000 709.250 3133.060 ;
        RECT 2900.830 3133.000 2901.150 3133.060 ;
        RECT 708.930 3132.860 2901.150 3133.000 ;
        RECT 708.930 3132.800 709.250 3132.860 ;
        RECT 2900.830 3132.800 2901.150 3132.860 ;
      LAYER via ;
        RECT 708.960 3132.800 709.220 3133.060 ;
        RECT 2900.860 3132.800 2901.120 3133.060 ;
      LAYER met2 ;
        RECT 2900.850 3138.355 2901.130 3138.725 ;
        RECT 2900.920 3133.090 2901.060 3138.355 ;
        RECT 708.960 3132.770 709.220 3133.090 ;
        RECT 2900.860 3132.770 2901.120 3133.090 ;
        RECT 709.020 1908.605 709.160 3132.770 ;
        RECT 708.950 1908.235 709.230 1908.605 ;
      LAYER via2 ;
        RECT 2900.850 3138.400 2901.130 3138.680 ;
        RECT 708.950 1908.280 709.230 1908.560 ;
      LAYER met3 ;
        RECT 2900.825 3138.690 2901.155 3138.705 ;
        RECT 2917.600 3138.690 2924.800 3139.140 ;
        RECT 2900.825 3138.390 2924.800 3138.690 ;
        RECT 2900.825 3138.375 2901.155 3138.390 ;
        RECT 2917.600 3137.940 2924.800 3138.390 ;
        RECT 708.925 1908.570 709.255 1908.585 ;
        RECT 715.810 1908.570 719.810 1908.575 ;
        RECT 708.925 1908.270 719.810 1908.570 ;
        RECT 708.925 1908.255 709.255 1908.270 ;
        RECT 715.810 1907.975 719.810 1908.270 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2415.070 3368.960 2415.390 3369.020 ;
        RECT 2429.330 3368.960 2429.650 3369.020 ;
        RECT 2415.070 3368.820 2429.650 3368.960 ;
        RECT 2415.070 3368.760 2415.390 3368.820 ;
        RECT 2429.330 3368.760 2429.650 3368.820 ;
      LAYER via ;
        RECT 2415.100 3368.760 2415.360 3369.020 ;
        RECT 2429.360 3368.760 2429.620 3369.020 ;
      LAYER met2 ;
        RECT 2415.090 3368.875 2415.370 3369.245 ;
        RECT 2415.100 3368.730 2415.360 3368.875 ;
        RECT 2429.360 3368.730 2429.620 3369.050 ;
        RECT 1800.530 3368.195 1800.810 3368.565 ;
        RECT 1800.600 3367.770 1800.740 3368.195 ;
        RECT 2429.420 3367.885 2429.560 3368.730 ;
        RECT 1800.990 3367.770 1801.270 3367.885 ;
        RECT 1800.600 3367.630 1801.270 3367.770 ;
        RECT 1800.990 3367.515 1801.270 3367.630 ;
        RECT 2429.350 3367.515 2429.630 3367.885 ;
      LAYER via2 ;
        RECT 2415.090 3368.920 2415.370 3369.200 ;
        RECT 1800.530 3368.240 1800.810 3368.520 ;
        RECT 1800.990 3367.560 1801.270 3367.840 ;
        RECT 2429.350 3367.560 2429.630 3367.840 ;
      LAYER met3 ;
        RECT 2917.600 3373.290 2924.800 3373.740 ;
        RECT 2916.710 3372.990 2924.800 3373.290 ;
        RECT 695.790 3369.210 696.170 3369.220 ;
        RECT 2415.065 3369.210 2415.395 3369.225 ;
        RECT 695.790 3368.910 710.850 3369.210 ;
        RECT 695.790 3368.900 696.170 3368.910 ;
        RECT 710.550 3368.530 710.850 3368.910 ;
        RECT 759.310 3368.910 807.450 3369.210 ;
        RECT 710.550 3368.230 758.690 3368.530 ;
        RECT 758.390 3367.850 758.690 3368.230 ;
        RECT 759.310 3367.850 759.610 3368.910 ;
        RECT 807.150 3368.530 807.450 3368.910 ;
        RECT 855.910 3368.910 904.050 3369.210 ;
        RECT 807.150 3368.230 855.290 3368.530 ;
        RECT 758.390 3367.550 759.610 3367.850 ;
        RECT 854.990 3367.850 855.290 3368.230 ;
        RECT 855.910 3367.850 856.210 3368.910 ;
        RECT 903.750 3368.530 904.050 3368.910 ;
        RECT 952.510 3368.910 1000.650 3369.210 ;
        RECT 903.750 3368.230 951.890 3368.530 ;
        RECT 854.990 3367.550 856.210 3367.850 ;
        RECT 951.590 3367.850 951.890 3368.230 ;
        RECT 952.510 3367.850 952.810 3368.910 ;
        RECT 1000.350 3368.530 1000.650 3368.910 ;
        RECT 1049.110 3368.910 1097.250 3369.210 ;
        RECT 1000.350 3368.230 1048.490 3368.530 ;
        RECT 951.590 3367.550 952.810 3367.850 ;
        RECT 1048.190 3367.850 1048.490 3368.230 ;
        RECT 1049.110 3367.850 1049.410 3368.910 ;
        RECT 1096.950 3368.530 1097.250 3368.910 ;
        RECT 1145.710 3368.910 1193.850 3369.210 ;
        RECT 1096.950 3368.230 1145.090 3368.530 ;
        RECT 1048.190 3367.550 1049.410 3367.850 ;
        RECT 1144.790 3367.850 1145.090 3368.230 ;
        RECT 1145.710 3367.850 1146.010 3368.910 ;
        RECT 1193.550 3368.530 1193.850 3368.910 ;
        RECT 1242.310 3368.910 1290.450 3369.210 ;
        RECT 1193.550 3368.230 1241.690 3368.530 ;
        RECT 1144.790 3367.550 1146.010 3367.850 ;
        RECT 1241.390 3367.850 1241.690 3368.230 ;
        RECT 1242.310 3367.850 1242.610 3368.910 ;
        RECT 1290.150 3368.530 1290.450 3368.910 ;
        RECT 1338.910 3368.910 1387.050 3369.210 ;
        RECT 1290.150 3368.230 1338.290 3368.530 ;
        RECT 1241.390 3367.550 1242.610 3367.850 ;
        RECT 1337.990 3367.850 1338.290 3368.230 ;
        RECT 1338.910 3367.850 1339.210 3368.910 ;
        RECT 1386.750 3368.530 1387.050 3368.910 ;
        RECT 1435.510 3368.910 1483.650 3369.210 ;
        RECT 1386.750 3368.230 1434.890 3368.530 ;
        RECT 1337.990 3367.550 1339.210 3367.850 ;
        RECT 1434.590 3367.850 1434.890 3368.230 ;
        RECT 1435.510 3367.850 1435.810 3368.910 ;
        RECT 1483.350 3368.530 1483.650 3368.910 ;
        RECT 1532.110 3368.910 1580.250 3369.210 ;
        RECT 1483.350 3368.230 1531.490 3368.530 ;
        RECT 1434.590 3367.550 1435.810 3367.850 ;
        RECT 1531.190 3367.850 1531.490 3368.230 ;
        RECT 1532.110 3367.850 1532.410 3368.910 ;
        RECT 1579.950 3368.530 1580.250 3368.910 ;
        RECT 1628.710 3368.910 1676.850 3369.210 ;
        RECT 1579.950 3368.230 1628.090 3368.530 ;
        RECT 1531.190 3367.550 1532.410 3367.850 ;
        RECT 1627.790 3367.850 1628.090 3368.230 ;
        RECT 1628.710 3367.850 1629.010 3368.910 ;
        RECT 1676.550 3368.530 1676.850 3368.910 ;
        RECT 1725.310 3368.910 1787.250 3369.210 ;
        RECT 1676.550 3368.230 1724.690 3368.530 ;
        RECT 1627.790 3367.550 1629.010 3367.850 ;
        RECT 1724.390 3367.850 1724.690 3368.230 ;
        RECT 1725.310 3367.850 1725.610 3368.910 ;
        RECT 1786.950 3368.530 1787.250 3368.910 ;
        RECT 1869.750 3368.910 1917.890 3369.210 ;
        RECT 1800.505 3368.530 1800.835 3368.545 ;
        RECT 1786.950 3368.230 1800.835 3368.530 ;
        RECT 1800.505 3368.215 1800.835 3368.230 ;
        RECT 1724.390 3367.550 1725.610 3367.850 ;
        RECT 1800.965 3367.850 1801.295 3367.865 ;
        RECT 1869.750 3367.850 1870.050 3368.910 ;
        RECT 1800.965 3367.550 1870.050 3367.850 ;
        RECT 1917.590 3367.850 1917.890 3368.910 ;
        RECT 1918.510 3368.910 1966.650 3369.210 ;
        RECT 1918.510 3367.850 1918.810 3368.910 ;
        RECT 1966.350 3368.530 1966.650 3368.910 ;
        RECT 2015.110 3368.910 2063.250 3369.210 ;
        RECT 1966.350 3368.230 2014.490 3368.530 ;
        RECT 1917.590 3367.550 1918.810 3367.850 ;
        RECT 2014.190 3367.850 2014.490 3368.230 ;
        RECT 2015.110 3367.850 2015.410 3368.910 ;
        RECT 2062.950 3368.530 2063.250 3368.910 ;
        RECT 2111.710 3368.910 2159.850 3369.210 ;
        RECT 2062.950 3368.230 2111.090 3368.530 ;
        RECT 2014.190 3367.550 2015.410 3367.850 ;
        RECT 2110.790 3367.850 2111.090 3368.230 ;
        RECT 2111.710 3367.850 2112.010 3368.910 ;
        RECT 2159.550 3368.530 2159.850 3368.910 ;
        RECT 2208.310 3368.910 2256.450 3369.210 ;
        RECT 2159.550 3368.230 2207.690 3368.530 ;
        RECT 2110.790 3367.550 2112.010 3367.850 ;
        RECT 2207.390 3367.850 2207.690 3368.230 ;
        RECT 2208.310 3367.850 2208.610 3368.910 ;
        RECT 2256.150 3368.530 2256.450 3368.910 ;
        RECT 2304.910 3368.910 2353.050 3369.210 ;
        RECT 2256.150 3368.230 2304.290 3368.530 ;
        RECT 2207.390 3367.550 2208.610 3367.850 ;
        RECT 2303.990 3367.850 2304.290 3368.230 ;
        RECT 2304.910 3367.850 2305.210 3368.910 ;
        RECT 2352.750 3368.530 2353.050 3368.910 ;
        RECT 2401.510 3368.910 2415.395 3369.210 ;
        RECT 2352.750 3368.230 2400.890 3368.530 ;
        RECT 2303.990 3367.550 2305.210 3367.850 ;
        RECT 2400.590 3367.850 2400.890 3368.230 ;
        RECT 2401.510 3367.850 2401.810 3368.910 ;
        RECT 2415.065 3368.895 2415.395 3368.910 ;
        RECT 2463.110 3369.210 2463.490 3369.220 ;
        RECT 2463.110 3368.910 2546.250 3369.210 ;
        RECT 2463.110 3368.900 2463.490 3368.910 ;
        RECT 2545.950 3368.530 2546.250 3368.910 ;
        RECT 2594.710 3368.910 2642.850 3369.210 ;
        RECT 2545.950 3368.230 2594.090 3368.530 ;
        RECT 2400.590 3367.550 2401.810 3367.850 ;
        RECT 2429.325 3367.850 2429.655 3367.865 ;
        RECT 2463.110 3367.850 2463.490 3367.860 ;
        RECT 2429.325 3367.550 2463.490 3367.850 ;
        RECT 2593.790 3367.850 2594.090 3368.230 ;
        RECT 2594.710 3367.850 2595.010 3368.910 ;
        RECT 2642.550 3368.530 2642.850 3368.910 ;
        RECT 2691.310 3368.910 2739.450 3369.210 ;
        RECT 2642.550 3368.230 2690.690 3368.530 ;
        RECT 2593.790 3367.550 2595.010 3367.850 ;
        RECT 2690.390 3367.850 2690.690 3368.230 ;
        RECT 2691.310 3367.850 2691.610 3368.910 ;
        RECT 2739.150 3368.530 2739.450 3368.910 ;
        RECT 2787.910 3368.910 2836.050 3369.210 ;
        RECT 2739.150 3368.230 2787.290 3368.530 ;
        RECT 2690.390 3367.550 2691.610 3367.850 ;
        RECT 2786.990 3367.850 2787.290 3368.230 ;
        RECT 2787.910 3367.850 2788.210 3368.910 ;
        RECT 2835.750 3368.530 2836.050 3368.910 ;
        RECT 2916.710 3368.530 2917.010 3372.990 ;
        RECT 2917.600 3372.540 2924.800 3372.990 ;
        RECT 2835.750 3368.230 2883.890 3368.530 ;
        RECT 2786.990 3367.550 2788.210 3367.850 ;
        RECT 2883.590 3367.850 2883.890 3368.230 ;
        RECT 2884.510 3368.230 2917.010 3368.530 ;
        RECT 2884.510 3367.850 2884.810 3368.230 ;
        RECT 2883.590 3367.550 2884.810 3367.850 ;
        RECT 1800.965 3367.535 1801.295 3367.550 ;
        RECT 2429.325 3367.535 2429.655 3367.550 ;
        RECT 2463.110 3367.540 2463.490 3367.550 ;
        RECT 695.790 1497.850 696.170 1497.860 ;
        RECT 715.810 1497.850 719.810 1497.855 ;
        RECT 695.790 1497.550 719.810 1497.850 ;
        RECT 695.790 1497.540 696.170 1497.550 ;
        RECT 715.810 1497.255 719.810 1497.550 ;
      LAYER via3 ;
        RECT 695.820 3368.900 696.140 3369.220 ;
        RECT 2463.140 3368.900 2463.460 3369.220 ;
        RECT 2463.140 3367.540 2463.460 3367.860 ;
        RECT 695.820 1497.540 696.140 1497.860 ;
      LAYER met4 ;
        RECT 695.815 3368.895 696.145 3369.225 ;
        RECT 2463.135 3368.895 2463.465 3369.225 ;
        RECT 695.830 1497.865 696.130 3368.895 ;
        RECT 2463.150 3367.865 2463.450 3368.895 ;
        RECT 2463.135 3367.535 2463.465 3367.865 ;
        RECT 695.815 1497.535 696.145 1497.865 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 862.110 3501.560 862.430 3501.620 ;
        RECT 2798.250 3501.560 2798.570 3501.620 ;
        RECT 862.110 3501.420 2798.570 3501.560 ;
        RECT 862.110 3501.360 862.430 3501.420 ;
        RECT 2798.250 3501.360 2798.570 3501.420 ;
      LAYER via ;
        RECT 862.140 3501.360 862.400 3501.620 ;
        RECT 2798.280 3501.360 2798.540 3501.620 ;
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
        RECT 2798.340 3501.650 2798.480 3517.600 ;
        RECT 862.140 3501.330 862.400 3501.650 ;
        RECT 2798.280 3501.330 2798.540 3501.650 ;
        RECT 860.340 2377.690 860.620 2377.880 ;
        RECT 862.200 2377.690 862.340 3501.330 ;
        RECT 860.340 2377.550 862.340 2377.690 ;
        RECT 860.340 2373.880 860.620 2377.550 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2470.345 3332.765 2470.515 3380.875 ;
        RECT 2470.345 3236.205 2470.515 3284.315 ;
        RECT 2471.265 3139.645 2471.435 3187.755 ;
        RECT 2471.265 3043.085 2471.435 3091.195 ;
        RECT 2471.265 2946.525 2471.435 2994.635 ;
        RECT 2470.805 2815.285 2470.975 2849.455 ;
        RECT 2471.725 2214.845 2471.895 2270.095 ;
        RECT 2472.185 2118.285 2472.355 2166.395 ;
        RECT 2471.265 2021.725 2471.435 2069.835 ;
        RECT 2471.265 1883.685 2471.435 1931.795 ;
        RECT 2472.185 1787.125 2472.355 1835.235 ;
        RECT 2471.725 1690.565 2471.895 1738.675 ;
        RECT 2471.265 1594.005 2471.435 1642.115 ;
        RECT 2470.805 1497.445 2470.975 1545.555 ;
      LAYER mcon ;
        RECT 2470.345 3380.705 2470.515 3380.875 ;
        RECT 2470.345 3284.145 2470.515 3284.315 ;
        RECT 2471.265 3187.585 2471.435 3187.755 ;
        RECT 2471.265 3091.025 2471.435 3091.195 ;
        RECT 2471.265 2994.465 2471.435 2994.635 ;
        RECT 2470.805 2849.285 2470.975 2849.455 ;
        RECT 2471.725 2269.925 2471.895 2270.095 ;
        RECT 2472.185 2166.225 2472.355 2166.395 ;
        RECT 2471.265 2069.665 2471.435 2069.835 ;
        RECT 2471.265 1931.625 2471.435 1931.795 ;
        RECT 2472.185 1835.065 2472.355 1835.235 ;
        RECT 2471.725 1738.505 2471.895 1738.675 ;
        RECT 2471.265 1641.945 2471.435 1642.115 ;
        RECT 2470.805 1545.385 2470.975 1545.555 ;
      LAYER met1 ;
        RECT 2470.270 3380.860 2470.590 3380.920 ;
        RECT 2470.075 3380.720 2470.590 3380.860 ;
        RECT 2470.270 3380.660 2470.590 3380.720 ;
        RECT 2470.285 3332.920 2470.575 3332.965 ;
        RECT 2471.190 3332.920 2471.510 3332.980 ;
        RECT 2470.285 3332.780 2471.510 3332.920 ;
        RECT 2470.285 3332.735 2470.575 3332.780 ;
        RECT 2471.190 3332.720 2471.510 3332.780 ;
        RECT 2470.270 3284.300 2470.590 3284.360 ;
        RECT 2470.075 3284.160 2470.590 3284.300 ;
        RECT 2470.270 3284.100 2470.590 3284.160 ;
        RECT 2470.285 3236.360 2470.575 3236.405 ;
        RECT 2470.730 3236.360 2471.050 3236.420 ;
        RECT 2470.285 3236.220 2471.050 3236.360 ;
        RECT 2470.285 3236.175 2470.575 3236.220 ;
        RECT 2470.730 3236.160 2471.050 3236.220 ;
        RECT 2471.205 3187.740 2471.495 3187.785 ;
        RECT 2471.650 3187.740 2471.970 3187.800 ;
        RECT 2471.205 3187.600 2471.970 3187.740 ;
        RECT 2471.205 3187.555 2471.495 3187.600 ;
        RECT 2471.650 3187.540 2471.970 3187.600 ;
        RECT 2471.190 3139.800 2471.510 3139.860 ;
        RECT 2470.995 3139.660 2471.510 3139.800 ;
        RECT 2471.190 3139.600 2471.510 3139.660 ;
        RECT 2471.205 3091.180 2471.495 3091.225 ;
        RECT 2471.650 3091.180 2471.970 3091.240 ;
        RECT 2471.205 3091.040 2471.970 3091.180 ;
        RECT 2471.205 3090.995 2471.495 3091.040 ;
        RECT 2471.650 3090.980 2471.970 3091.040 ;
        RECT 2471.190 3043.240 2471.510 3043.300 ;
        RECT 2470.995 3043.100 2471.510 3043.240 ;
        RECT 2471.190 3043.040 2471.510 3043.100 ;
        RECT 2471.205 2994.620 2471.495 2994.665 ;
        RECT 2471.650 2994.620 2471.970 2994.680 ;
        RECT 2471.205 2994.480 2471.970 2994.620 ;
        RECT 2471.205 2994.435 2471.495 2994.480 ;
        RECT 2471.650 2994.420 2471.970 2994.480 ;
        RECT 2471.190 2946.680 2471.510 2946.740 ;
        RECT 2470.995 2946.540 2471.510 2946.680 ;
        RECT 2471.190 2946.480 2471.510 2946.540 ;
        RECT 2470.270 2900.440 2470.590 2900.500 ;
        RECT 2471.190 2900.440 2471.510 2900.500 ;
        RECT 2470.270 2900.300 2471.510 2900.440 ;
        RECT 2470.270 2900.240 2470.590 2900.300 ;
        RECT 2471.190 2900.240 2471.510 2900.300 ;
        RECT 2470.730 2849.440 2471.050 2849.500 ;
        RECT 2470.535 2849.300 2471.050 2849.440 ;
        RECT 2470.730 2849.240 2471.050 2849.300 ;
        RECT 2470.745 2815.440 2471.035 2815.485 ;
        RECT 2471.650 2815.440 2471.970 2815.500 ;
        RECT 2470.745 2815.300 2471.970 2815.440 ;
        RECT 2470.745 2815.255 2471.035 2815.300 ;
        RECT 2471.650 2815.240 2471.970 2815.300 ;
        RECT 2470.730 2753.220 2471.050 2753.280 ;
        RECT 2472.110 2753.220 2472.430 2753.280 ;
        RECT 2470.730 2753.080 2472.430 2753.220 ;
        RECT 2470.730 2753.020 2471.050 2753.080 ;
        RECT 2472.110 2753.020 2472.430 2753.080 ;
        RECT 2472.110 2719.220 2472.430 2719.280 ;
        RECT 2471.740 2719.080 2472.430 2719.220 ;
        RECT 2471.740 2718.600 2471.880 2719.080 ;
        RECT 2472.110 2719.020 2472.430 2719.080 ;
        RECT 2471.650 2718.340 2471.970 2718.600 ;
        RECT 2470.730 2656.660 2471.050 2656.720 ;
        RECT 2472.110 2656.660 2472.430 2656.720 ;
        RECT 2470.730 2656.520 2472.430 2656.660 ;
        RECT 2470.730 2656.460 2471.050 2656.520 ;
        RECT 2472.110 2656.460 2472.430 2656.520 ;
        RECT 2472.110 2622.660 2472.430 2622.720 ;
        RECT 2471.740 2622.520 2472.430 2622.660 ;
        RECT 2471.740 2622.040 2471.880 2622.520 ;
        RECT 2472.110 2622.460 2472.430 2622.520 ;
        RECT 2471.650 2621.780 2471.970 2622.040 ;
        RECT 2470.730 2560.100 2471.050 2560.160 ;
        RECT 2472.110 2560.100 2472.430 2560.160 ;
        RECT 2470.730 2559.960 2472.430 2560.100 ;
        RECT 2470.730 2559.900 2471.050 2559.960 ;
        RECT 2472.110 2559.900 2472.430 2559.960 ;
        RECT 2472.110 2526.100 2472.430 2526.160 ;
        RECT 2471.740 2525.960 2472.430 2526.100 ;
        RECT 2471.740 2525.480 2471.880 2525.960 ;
        RECT 2472.110 2525.900 2472.430 2525.960 ;
        RECT 2471.650 2525.220 2471.970 2525.480 ;
        RECT 2471.190 2428.860 2471.510 2428.920 ;
        RECT 2471.190 2428.720 2471.880 2428.860 ;
        RECT 2471.190 2428.660 2471.510 2428.720 ;
        RECT 2471.740 2428.580 2471.880 2428.720 ;
        RECT 2471.650 2428.320 2471.970 2428.580 ;
        RECT 2471.650 2414.920 2471.970 2414.980 ;
        RECT 2472.570 2414.920 2472.890 2414.980 ;
        RECT 2471.650 2414.780 2472.890 2414.920 ;
        RECT 2471.650 2414.720 2471.970 2414.780 ;
        RECT 2472.570 2414.720 2472.890 2414.780 ;
        RECT 2471.190 2332.100 2471.510 2332.360 ;
        RECT 2471.280 2331.960 2471.420 2332.100 ;
        RECT 2472.110 2331.960 2472.430 2332.020 ;
        RECT 2471.280 2331.820 2472.430 2331.960 ;
        RECT 2472.110 2331.760 2472.430 2331.820 ;
        RECT 2471.190 2284.020 2471.510 2284.080 ;
        RECT 2472.110 2284.020 2472.430 2284.080 ;
        RECT 2471.190 2283.880 2472.430 2284.020 ;
        RECT 2471.190 2283.820 2471.510 2283.880 ;
        RECT 2472.110 2283.820 2472.430 2283.880 ;
        RECT 2471.650 2270.080 2471.970 2270.140 ;
        RECT 2471.455 2269.940 2471.970 2270.080 ;
        RECT 2471.650 2269.880 2471.970 2269.940 ;
        RECT 2471.665 2215.000 2471.955 2215.045 ;
        RECT 2472.110 2215.000 2472.430 2215.060 ;
        RECT 2471.665 2214.860 2472.430 2215.000 ;
        RECT 2471.665 2214.815 2471.955 2214.860 ;
        RECT 2472.110 2214.800 2472.430 2214.860 ;
        RECT 2471.190 2187.460 2471.510 2187.520 ;
        RECT 2472.110 2187.460 2472.430 2187.520 ;
        RECT 2471.190 2187.320 2472.430 2187.460 ;
        RECT 2471.190 2187.260 2471.510 2187.320 ;
        RECT 2472.110 2187.260 2472.430 2187.320 ;
        RECT 2472.110 2166.380 2472.430 2166.440 ;
        RECT 2471.915 2166.240 2472.430 2166.380 ;
        RECT 2472.110 2166.180 2472.430 2166.240 ;
        RECT 2472.125 2118.440 2472.415 2118.485 ;
        RECT 2472.570 2118.440 2472.890 2118.500 ;
        RECT 2472.125 2118.300 2472.890 2118.440 ;
        RECT 2472.125 2118.255 2472.415 2118.300 ;
        RECT 2472.570 2118.240 2472.890 2118.300 ;
        RECT 2471.190 2077.640 2471.510 2077.700 ;
        RECT 2472.570 2077.640 2472.890 2077.700 ;
        RECT 2471.190 2077.500 2472.890 2077.640 ;
        RECT 2471.190 2077.440 2471.510 2077.500 ;
        RECT 2472.570 2077.440 2472.890 2077.500 ;
        RECT 2471.190 2069.820 2471.510 2069.880 ;
        RECT 2470.995 2069.680 2471.510 2069.820 ;
        RECT 2471.190 2069.620 2471.510 2069.680 ;
        RECT 2471.205 2021.880 2471.495 2021.925 ;
        RECT 2472.110 2021.880 2472.430 2021.940 ;
        RECT 2471.205 2021.740 2472.430 2021.880 ;
        RECT 2471.205 2021.695 2471.495 2021.740 ;
        RECT 2472.110 2021.680 2472.430 2021.740 ;
        RECT 2471.190 1931.780 2471.510 1931.840 ;
        RECT 2470.995 1931.640 2471.510 1931.780 ;
        RECT 2471.190 1931.580 2471.510 1931.640 ;
        RECT 2471.205 1883.840 2471.495 1883.885 ;
        RECT 2472.570 1883.840 2472.890 1883.900 ;
        RECT 2471.205 1883.700 2472.890 1883.840 ;
        RECT 2471.205 1883.655 2471.495 1883.700 ;
        RECT 2472.570 1883.640 2472.890 1883.700 ;
        RECT 2471.650 1849.160 2471.970 1849.220 ;
        RECT 2472.570 1849.160 2472.890 1849.220 ;
        RECT 2471.650 1849.020 2472.890 1849.160 ;
        RECT 2471.650 1848.960 2471.970 1849.020 ;
        RECT 2472.570 1848.960 2472.890 1849.020 ;
        RECT 2472.125 1835.220 2472.415 1835.265 ;
        RECT 2472.570 1835.220 2472.890 1835.280 ;
        RECT 2472.125 1835.080 2472.890 1835.220 ;
        RECT 2472.125 1835.035 2472.415 1835.080 ;
        RECT 2472.570 1835.020 2472.890 1835.080 ;
        RECT 2472.110 1787.280 2472.430 1787.340 ;
        RECT 2471.915 1787.140 2472.430 1787.280 ;
        RECT 2472.110 1787.080 2472.430 1787.140 ;
        RECT 2471.190 1752.600 2471.510 1752.660 ;
        RECT 2472.110 1752.600 2472.430 1752.660 ;
        RECT 2471.190 1752.460 2472.430 1752.600 ;
        RECT 2471.190 1752.400 2471.510 1752.460 ;
        RECT 2472.110 1752.400 2472.430 1752.460 ;
        RECT 2471.665 1738.660 2471.955 1738.705 ;
        RECT 2472.110 1738.660 2472.430 1738.720 ;
        RECT 2471.665 1738.520 2472.430 1738.660 ;
        RECT 2471.665 1738.475 2471.955 1738.520 ;
        RECT 2472.110 1738.460 2472.430 1738.520 ;
        RECT 2471.650 1690.720 2471.970 1690.780 ;
        RECT 2471.455 1690.580 2471.970 1690.720 ;
        RECT 2471.650 1690.520 2471.970 1690.580 ;
        RECT 2471.190 1642.100 2471.510 1642.160 ;
        RECT 2470.995 1641.960 2471.510 1642.100 ;
        RECT 2471.190 1641.900 2471.510 1641.960 ;
        RECT 2471.205 1594.160 2471.495 1594.205 ;
        RECT 2472.110 1594.160 2472.430 1594.220 ;
        RECT 2471.205 1594.020 2472.430 1594.160 ;
        RECT 2471.205 1593.975 2471.495 1594.020 ;
        RECT 2472.110 1593.960 2472.430 1594.020 ;
        RECT 2470.730 1559.480 2471.050 1559.540 ;
        RECT 2472.110 1559.480 2472.430 1559.540 ;
        RECT 2470.730 1559.340 2472.430 1559.480 ;
        RECT 2470.730 1559.280 2471.050 1559.340 ;
        RECT 2472.110 1559.280 2472.430 1559.340 ;
        RECT 2470.730 1545.540 2471.050 1545.600 ;
        RECT 2470.730 1545.400 2471.245 1545.540 ;
        RECT 2470.730 1545.340 2471.050 1545.400 ;
        RECT 2470.745 1497.600 2471.035 1497.645 ;
        RECT 2472.110 1497.600 2472.430 1497.660 ;
        RECT 2470.745 1497.460 2472.430 1497.600 ;
        RECT 2470.745 1497.415 2471.035 1497.460 ;
        RECT 2472.110 1497.400 2472.430 1497.460 ;
        RECT 2471.190 1462.920 2471.510 1462.980 ;
        RECT 2472.110 1462.920 2472.430 1462.980 ;
        RECT 2471.190 1462.780 2472.430 1462.920 ;
        RECT 2471.190 1462.720 2471.510 1462.780 ;
        RECT 2472.110 1462.720 2472.430 1462.780 ;
        RECT 926.510 1320.460 926.830 1320.520 ;
        RECT 2471.650 1320.460 2471.970 1320.520 ;
        RECT 926.510 1320.320 2471.970 1320.460 ;
        RECT 926.510 1320.260 926.830 1320.320 ;
        RECT 2471.650 1320.260 2471.970 1320.320 ;
      LAYER via ;
        RECT 2470.300 3380.660 2470.560 3380.920 ;
        RECT 2471.220 3332.720 2471.480 3332.980 ;
        RECT 2470.300 3284.100 2470.560 3284.360 ;
        RECT 2470.760 3236.160 2471.020 3236.420 ;
        RECT 2471.680 3187.540 2471.940 3187.800 ;
        RECT 2471.220 3139.600 2471.480 3139.860 ;
        RECT 2471.680 3090.980 2471.940 3091.240 ;
        RECT 2471.220 3043.040 2471.480 3043.300 ;
        RECT 2471.680 2994.420 2471.940 2994.680 ;
        RECT 2471.220 2946.480 2471.480 2946.740 ;
        RECT 2470.300 2900.240 2470.560 2900.500 ;
        RECT 2471.220 2900.240 2471.480 2900.500 ;
        RECT 2470.760 2849.240 2471.020 2849.500 ;
        RECT 2471.680 2815.240 2471.940 2815.500 ;
        RECT 2470.760 2753.020 2471.020 2753.280 ;
        RECT 2472.140 2753.020 2472.400 2753.280 ;
        RECT 2472.140 2719.020 2472.400 2719.280 ;
        RECT 2471.680 2718.340 2471.940 2718.600 ;
        RECT 2470.760 2656.460 2471.020 2656.720 ;
        RECT 2472.140 2656.460 2472.400 2656.720 ;
        RECT 2472.140 2622.460 2472.400 2622.720 ;
        RECT 2471.680 2621.780 2471.940 2622.040 ;
        RECT 2470.760 2559.900 2471.020 2560.160 ;
        RECT 2472.140 2559.900 2472.400 2560.160 ;
        RECT 2472.140 2525.900 2472.400 2526.160 ;
        RECT 2471.680 2525.220 2471.940 2525.480 ;
        RECT 2471.220 2428.660 2471.480 2428.920 ;
        RECT 2471.680 2428.320 2471.940 2428.580 ;
        RECT 2471.680 2414.720 2471.940 2414.980 ;
        RECT 2472.600 2414.720 2472.860 2414.980 ;
        RECT 2471.220 2332.100 2471.480 2332.360 ;
        RECT 2472.140 2331.760 2472.400 2332.020 ;
        RECT 2471.220 2283.820 2471.480 2284.080 ;
        RECT 2472.140 2283.820 2472.400 2284.080 ;
        RECT 2471.680 2269.880 2471.940 2270.140 ;
        RECT 2472.140 2214.800 2472.400 2215.060 ;
        RECT 2471.220 2187.260 2471.480 2187.520 ;
        RECT 2472.140 2187.260 2472.400 2187.520 ;
        RECT 2472.140 2166.180 2472.400 2166.440 ;
        RECT 2472.600 2118.240 2472.860 2118.500 ;
        RECT 2471.220 2077.440 2471.480 2077.700 ;
        RECT 2472.600 2077.440 2472.860 2077.700 ;
        RECT 2471.220 2069.620 2471.480 2069.880 ;
        RECT 2472.140 2021.680 2472.400 2021.940 ;
        RECT 2471.220 1931.580 2471.480 1931.840 ;
        RECT 2472.600 1883.640 2472.860 1883.900 ;
        RECT 2471.680 1848.960 2471.940 1849.220 ;
        RECT 2472.600 1848.960 2472.860 1849.220 ;
        RECT 2472.600 1835.020 2472.860 1835.280 ;
        RECT 2472.140 1787.080 2472.400 1787.340 ;
        RECT 2471.220 1752.400 2471.480 1752.660 ;
        RECT 2472.140 1752.400 2472.400 1752.660 ;
        RECT 2472.140 1738.460 2472.400 1738.720 ;
        RECT 2471.680 1690.520 2471.940 1690.780 ;
        RECT 2471.220 1641.900 2471.480 1642.160 ;
        RECT 2472.140 1593.960 2472.400 1594.220 ;
        RECT 2470.760 1559.280 2471.020 1559.540 ;
        RECT 2472.140 1559.280 2472.400 1559.540 ;
        RECT 2470.760 1545.340 2471.020 1545.600 ;
        RECT 2472.140 1497.400 2472.400 1497.660 ;
        RECT 2471.220 1462.720 2471.480 1462.980 ;
        RECT 2472.140 1462.720 2472.400 1462.980 ;
        RECT 926.540 1320.260 926.800 1320.520 ;
        RECT 2471.680 1320.260 2471.940 1320.520 ;
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
        RECT 2474.040 3517.370 2474.180 3517.600 ;
        RECT 2474.040 3517.230 2475.100 3517.370 ;
        RECT 2474.960 3430.445 2475.100 3517.230 ;
        RECT 2474.890 3430.075 2475.170 3430.445 ;
        RECT 2471.210 3429.395 2471.490 3429.765 ;
        RECT 2471.280 3394.970 2471.420 3429.395 ;
        RECT 2470.360 3394.830 2471.420 3394.970 ;
        RECT 2470.360 3380.950 2470.500 3394.830 ;
        RECT 2470.300 3380.630 2470.560 3380.950 ;
        RECT 2471.220 3332.690 2471.480 3333.010 ;
        RECT 2471.280 3298.410 2471.420 3332.690 ;
        RECT 2470.360 3298.270 2471.420 3298.410 ;
        RECT 2470.360 3284.390 2470.500 3298.270 ;
        RECT 2470.300 3284.070 2470.560 3284.390 ;
        RECT 2470.760 3236.130 2471.020 3236.450 ;
        RECT 2470.820 3201.850 2470.960 3236.130 ;
        RECT 2470.820 3201.710 2471.880 3201.850 ;
        RECT 2471.740 3187.830 2471.880 3201.710 ;
        RECT 2471.680 3187.510 2471.940 3187.830 ;
        RECT 2471.220 3139.570 2471.480 3139.890 ;
        RECT 2471.280 3105.290 2471.420 3139.570 ;
        RECT 2471.280 3105.150 2471.880 3105.290 ;
        RECT 2471.740 3091.270 2471.880 3105.150 ;
        RECT 2471.680 3090.950 2471.940 3091.270 ;
        RECT 2471.220 3043.010 2471.480 3043.330 ;
        RECT 2471.280 3008.730 2471.420 3043.010 ;
        RECT 2471.280 3008.590 2471.880 3008.730 ;
        RECT 2471.740 2994.710 2471.880 3008.590 ;
        RECT 2471.680 2994.390 2471.940 2994.710 ;
        RECT 2471.220 2946.450 2471.480 2946.770 ;
        RECT 2471.280 2900.530 2471.420 2946.450 ;
        RECT 2470.300 2900.210 2470.560 2900.530 ;
        RECT 2471.220 2900.210 2471.480 2900.530 ;
        RECT 2470.360 2863.210 2470.500 2900.210 ;
        RECT 2470.360 2863.070 2470.960 2863.210 ;
        RECT 2470.820 2849.530 2470.960 2863.070 ;
        RECT 2470.760 2849.210 2471.020 2849.530 ;
        RECT 2471.680 2815.210 2471.940 2815.530 ;
        RECT 2471.740 2801.445 2471.880 2815.210 ;
        RECT 2470.750 2801.075 2471.030 2801.445 ;
        RECT 2471.670 2801.075 2471.950 2801.445 ;
        RECT 2470.820 2753.310 2470.960 2801.075 ;
        RECT 2470.760 2752.990 2471.020 2753.310 ;
        RECT 2472.140 2752.990 2472.400 2753.310 ;
        RECT 2472.200 2719.310 2472.340 2752.990 ;
        RECT 2472.140 2718.990 2472.400 2719.310 ;
        RECT 2471.680 2718.310 2471.940 2718.630 ;
        RECT 2471.740 2704.885 2471.880 2718.310 ;
        RECT 2470.750 2704.515 2471.030 2704.885 ;
        RECT 2471.670 2704.515 2471.950 2704.885 ;
        RECT 2470.820 2656.750 2470.960 2704.515 ;
        RECT 2470.760 2656.430 2471.020 2656.750 ;
        RECT 2472.140 2656.430 2472.400 2656.750 ;
        RECT 2472.200 2622.750 2472.340 2656.430 ;
        RECT 2472.140 2622.430 2472.400 2622.750 ;
        RECT 2471.680 2621.750 2471.940 2622.070 ;
        RECT 2471.740 2608.325 2471.880 2621.750 ;
        RECT 2470.750 2607.955 2471.030 2608.325 ;
        RECT 2471.670 2607.955 2471.950 2608.325 ;
        RECT 2470.820 2560.190 2470.960 2607.955 ;
        RECT 2470.760 2559.870 2471.020 2560.190 ;
        RECT 2472.140 2559.870 2472.400 2560.190 ;
        RECT 2472.200 2526.190 2472.340 2559.870 ;
        RECT 2472.140 2525.870 2472.400 2526.190 ;
        RECT 2471.680 2525.190 2471.940 2525.510 ;
        RECT 2471.740 2476.970 2471.880 2525.190 ;
        RECT 2470.820 2476.830 2471.880 2476.970 ;
        RECT 2470.820 2438.890 2470.960 2476.830 ;
        RECT 2470.820 2438.750 2471.420 2438.890 ;
        RECT 2471.280 2428.950 2471.420 2438.750 ;
        RECT 2471.220 2428.630 2471.480 2428.950 ;
        RECT 2471.680 2428.290 2471.940 2428.610 ;
        RECT 2471.740 2415.010 2471.880 2428.290 ;
        RECT 2471.680 2414.690 2471.940 2415.010 ;
        RECT 2472.600 2414.690 2472.860 2415.010 ;
        RECT 2472.660 2366.925 2472.800 2414.690 ;
        RECT 2471.210 2366.555 2471.490 2366.925 ;
        RECT 2472.590 2366.555 2472.870 2366.925 ;
        RECT 2471.280 2332.390 2471.420 2366.555 ;
        RECT 2471.220 2332.070 2471.480 2332.390 ;
        RECT 2472.140 2331.730 2472.400 2332.050 ;
        RECT 2472.200 2284.110 2472.340 2331.730 ;
        RECT 2471.220 2283.850 2471.480 2284.110 ;
        RECT 2471.220 2283.790 2471.880 2283.850 ;
        RECT 2472.140 2283.790 2472.400 2284.110 ;
        RECT 2471.280 2283.710 2471.880 2283.790 ;
        RECT 2471.740 2270.170 2471.880 2283.710 ;
        RECT 2471.680 2269.850 2471.940 2270.170 ;
        RECT 2472.140 2214.770 2472.400 2215.090 ;
        RECT 2472.200 2187.550 2472.340 2214.770 ;
        RECT 2471.220 2187.290 2471.480 2187.550 ;
        RECT 2472.140 2187.290 2472.400 2187.550 ;
        RECT 2471.220 2187.230 2472.400 2187.290 ;
        RECT 2471.280 2187.150 2472.340 2187.230 ;
        RECT 2472.200 2166.470 2472.340 2187.150 ;
        RECT 2472.140 2166.150 2472.400 2166.470 ;
        RECT 2472.600 2118.210 2472.860 2118.530 ;
        RECT 2472.660 2077.730 2472.800 2118.210 ;
        RECT 2471.220 2077.410 2471.480 2077.730 ;
        RECT 2472.600 2077.410 2472.860 2077.730 ;
        RECT 2471.280 2069.910 2471.420 2077.410 ;
        RECT 2471.220 2069.590 2471.480 2069.910 ;
        RECT 2472.140 2021.650 2472.400 2021.970 ;
        RECT 2472.200 1994.170 2472.340 2021.650 ;
        RECT 2471.280 1994.030 2472.340 1994.170 ;
        RECT 2471.280 1931.870 2471.420 1994.030 ;
        RECT 2471.220 1931.550 2471.480 1931.870 ;
        RECT 2472.600 1883.610 2472.860 1883.930 ;
        RECT 2472.660 1849.330 2472.800 1883.610 ;
        RECT 2471.740 1849.250 2472.800 1849.330 ;
        RECT 2471.680 1849.190 2472.860 1849.250 ;
        RECT 2471.680 1848.930 2471.940 1849.190 ;
        RECT 2472.600 1848.930 2472.860 1849.190 ;
        RECT 2472.660 1835.310 2472.800 1848.930 ;
        RECT 2472.600 1834.990 2472.860 1835.310 ;
        RECT 2472.140 1787.050 2472.400 1787.370 ;
        RECT 2472.200 1752.770 2472.340 1787.050 ;
        RECT 2471.280 1752.690 2472.340 1752.770 ;
        RECT 2471.220 1752.630 2472.400 1752.690 ;
        RECT 2471.220 1752.370 2471.480 1752.630 ;
        RECT 2472.140 1752.370 2472.400 1752.630 ;
        RECT 2472.200 1738.750 2472.340 1752.370 ;
        RECT 2472.140 1738.430 2472.400 1738.750 ;
        RECT 2471.680 1690.490 2471.940 1690.810 ;
        RECT 2471.740 1656.210 2471.880 1690.490 ;
        RECT 2471.280 1656.070 2471.880 1656.210 ;
        RECT 2471.280 1642.190 2471.420 1656.070 ;
        RECT 2471.220 1641.870 2471.480 1642.190 ;
        RECT 2472.140 1593.930 2472.400 1594.250 ;
        RECT 2472.200 1559.570 2472.340 1593.930 ;
        RECT 2470.760 1559.250 2471.020 1559.570 ;
        RECT 2472.140 1559.250 2472.400 1559.570 ;
        RECT 2470.820 1545.630 2470.960 1559.250 ;
        RECT 2470.760 1545.310 2471.020 1545.630 ;
        RECT 2472.140 1497.370 2472.400 1497.690 ;
        RECT 2472.200 1463.010 2472.340 1497.370 ;
        RECT 2471.220 1462.690 2471.480 1463.010 ;
        RECT 2472.140 1462.690 2472.400 1463.010 ;
        RECT 2471.280 1414.810 2471.420 1462.690 ;
        RECT 2471.280 1414.670 2471.880 1414.810 ;
        RECT 926.580 1323.135 926.860 1327.135 ;
        RECT 926.600 1320.550 926.740 1323.135 ;
        RECT 2471.740 1320.550 2471.880 1414.670 ;
        RECT 926.540 1320.230 926.800 1320.550 ;
        RECT 2471.680 1320.230 2471.940 1320.550 ;
      LAYER via2 ;
        RECT 2474.890 3430.120 2475.170 3430.400 ;
        RECT 2471.210 3429.440 2471.490 3429.720 ;
        RECT 2470.750 2801.120 2471.030 2801.400 ;
        RECT 2471.670 2801.120 2471.950 2801.400 ;
        RECT 2470.750 2704.560 2471.030 2704.840 ;
        RECT 2471.670 2704.560 2471.950 2704.840 ;
        RECT 2470.750 2608.000 2471.030 2608.280 ;
        RECT 2471.670 2608.000 2471.950 2608.280 ;
        RECT 2471.210 2366.600 2471.490 2366.880 ;
        RECT 2472.590 2366.600 2472.870 2366.880 ;
      LAYER met3 ;
        RECT 2474.865 3430.410 2475.195 3430.425 ;
        RECT 2470.510 3430.110 2475.195 3430.410 ;
        RECT 2470.510 3429.730 2470.810 3430.110 ;
        RECT 2474.865 3430.095 2475.195 3430.110 ;
        RECT 2471.185 3429.730 2471.515 3429.745 ;
        RECT 2470.510 3429.430 2471.515 3429.730 ;
        RECT 2471.185 3429.415 2471.515 3429.430 ;
        RECT 2470.725 2801.410 2471.055 2801.425 ;
        RECT 2471.645 2801.410 2471.975 2801.425 ;
        RECT 2470.725 2801.110 2471.975 2801.410 ;
        RECT 2470.725 2801.095 2471.055 2801.110 ;
        RECT 2471.645 2801.095 2471.975 2801.110 ;
        RECT 2470.725 2704.850 2471.055 2704.865 ;
        RECT 2471.645 2704.850 2471.975 2704.865 ;
        RECT 2470.725 2704.550 2471.975 2704.850 ;
        RECT 2470.725 2704.535 2471.055 2704.550 ;
        RECT 2471.645 2704.535 2471.975 2704.550 ;
        RECT 2470.725 2608.290 2471.055 2608.305 ;
        RECT 2471.645 2608.290 2471.975 2608.305 ;
        RECT 2470.725 2607.990 2471.975 2608.290 ;
        RECT 2470.725 2607.975 2471.055 2607.990 ;
        RECT 2471.645 2607.975 2471.975 2607.990 ;
        RECT 2471.185 2366.890 2471.515 2366.905 ;
        RECT 2472.565 2366.890 2472.895 2366.905 ;
        RECT 2471.185 2366.590 2472.895 2366.890 ;
        RECT 2471.185 2366.575 2471.515 2366.590 ;
        RECT 2472.565 2366.575 2472.895 2366.590 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1331.310 3503.260 1331.630 3503.320 ;
        RECT 2149.190 3503.260 2149.510 3503.320 ;
        RECT 1331.310 3503.120 2149.510 3503.260 ;
        RECT 1331.310 3503.060 1331.630 3503.120 ;
        RECT 2149.190 3503.060 2149.510 3503.120 ;
      LAYER via ;
        RECT 1331.340 3503.060 1331.600 3503.320 ;
        RECT 2149.220 3503.060 2149.480 3503.320 ;
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
        RECT 2149.280 3503.350 2149.420 3517.600 ;
        RECT 1331.340 3503.030 1331.600 3503.350 ;
        RECT 2149.220 3503.030 2149.480 3503.350 ;
        RECT 1328.620 2377.010 1328.900 2377.880 ;
        RECT 1331.400 2377.010 1331.540 3503.030 ;
        RECT 1328.620 2376.870 1331.540 2377.010 ;
        RECT 1328.620 2373.880 1328.900 2376.870 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1822.205 3332.765 1822.375 3380.875 ;
        RECT 1821.745 3236.205 1821.915 3284.315 ;
        RECT 1822.665 3139.645 1822.835 3187.755 ;
        RECT 1822.665 3043.085 1822.835 3091.195 ;
        RECT 1822.665 2946.525 1822.835 2994.635 ;
        RECT 1822.205 2815.285 1822.375 2849.455 ;
        RECT 1822.205 2428.365 1822.375 2463.215 ;
        RECT 1822.205 2318.885 1822.375 2366.655 ;
        RECT 1822.665 2235.245 1822.835 2265.675 ;
        RECT 1824.045 2084.965 1824.215 2125.255 ;
        RECT 1824.045 2028.525 1824.215 2076.975 ;
        RECT 1822.665 1883.685 1822.835 1931.795 ;
        RECT 1823.125 1594.345 1823.295 1642.115 ;
        RECT 1823.125 1497.785 1823.295 1545.555 ;
        RECT 1822.665 1462.425 1822.835 1463.275 ;
      LAYER mcon ;
        RECT 1822.205 3380.705 1822.375 3380.875 ;
        RECT 1821.745 3284.145 1821.915 3284.315 ;
        RECT 1822.665 3187.585 1822.835 3187.755 ;
        RECT 1822.665 3091.025 1822.835 3091.195 ;
        RECT 1822.665 2994.465 1822.835 2994.635 ;
        RECT 1822.205 2849.285 1822.375 2849.455 ;
        RECT 1822.205 2463.045 1822.375 2463.215 ;
        RECT 1822.205 2366.485 1822.375 2366.655 ;
        RECT 1822.665 2265.505 1822.835 2265.675 ;
        RECT 1824.045 2125.085 1824.215 2125.255 ;
        RECT 1824.045 2076.805 1824.215 2076.975 ;
        RECT 1822.665 1931.625 1822.835 1931.795 ;
        RECT 1823.125 1641.945 1823.295 1642.115 ;
        RECT 1823.125 1545.385 1823.295 1545.555 ;
        RECT 1822.665 1463.105 1822.835 1463.275 ;
      LAYER met1 ;
        RECT 1822.130 3464.160 1822.450 3464.220 ;
        RECT 1825.350 3464.160 1825.670 3464.220 ;
        RECT 1822.130 3464.020 1825.670 3464.160 ;
        RECT 1822.130 3463.960 1822.450 3464.020 ;
        RECT 1825.350 3463.960 1825.670 3464.020 ;
        RECT 1822.130 3380.860 1822.450 3380.920 ;
        RECT 1821.935 3380.720 1822.450 3380.860 ;
        RECT 1822.130 3380.660 1822.450 3380.720 ;
        RECT 1822.145 3332.920 1822.435 3332.965 ;
        RECT 1822.590 3332.920 1822.910 3332.980 ;
        RECT 1822.145 3332.780 1822.910 3332.920 ;
        RECT 1822.145 3332.735 1822.435 3332.780 ;
        RECT 1822.590 3332.720 1822.910 3332.780 ;
        RECT 1821.670 3284.300 1821.990 3284.360 ;
        RECT 1821.475 3284.160 1821.990 3284.300 ;
        RECT 1821.670 3284.100 1821.990 3284.160 ;
        RECT 1821.685 3236.360 1821.975 3236.405 ;
        RECT 1822.130 3236.360 1822.450 3236.420 ;
        RECT 1821.685 3236.220 1822.450 3236.360 ;
        RECT 1821.685 3236.175 1821.975 3236.220 ;
        RECT 1822.130 3236.160 1822.450 3236.220 ;
        RECT 1822.605 3187.740 1822.895 3187.785 ;
        RECT 1823.050 3187.740 1823.370 3187.800 ;
        RECT 1822.605 3187.600 1823.370 3187.740 ;
        RECT 1822.605 3187.555 1822.895 3187.600 ;
        RECT 1823.050 3187.540 1823.370 3187.600 ;
        RECT 1822.590 3139.800 1822.910 3139.860 ;
        RECT 1822.395 3139.660 1822.910 3139.800 ;
        RECT 1822.590 3139.600 1822.910 3139.660 ;
        RECT 1822.605 3091.180 1822.895 3091.225 ;
        RECT 1823.050 3091.180 1823.370 3091.240 ;
        RECT 1822.605 3091.040 1823.370 3091.180 ;
        RECT 1822.605 3090.995 1822.895 3091.040 ;
        RECT 1823.050 3090.980 1823.370 3091.040 ;
        RECT 1822.590 3043.240 1822.910 3043.300 ;
        RECT 1822.395 3043.100 1822.910 3043.240 ;
        RECT 1822.590 3043.040 1822.910 3043.100 ;
        RECT 1822.605 2994.620 1822.895 2994.665 ;
        RECT 1823.050 2994.620 1823.370 2994.680 ;
        RECT 1822.605 2994.480 1823.370 2994.620 ;
        RECT 1822.605 2994.435 1822.895 2994.480 ;
        RECT 1823.050 2994.420 1823.370 2994.480 ;
        RECT 1822.590 2946.680 1822.910 2946.740 ;
        RECT 1822.395 2946.540 1822.910 2946.680 ;
        RECT 1822.590 2946.480 1822.910 2946.540 ;
        RECT 1821.670 2900.440 1821.990 2900.500 ;
        RECT 1822.590 2900.440 1822.910 2900.500 ;
        RECT 1821.670 2900.300 1822.910 2900.440 ;
        RECT 1821.670 2900.240 1821.990 2900.300 ;
        RECT 1822.590 2900.240 1822.910 2900.300 ;
        RECT 1822.130 2849.440 1822.450 2849.500 ;
        RECT 1821.935 2849.300 1822.450 2849.440 ;
        RECT 1822.130 2849.240 1822.450 2849.300 ;
        RECT 1822.145 2815.440 1822.435 2815.485 ;
        RECT 1823.050 2815.440 1823.370 2815.500 ;
        RECT 1822.145 2815.300 1823.370 2815.440 ;
        RECT 1822.145 2815.255 1822.435 2815.300 ;
        RECT 1823.050 2815.240 1823.370 2815.300 ;
        RECT 1822.130 2753.220 1822.450 2753.280 ;
        RECT 1823.510 2753.220 1823.830 2753.280 ;
        RECT 1822.130 2753.080 1823.830 2753.220 ;
        RECT 1822.130 2753.020 1822.450 2753.080 ;
        RECT 1823.510 2753.020 1823.830 2753.080 ;
        RECT 1823.510 2719.220 1823.830 2719.280 ;
        RECT 1823.140 2719.080 1823.830 2719.220 ;
        RECT 1823.140 2718.600 1823.280 2719.080 ;
        RECT 1823.510 2719.020 1823.830 2719.080 ;
        RECT 1823.050 2718.340 1823.370 2718.600 ;
        RECT 1822.130 2656.660 1822.450 2656.720 ;
        RECT 1823.510 2656.660 1823.830 2656.720 ;
        RECT 1822.130 2656.520 1823.830 2656.660 ;
        RECT 1822.130 2656.460 1822.450 2656.520 ;
        RECT 1823.510 2656.460 1823.830 2656.520 ;
        RECT 1823.510 2622.660 1823.830 2622.720 ;
        RECT 1823.140 2622.520 1823.830 2622.660 ;
        RECT 1823.140 2622.040 1823.280 2622.520 ;
        RECT 1823.510 2622.460 1823.830 2622.520 ;
        RECT 1823.050 2621.780 1823.370 2622.040 ;
        RECT 1822.130 2560.100 1822.450 2560.160 ;
        RECT 1823.510 2560.100 1823.830 2560.160 ;
        RECT 1822.130 2559.960 1823.830 2560.100 ;
        RECT 1822.130 2559.900 1822.450 2559.960 ;
        RECT 1823.510 2559.900 1823.830 2559.960 ;
        RECT 1823.510 2526.100 1823.830 2526.160 ;
        RECT 1823.140 2525.960 1823.830 2526.100 ;
        RECT 1823.140 2525.480 1823.280 2525.960 ;
        RECT 1823.510 2525.900 1823.830 2525.960 ;
        RECT 1823.050 2525.220 1823.370 2525.480 ;
        RECT 1822.130 2463.200 1822.450 2463.260 ;
        RECT 1821.935 2463.060 1822.450 2463.200 ;
        RECT 1822.130 2463.000 1822.450 2463.060 ;
        RECT 1822.145 2428.520 1822.435 2428.565 ;
        RECT 1822.590 2428.520 1822.910 2428.580 ;
        RECT 1822.145 2428.380 1822.910 2428.520 ;
        RECT 1822.145 2428.335 1822.435 2428.380 ;
        RECT 1822.590 2428.320 1822.910 2428.380 ;
        RECT 1822.145 2366.640 1822.435 2366.685 ;
        RECT 1823.050 2366.640 1823.370 2366.700 ;
        RECT 1822.145 2366.500 1823.370 2366.640 ;
        RECT 1822.145 2366.455 1822.435 2366.500 ;
        RECT 1823.050 2366.440 1823.370 2366.500 ;
        RECT 1822.130 2319.040 1822.450 2319.100 ;
        RECT 1821.935 2318.900 1822.450 2319.040 ;
        RECT 1822.130 2318.840 1822.450 2318.900 ;
        RECT 1821.210 2318.360 1821.530 2318.420 ;
        RECT 1822.130 2318.360 1822.450 2318.420 ;
        RECT 1821.210 2318.220 1822.450 2318.360 ;
        RECT 1821.210 2318.160 1821.530 2318.220 ;
        RECT 1822.130 2318.160 1822.450 2318.220 ;
        RECT 1822.590 2265.660 1822.910 2265.720 ;
        RECT 1822.395 2265.520 1822.910 2265.660 ;
        RECT 1822.590 2265.460 1822.910 2265.520 ;
        RECT 1822.605 2235.400 1822.895 2235.445 ;
        RECT 1823.510 2235.400 1823.830 2235.460 ;
        RECT 1822.605 2235.260 1823.830 2235.400 ;
        RECT 1822.605 2235.215 1822.895 2235.260 ;
        RECT 1823.510 2235.200 1823.830 2235.260 ;
        RECT 1824.430 2149.380 1824.750 2149.440 ;
        RECT 1825.350 2149.380 1825.670 2149.440 ;
        RECT 1824.430 2149.240 1825.670 2149.380 ;
        RECT 1824.430 2149.180 1824.750 2149.240 ;
        RECT 1825.350 2149.180 1825.670 2149.240 ;
        RECT 1823.970 2125.240 1824.290 2125.300 ;
        RECT 1823.775 2125.100 1824.290 2125.240 ;
        RECT 1823.970 2125.040 1824.290 2125.100 ;
        RECT 1823.970 2085.120 1824.290 2085.180 ;
        RECT 1823.775 2084.980 1824.290 2085.120 ;
        RECT 1823.970 2084.920 1824.290 2084.980 ;
        RECT 1823.970 2076.960 1824.290 2077.020 ;
        RECT 1823.775 2076.820 1824.290 2076.960 ;
        RECT 1823.970 2076.760 1824.290 2076.820 ;
        RECT 1823.970 2028.680 1824.290 2028.740 ;
        RECT 1823.775 2028.540 1824.290 2028.680 ;
        RECT 1823.970 2028.480 1824.290 2028.540 ;
        RECT 1823.970 1994.680 1824.290 1994.740 ;
        RECT 1823.600 1994.540 1824.290 1994.680 ;
        RECT 1823.600 1994.060 1823.740 1994.540 ;
        RECT 1823.970 1994.480 1824.290 1994.540 ;
        RECT 1823.510 1993.800 1823.830 1994.060 ;
        RECT 1822.590 1931.780 1822.910 1931.840 ;
        RECT 1822.395 1931.640 1822.910 1931.780 ;
        RECT 1822.590 1931.580 1822.910 1931.640 ;
        RECT 1822.605 1883.840 1822.895 1883.885 ;
        RECT 1823.050 1883.840 1823.370 1883.900 ;
        RECT 1822.605 1883.700 1823.370 1883.840 ;
        RECT 1822.605 1883.655 1822.895 1883.700 ;
        RECT 1823.050 1883.640 1823.370 1883.700 ;
        RECT 1823.050 1849.500 1823.370 1849.560 ;
        RECT 1823.510 1849.500 1823.830 1849.560 ;
        RECT 1823.050 1849.360 1823.830 1849.500 ;
        RECT 1823.050 1849.300 1823.370 1849.360 ;
        RECT 1823.510 1849.300 1823.830 1849.360 ;
        RECT 1823.065 1642.100 1823.355 1642.145 ;
        RECT 1823.510 1642.100 1823.830 1642.160 ;
        RECT 1823.065 1641.960 1823.830 1642.100 ;
        RECT 1823.065 1641.915 1823.355 1641.960 ;
        RECT 1823.510 1641.900 1823.830 1641.960 ;
        RECT 1823.050 1594.500 1823.370 1594.560 ;
        RECT 1822.855 1594.360 1823.370 1594.500 ;
        RECT 1823.050 1594.300 1823.370 1594.360 ;
        RECT 1823.050 1559.820 1823.370 1559.880 ;
        RECT 1823.510 1559.820 1823.830 1559.880 ;
        RECT 1823.050 1559.680 1823.830 1559.820 ;
        RECT 1823.050 1559.620 1823.370 1559.680 ;
        RECT 1823.510 1559.620 1823.830 1559.680 ;
        RECT 1823.065 1545.540 1823.355 1545.585 ;
        RECT 1823.510 1545.540 1823.830 1545.600 ;
        RECT 1823.065 1545.400 1823.830 1545.540 ;
        RECT 1823.065 1545.355 1823.355 1545.400 ;
        RECT 1823.510 1545.340 1823.830 1545.400 ;
        RECT 1823.050 1497.940 1823.370 1498.000 ;
        RECT 1822.855 1497.800 1823.370 1497.940 ;
        RECT 1823.050 1497.740 1823.370 1497.800 ;
        RECT 1822.605 1463.260 1822.895 1463.305 ;
        RECT 1823.050 1463.260 1823.370 1463.320 ;
        RECT 1822.605 1463.120 1823.370 1463.260 ;
        RECT 1822.605 1463.075 1822.895 1463.120 ;
        RECT 1823.050 1463.060 1823.370 1463.120 ;
        RECT 1822.590 1462.580 1822.910 1462.640 ;
        RECT 1822.395 1462.440 1822.910 1462.580 ;
        RECT 1822.590 1462.380 1822.910 1462.440 ;
        RECT 1637.670 1320.120 1637.990 1320.180 ;
        RECT 1823.050 1320.120 1823.370 1320.180 ;
        RECT 1637.670 1319.980 1823.370 1320.120 ;
        RECT 1637.670 1319.920 1637.990 1319.980 ;
        RECT 1823.050 1319.920 1823.370 1319.980 ;
      LAYER via ;
        RECT 1822.160 3463.960 1822.420 3464.220 ;
        RECT 1825.380 3463.960 1825.640 3464.220 ;
        RECT 1822.160 3380.660 1822.420 3380.920 ;
        RECT 1822.620 3332.720 1822.880 3332.980 ;
        RECT 1821.700 3284.100 1821.960 3284.360 ;
        RECT 1822.160 3236.160 1822.420 3236.420 ;
        RECT 1823.080 3187.540 1823.340 3187.800 ;
        RECT 1822.620 3139.600 1822.880 3139.860 ;
        RECT 1823.080 3090.980 1823.340 3091.240 ;
        RECT 1822.620 3043.040 1822.880 3043.300 ;
        RECT 1823.080 2994.420 1823.340 2994.680 ;
        RECT 1822.620 2946.480 1822.880 2946.740 ;
        RECT 1821.700 2900.240 1821.960 2900.500 ;
        RECT 1822.620 2900.240 1822.880 2900.500 ;
        RECT 1822.160 2849.240 1822.420 2849.500 ;
        RECT 1823.080 2815.240 1823.340 2815.500 ;
        RECT 1822.160 2753.020 1822.420 2753.280 ;
        RECT 1823.540 2753.020 1823.800 2753.280 ;
        RECT 1823.540 2719.020 1823.800 2719.280 ;
        RECT 1823.080 2718.340 1823.340 2718.600 ;
        RECT 1822.160 2656.460 1822.420 2656.720 ;
        RECT 1823.540 2656.460 1823.800 2656.720 ;
        RECT 1823.540 2622.460 1823.800 2622.720 ;
        RECT 1823.080 2621.780 1823.340 2622.040 ;
        RECT 1822.160 2559.900 1822.420 2560.160 ;
        RECT 1823.540 2559.900 1823.800 2560.160 ;
        RECT 1823.540 2525.900 1823.800 2526.160 ;
        RECT 1823.080 2525.220 1823.340 2525.480 ;
        RECT 1822.160 2463.000 1822.420 2463.260 ;
        RECT 1822.620 2428.320 1822.880 2428.580 ;
        RECT 1823.080 2366.440 1823.340 2366.700 ;
        RECT 1822.160 2318.840 1822.420 2319.100 ;
        RECT 1821.240 2318.160 1821.500 2318.420 ;
        RECT 1822.160 2318.160 1822.420 2318.420 ;
        RECT 1822.620 2265.460 1822.880 2265.720 ;
        RECT 1823.540 2235.200 1823.800 2235.460 ;
        RECT 1824.460 2149.180 1824.720 2149.440 ;
        RECT 1825.380 2149.180 1825.640 2149.440 ;
        RECT 1824.000 2125.040 1824.260 2125.300 ;
        RECT 1824.000 2084.920 1824.260 2085.180 ;
        RECT 1824.000 2076.760 1824.260 2077.020 ;
        RECT 1824.000 2028.480 1824.260 2028.740 ;
        RECT 1824.000 1994.480 1824.260 1994.740 ;
        RECT 1823.540 1993.800 1823.800 1994.060 ;
        RECT 1822.620 1931.580 1822.880 1931.840 ;
        RECT 1823.080 1883.640 1823.340 1883.900 ;
        RECT 1823.080 1849.300 1823.340 1849.560 ;
        RECT 1823.540 1849.300 1823.800 1849.560 ;
        RECT 1823.540 1641.900 1823.800 1642.160 ;
        RECT 1823.080 1594.300 1823.340 1594.560 ;
        RECT 1823.080 1559.620 1823.340 1559.880 ;
        RECT 1823.540 1559.620 1823.800 1559.880 ;
        RECT 1823.540 1545.340 1823.800 1545.600 ;
        RECT 1823.080 1497.740 1823.340 1498.000 ;
        RECT 1823.080 1463.060 1823.340 1463.320 ;
        RECT 1822.620 1462.380 1822.880 1462.640 ;
        RECT 1637.700 1319.920 1637.960 1320.180 ;
        RECT 1823.080 1319.920 1823.340 1320.180 ;
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
        RECT 1824.980 3517.370 1825.120 3517.600 ;
        RECT 1824.980 3517.230 1825.580 3517.370 ;
        RECT 1825.440 3464.250 1825.580 3517.230 ;
        RECT 1822.160 3463.930 1822.420 3464.250 ;
        RECT 1825.380 3463.930 1825.640 3464.250 ;
        RECT 1822.220 3380.950 1822.360 3463.930 ;
        RECT 1822.160 3380.630 1822.420 3380.950 ;
        RECT 1822.620 3332.690 1822.880 3333.010 ;
        RECT 1822.680 3298.410 1822.820 3332.690 ;
        RECT 1821.760 3298.270 1822.820 3298.410 ;
        RECT 1821.760 3284.390 1821.900 3298.270 ;
        RECT 1821.700 3284.070 1821.960 3284.390 ;
        RECT 1822.160 3236.130 1822.420 3236.450 ;
        RECT 1822.220 3201.850 1822.360 3236.130 ;
        RECT 1822.220 3201.710 1823.280 3201.850 ;
        RECT 1823.140 3187.830 1823.280 3201.710 ;
        RECT 1823.080 3187.510 1823.340 3187.830 ;
        RECT 1822.620 3139.570 1822.880 3139.890 ;
        RECT 1822.680 3105.290 1822.820 3139.570 ;
        RECT 1822.680 3105.150 1823.280 3105.290 ;
        RECT 1823.140 3091.270 1823.280 3105.150 ;
        RECT 1823.080 3090.950 1823.340 3091.270 ;
        RECT 1822.620 3043.010 1822.880 3043.330 ;
        RECT 1822.680 3008.730 1822.820 3043.010 ;
        RECT 1822.680 3008.590 1823.280 3008.730 ;
        RECT 1823.140 2994.710 1823.280 3008.590 ;
        RECT 1823.080 2994.390 1823.340 2994.710 ;
        RECT 1822.620 2946.450 1822.880 2946.770 ;
        RECT 1822.680 2900.530 1822.820 2946.450 ;
        RECT 1821.700 2900.210 1821.960 2900.530 ;
        RECT 1822.620 2900.210 1822.880 2900.530 ;
        RECT 1821.760 2863.210 1821.900 2900.210 ;
        RECT 1821.760 2863.070 1822.360 2863.210 ;
        RECT 1822.220 2849.530 1822.360 2863.070 ;
        RECT 1822.160 2849.210 1822.420 2849.530 ;
        RECT 1823.080 2815.210 1823.340 2815.530 ;
        RECT 1823.140 2801.445 1823.280 2815.210 ;
        RECT 1822.150 2801.075 1822.430 2801.445 ;
        RECT 1823.070 2801.075 1823.350 2801.445 ;
        RECT 1822.220 2753.310 1822.360 2801.075 ;
        RECT 1822.160 2752.990 1822.420 2753.310 ;
        RECT 1823.540 2752.990 1823.800 2753.310 ;
        RECT 1823.600 2719.310 1823.740 2752.990 ;
        RECT 1823.540 2718.990 1823.800 2719.310 ;
        RECT 1823.080 2718.310 1823.340 2718.630 ;
        RECT 1823.140 2704.885 1823.280 2718.310 ;
        RECT 1822.150 2704.515 1822.430 2704.885 ;
        RECT 1823.070 2704.515 1823.350 2704.885 ;
        RECT 1822.220 2656.750 1822.360 2704.515 ;
        RECT 1822.160 2656.430 1822.420 2656.750 ;
        RECT 1823.540 2656.430 1823.800 2656.750 ;
        RECT 1823.600 2622.750 1823.740 2656.430 ;
        RECT 1823.540 2622.430 1823.800 2622.750 ;
        RECT 1823.080 2621.750 1823.340 2622.070 ;
        RECT 1823.140 2608.325 1823.280 2621.750 ;
        RECT 1822.150 2607.955 1822.430 2608.325 ;
        RECT 1823.070 2607.955 1823.350 2608.325 ;
        RECT 1822.220 2560.190 1822.360 2607.955 ;
        RECT 1822.160 2559.870 1822.420 2560.190 ;
        RECT 1823.540 2559.870 1823.800 2560.190 ;
        RECT 1823.600 2526.190 1823.740 2559.870 ;
        RECT 1823.540 2525.870 1823.800 2526.190 ;
        RECT 1823.080 2525.190 1823.340 2525.510 ;
        RECT 1823.140 2476.970 1823.280 2525.190 ;
        RECT 1822.220 2476.830 1823.280 2476.970 ;
        RECT 1822.220 2463.290 1822.360 2476.830 ;
        RECT 1822.160 2462.970 1822.420 2463.290 ;
        RECT 1822.620 2428.290 1822.880 2428.610 ;
        RECT 1822.680 2415.090 1822.820 2428.290 ;
        RECT 1822.680 2414.950 1823.280 2415.090 ;
        RECT 1823.140 2366.730 1823.280 2414.950 ;
        RECT 1823.080 2366.410 1823.340 2366.730 ;
        RECT 1822.160 2318.810 1822.420 2319.130 ;
        RECT 1822.220 2318.450 1822.360 2318.810 ;
        RECT 1821.240 2318.130 1821.500 2318.450 ;
        RECT 1822.160 2318.130 1822.420 2318.450 ;
        RECT 1821.300 2270.365 1821.440 2318.130 ;
        RECT 1821.230 2269.995 1821.510 2270.365 ;
        RECT 1822.610 2269.995 1822.890 2270.365 ;
        RECT 1822.680 2265.750 1822.820 2269.995 ;
        RECT 1822.620 2265.430 1822.880 2265.750 ;
        RECT 1823.540 2235.170 1823.800 2235.490 ;
        RECT 1823.600 2187.290 1823.740 2235.170 ;
        RECT 1823.600 2187.150 1824.660 2187.290 ;
        RECT 1824.520 2149.470 1824.660 2187.150 ;
        RECT 1824.460 2149.150 1824.720 2149.470 ;
        RECT 1825.380 2149.150 1825.640 2149.470 ;
        RECT 1825.440 2125.525 1825.580 2149.150 ;
        RECT 1824.450 2125.410 1824.730 2125.525 ;
        RECT 1824.060 2125.330 1824.730 2125.410 ;
        RECT 1824.000 2125.270 1824.730 2125.330 ;
        RECT 1824.000 2125.010 1824.260 2125.270 ;
        RECT 1824.450 2125.155 1824.730 2125.270 ;
        RECT 1825.370 2125.155 1825.650 2125.525 ;
        RECT 1824.060 2124.855 1824.200 2125.010 ;
        RECT 1824.000 2084.890 1824.260 2085.210 ;
        RECT 1824.060 2077.050 1824.200 2084.890 ;
        RECT 1824.000 2076.730 1824.260 2077.050 ;
        RECT 1824.000 2028.450 1824.260 2028.770 ;
        RECT 1824.060 1994.770 1824.200 2028.450 ;
        RECT 1824.000 1994.450 1824.260 1994.770 ;
        RECT 1823.540 1993.770 1823.800 1994.090 ;
        RECT 1823.600 1945.890 1823.740 1993.770 ;
        RECT 1822.680 1945.750 1823.740 1945.890 ;
        RECT 1822.680 1931.870 1822.820 1945.750 ;
        RECT 1822.620 1931.550 1822.880 1931.870 ;
        RECT 1823.080 1883.610 1823.340 1883.930 ;
        RECT 1823.140 1849.590 1823.280 1883.610 ;
        RECT 1823.080 1849.270 1823.340 1849.590 ;
        RECT 1823.540 1849.270 1823.800 1849.590 ;
        RECT 1823.600 1801.050 1823.740 1849.270 ;
        RECT 1822.680 1800.910 1823.740 1801.050 ;
        RECT 1822.680 1704.490 1822.820 1800.910 ;
        RECT 1822.680 1704.350 1823.740 1704.490 ;
        RECT 1823.600 1642.190 1823.740 1704.350 ;
        RECT 1823.540 1641.870 1823.800 1642.190 ;
        RECT 1823.080 1594.270 1823.340 1594.590 ;
        RECT 1823.140 1559.910 1823.280 1594.270 ;
        RECT 1823.080 1559.590 1823.340 1559.910 ;
        RECT 1823.540 1559.590 1823.800 1559.910 ;
        RECT 1823.600 1545.630 1823.740 1559.590 ;
        RECT 1823.540 1545.310 1823.800 1545.630 ;
        RECT 1823.080 1497.710 1823.340 1498.030 ;
        RECT 1823.140 1463.350 1823.280 1497.710 ;
        RECT 1823.080 1463.030 1823.340 1463.350 ;
        RECT 1822.620 1462.350 1822.880 1462.670 ;
        RECT 1822.680 1414.810 1822.820 1462.350 ;
        RECT 1822.680 1414.670 1823.280 1414.810 ;
        RECT 1637.740 1323.135 1638.020 1327.135 ;
        RECT 1637.760 1320.210 1637.900 1323.135 ;
        RECT 1823.140 1320.210 1823.280 1414.670 ;
        RECT 1637.700 1319.890 1637.960 1320.210 ;
        RECT 1823.080 1319.890 1823.340 1320.210 ;
      LAYER via2 ;
        RECT 1822.150 2801.120 1822.430 2801.400 ;
        RECT 1823.070 2801.120 1823.350 2801.400 ;
        RECT 1822.150 2704.560 1822.430 2704.840 ;
        RECT 1823.070 2704.560 1823.350 2704.840 ;
        RECT 1822.150 2608.000 1822.430 2608.280 ;
        RECT 1823.070 2608.000 1823.350 2608.280 ;
        RECT 1821.230 2270.040 1821.510 2270.320 ;
        RECT 1822.610 2270.040 1822.890 2270.320 ;
        RECT 1824.450 2125.200 1824.730 2125.480 ;
        RECT 1825.370 2125.200 1825.650 2125.480 ;
      LAYER met3 ;
        RECT 1822.125 2801.410 1822.455 2801.425 ;
        RECT 1823.045 2801.410 1823.375 2801.425 ;
        RECT 1822.125 2801.110 1823.375 2801.410 ;
        RECT 1822.125 2801.095 1822.455 2801.110 ;
        RECT 1823.045 2801.095 1823.375 2801.110 ;
        RECT 1822.125 2704.850 1822.455 2704.865 ;
        RECT 1823.045 2704.850 1823.375 2704.865 ;
        RECT 1822.125 2704.550 1823.375 2704.850 ;
        RECT 1822.125 2704.535 1822.455 2704.550 ;
        RECT 1823.045 2704.535 1823.375 2704.550 ;
        RECT 1822.125 2608.290 1822.455 2608.305 ;
        RECT 1823.045 2608.290 1823.375 2608.305 ;
        RECT 1822.125 2607.990 1823.375 2608.290 ;
        RECT 1822.125 2607.975 1822.455 2607.990 ;
        RECT 1823.045 2607.975 1823.375 2607.990 ;
        RECT 1821.205 2270.330 1821.535 2270.345 ;
        RECT 1822.585 2270.330 1822.915 2270.345 ;
        RECT 1821.205 2270.030 1822.915 2270.330 ;
        RECT 1821.205 2270.015 1821.535 2270.030 ;
        RECT 1822.585 2270.015 1822.915 2270.030 ;
        RECT 1824.425 2125.490 1824.755 2125.505 ;
        RECT 1825.345 2125.490 1825.675 2125.505 ;
        RECT 1824.425 2125.190 1825.675 2125.490 ;
        RECT 1824.425 2125.175 1824.755 2125.190 ;
        RECT 1825.345 2125.175 1825.675 2125.190 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1172.610 3504.620 1172.930 3504.680 ;
        RECT 1500.590 3504.620 1500.910 3504.680 ;
        RECT 1172.610 3504.480 1500.910 3504.620 ;
        RECT 1172.610 3504.420 1172.930 3504.480 ;
        RECT 1500.590 3504.420 1500.910 3504.480 ;
        RECT 1166.630 2388.740 1166.950 2388.800 ;
        RECT 1172.610 2388.740 1172.930 2388.800 ;
        RECT 1166.630 2388.600 1172.930 2388.740 ;
        RECT 1166.630 2388.540 1166.950 2388.600 ;
        RECT 1172.610 2388.540 1172.930 2388.600 ;
      LAYER via ;
        RECT 1172.640 3504.420 1172.900 3504.680 ;
        RECT 1500.620 3504.420 1500.880 3504.680 ;
        RECT 1166.660 2388.540 1166.920 2388.800 ;
        RECT 1172.640 2388.540 1172.900 2388.800 ;
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
        RECT 1500.680 3504.710 1500.820 3517.600 ;
        RECT 1172.640 3504.390 1172.900 3504.710 ;
        RECT 1500.620 3504.390 1500.880 3504.710 ;
        RECT 1172.700 2388.830 1172.840 3504.390 ;
        RECT 1166.660 2388.510 1166.920 2388.830 ;
        RECT 1172.640 2388.510 1172.900 2388.830 ;
        RECT 1166.720 2377.880 1166.860 2388.510 ;
        RECT 1166.700 2373.880 1166.980 2377.880 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1771.530 1539.080 1771.850 1539.140 ;
        RECT 1777.510 1539.080 1777.830 1539.140 ;
        RECT 1771.530 1538.940 1777.830 1539.080 ;
        RECT 1771.530 1538.880 1771.850 1538.940 ;
        RECT 1777.510 1538.880 1777.830 1538.940 ;
        RECT 1777.510 324.260 1777.830 324.320 ;
        RECT 2900.370 324.260 2900.690 324.320 ;
        RECT 1777.510 324.120 2900.690 324.260 ;
        RECT 1777.510 324.060 1777.830 324.120 ;
        RECT 2900.370 324.060 2900.690 324.120 ;
      LAYER via ;
        RECT 1771.560 1538.880 1771.820 1539.140 ;
        RECT 1777.540 1538.880 1777.800 1539.140 ;
        RECT 1777.540 324.060 1777.800 324.320 ;
        RECT 2900.400 324.060 2900.660 324.320 ;
      LAYER met2 ;
        RECT 1771.550 1545.115 1771.830 1545.485 ;
        RECT 1771.620 1539.170 1771.760 1545.115 ;
        RECT 1771.560 1538.850 1771.820 1539.170 ;
        RECT 1777.540 1538.850 1777.800 1539.170 ;
        RECT 1777.600 324.350 1777.740 1538.850 ;
        RECT 1777.540 324.030 1777.800 324.350 ;
        RECT 2900.400 324.030 2900.660 324.350 ;
        RECT 2900.460 322.845 2900.600 324.030 ;
        RECT 2900.390 322.475 2900.670 322.845 ;
      LAYER via2 ;
        RECT 1771.550 1545.160 1771.830 1545.440 ;
        RECT 2900.390 322.520 2900.670 322.800 ;
      LAYER met3 ;
        RECT 1755.835 1545.450 1759.835 1545.455 ;
        RECT 1771.525 1545.450 1771.855 1545.465 ;
        RECT 1755.835 1545.150 1771.855 1545.450 ;
        RECT 1755.835 1544.855 1759.835 1545.150 ;
        RECT 1771.525 1545.135 1771.855 1545.150 ;
        RECT 2900.365 322.810 2900.695 322.825 ;
        RECT 2917.600 322.810 2924.800 323.260 ;
        RECT 2900.365 322.510 2924.800 322.810 ;
        RECT 2900.365 322.495 2900.695 322.510 ;
        RECT 2917.600 322.060 2924.800 322.510 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 694.285 1368.925 694.455 1393.575 ;
      LAYER mcon ;
        RECT 694.285 1393.405 694.455 1393.575 ;
      LAYER met1 ;
        RECT 694.210 3503.260 694.530 3503.320 ;
        RECT 1175.830 3503.260 1176.150 3503.320 ;
        RECT 694.210 3503.120 1176.150 3503.260 ;
        RECT 694.210 3503.060 694.530 3503.120 ;
        RECT 1175.830 3503.060 1176.150 3503.120 ;
        RECT 694.210 1393.560 694.530 1393.620 ;
        RECT 694.210 1393.420 694.725 1393.560 ;
        RECT 694.210 1393.360 694.530 1393.420 ;
        RECT 694.210 1369.080 694.530 1369.140 ;
        RECT 694.015 1368.940 694.530 1369.080 ;
        RECT 694.210 1368.880 694.530 1368.940 ;
        RECT 694.210 1325.560 694.530 1325.620 ;
        RECT 786.670 1325.560 786.990 1325.620 ;
        RECT 694.210 1325.420 786.990 1325.560 ;
        RECT 694.210 1325.360 694.530 1325.420 ;
        RECT 786.670 1325.360 786.990 1325.420 ;
      LAYER via ;
        RECT 694.240 3503.060 694.500 3503.320 ;
        RECT 1175.860 3503.060 1176.120 3503.320 ;
        RECT 694.240 1393.360 694.500 1393.620 ;
        RECT 694.240 1368.880 694.500 1369.140 ;
        RECT 694.240 1325.360 694.500 1325.620 ;
        RECT 786.700 1325.360 786.960 1325.620 ;
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
        RECT 1175.920 3503.350 1176.060 3517.600 ;
        RECT 694.240 3503.030 694.500 3503.350 ;
        RECT 1175.860 3503.030 1176.120 3503.350 ;
        RECT 694.300 1393.650 694.440 3503.030 ;
        RECT 694.240 1393.330 694.500 1393.650 ;
        RECT 694.240 1368.850 694.500 1369.170 ;
        RECT 694.300 1325.650 694.440 1368.850 ;
        RECT 787.660 1325.730 787.940 1327.135 ;
        RECT 786.760 1325.650 787.940 1325.730 ;
        RECT 694.240 1325.330 694.500 1325.650 ;
        RECT 786.700 1325.590 787.940 1325.650 ;
        RECT 786.700 1325.330 786.960 1325.590 ;
        RECT 787.660 1323.135 787.940 1325.590 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 712.150 3501.560 712.470 3501.620 ;
        RECT 851.530 3501.560 851.850 3501.620 ;
        RECT 712.150 3501.420 851.850 3501.560 ;
        RECT 712.150 3501.360 712.470 3501.420 ;
        RECT 851.530 3501.360 851.850 3501.420 ;
      LAYER via ;
        RECT 712.180 3501.360 712.440 3501.620 ;
        RECT 851.560 3501.360 851.820 3501.620 ;
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
        RECT 851.620 3501.650 851.760 3517.600 ;
        RECT 712.180 3501.330 712.440 3501.650 ;
        RECT 851.560 3501.330 851.820 3501.650 ;
        RECT 712.240 1754.925 712.380 3501.330 ;
        RECT 712.170 1754.555 712.450 1754.925 ;
      LAYER via2 ;
        RECT 712.170 1754.600 712.450 1754.880 ;
      LAYER met3 ;
        RECT 712.145 1754.890 712.475 1754.905 ;
        RECT 715.810 1754.890 719.810 1754.895 ;
        RECT 712.145 1754.590 719.810 1754.890 ;
        RECT 712.145 1754.575 712.475 1754.590 ;
        RECT 715.810 1754.295 719.810 1754.590 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 527.230 3498.500 527.550 3498.560 ;
        RECT 530.910 3498.500 531.230 3498.560 ;
        RECT 527.230 3498.360 531.230 3498.500 ;
        RECT 527.230 3498.300 527.550 3498.360 ;
        RECT 530.910 3498.300 531.230 3498.360 ;
        RECT 530.910 1320.460 531.230 1320.520 ;
        RECT 909.030 1320.460 909.350 1320.520 ;
        RECT 530.910 1320.320 909.350 1320.460 ;
        RECT 530.910 1320.260 531.230 1320.320 ;
        RECT 909.030 1320.260 909.350 1320.320 ;
      LAYER via ;
        RECT 527.260 3498.300 527.520 3498.560 ;
        RECT 530.940 3498.300 531.200 3498.560 ;
        RECT 530.940 1320.260 531.200 1320.520 ;
        RECT 909.060 1320.260 909.320 1320.520 ;
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
        RECT 527.320 3498.590 527.460 3517.600 ;
        RECT 527.260 3498.270 527.520 3498.590 ;
        RECT 530.940 3498.270 531.200 3498.590 ;
        RECT 531.000 1320.550 531.140 3498.270 ;
        RECT 909.100 1323.135 909.380 1327.135 ;
        RECT 909.120 1320.550 909.260 1323.135 ;
        RECT 530.940 1320.230 531.200 1320.550 ;
        RECT 909.060 1320.230 909.320 1320.550 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 202.470 3502.920 202.790 3502.980 ;
        RECT 1491.390 3502.920 1491.710 3502.980 ;
        RECT 202.470 3502.780 1491.710 3502.920 ;
        RECT 202.470 3502.720 202.790 3502.780 ;
        RECT 1491.390 3502.720 1491.710 3502.780 ;
      LAYER via ;
        RECT 202.500 3502.720 202.760 3502.980 ;
        RECT 1491.420 3502.720 1491.680 3502.980 ;
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
        RECT 202.560 3503.010 202.700 3517.600 ;
        RECT 202.500 3502.690 202.760 3503.010 ;
        RECT 1491.420 3502.690 1491.680 3503.010 ;
        RECT 1491.480 2377.010 1491.620 3502.690 ;
        RECT 1496.980 2377.010 1497.260 2377.880 ;
        RECT 1491.480 2376.870 1497.260 2377.010 ;
        RECT 1496.980 2373.880 1497.260 2376.870 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 18.930 3408.740 19.250 3408.800 ;
        RECT 679.490 3408.740 679.810 3408.800 ;
        RECT 18.930 3408.600 679.810 3408.740 ;
        RECT 18.930 3408.540 19.250 3408.600 ;
        RECT 679.490 3408.540 679.810 3408.600 ;
        RECT 679.490 1321.820 679.810 1321.880 ;
        RECT 1718.630 1321.820 1718.950 1321.880 ;
        RECT 679.490 1321.680 1718.950 1321.820 ;
        RECT 679.490 1321.620 679.810 1321.680 ;
        RECT 1718.630 1321.620 1718.950 1321.680 ;
      LAYER via ;
        RECT 18.960 3408.540 19.220 3408.800 ;
        RECT 679.520 3408.540 679.780 3408.800 ;
        RECT 679.520 1321.620 679.780 1321.880 ;
        RECT 1718.660 1321.620 1718.920 1321.880 ;
      LAYER met2 ;
        RECT 18.950 3411.035 19.230 3411.405 ;
        RECT 19.020 3408.830 19.160 3411.035 ;
        RECT 18.960 3408.510 19.220 3408.830 ;
        RECT 679.520 3408.510 679.780 3408.830 ;
        RECT 679.580 1321.910 679.720 3408.510 ;
        RECT 1718.700 1323.135 1718.980 1327.135 ;
        RECT 1718.720 1321.910 1718.860 1323.135 ;
        RECT 679.520 1321.590 679.780 1321.910 ;
        RECT 1718.660 1321.590 1718.920 1321.910 ;
      LAYER via2 ;
        RECT 18.950 3411.080 19.230 3411.360 ;
      LAYER met3 ;
        RECT -4.800 3411.370 2.400 3411.820 ;
        RECT 18.925 3411.370 19.255 3411.385 ;
        RECT -4.800 3411.070 19.255 3411.370 ;
        RECT -4.800 3410.620 2.400 3411.070 ;
        RECT 18.925 3411.055 19.255 3411.070 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 19.390 3119.060 19.710 3119.120 ;
        RECT 24.910 3119.060 25.230 3119.120 ;
        RECT 19.390 3118.920 25.230 3119.060 ;
        RECT 19.390 3118.860 19.710 3118.920 ;
        RECT 24.910 3118.860 25.230 3118.920 ;
        RECT 24.910 1635.300 25.230 1635.360 ;
        RECT 707.550 1635.300 707.870 1635.360 ;
        RECT 24.910 1635.160 707.870 1635.300 ;
        RECT 24.910 1635.100 25.230 1635.160 ;
        RECT 707.550 1635.100 707.870 1635.160 ;
      LAYER via ;
        RECT 19.420 3118.860 19.680 3119.120 ;
        RECT 24.940 3118.860 25.200 3119.120 ;
        RECT 24.940 1635.100 25.200 1635.360 ;
        RECT 707.580 1635.100 707.840 1635.360 ;
      LAYER met2 ;
        RECT 19.410 3124.075 19.690 3124.445 ;
        RECT 19.480 3119.150 19.620 3124.075 ;
        RECT 19.420 3118.830 19.680 3119.150 ;
        RECT 24.940 3118.830 25.200 3119.150 ;
        RECT 25.000 1635.390 25.140 3118.830 ;
        RECT 24.940 1635.070 25.200 1635.390 ;
        RECT 707.580 1635.245 707.840 1635.390 ;
        RECT 707.570 1634.875 707.850 1635.245 ;
      LAYER via2 ;
        RECT 19.410 3124.120 19.690 3124.400 ;
        RECT 707.570 1634.920 707.850 1635.200 ;
      LAYER met3 ;
        RECT -4.800 3124.410 2.400 3124.860 ;
        RECT 19.385 3124.410 19.715 3124.425 ;
        RECT -4.800 3124.110 19.715 3124.410 ;
        RECT -4.800 3123.660 2.400 3124.110 ;
        RECT 19.385 3124.095 19.715 3124.110 ;
        RECT 707.545 1635.210 707.875 1635.225 ;
        RECT 715.810 1635.210 719.810 1635.215 ;
        RECT 707.545 1634.910 719.810 1635.210 ;
        RECT 707.545 1634.895 707.875 1634.910 ;
        RECT 715.810 1634.615 719.810 1634.910 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 18.010 1319.100 18.330 1319.160 ;
        RECT 828.070 1319.100 828.390 1319.160 ;
        RECT 18.010 1318.960 828.390 1319.100 ;
        RECT 18.010 1318.900 18.330 1318.960 ;
        RECT 828.070 1318.900 828.390 1318.960 ;
      LAYER via ;
        RECT 18.040 1318.900 18.300 1319.160 ;
        RECT 828.100 1318.900 828.360 1319.160 ;
      LAYER met2 ;
        RECT 18.030 2836.435 18.310 2836.805 ;
        RECT 18.100 1319.190 18.240 2836.435 ;
        RECT 828.140 1323.135 828.420 1327.135 ;
        RECT 828.160 1319.190 828.300 1323.135 ;
        RECT 18.040 1318.870 18.300 1319.190 ;
        RECT 828.100 1318.870 828.360 1319.190 ;
      LAYER via2 ;
        RECT 18.030 2836.480 18.310 2836.760 ;
      LAYER met3 ;
        RECT -4.800 2836.770 2.400 2837.220 ;
        RECT 18.005 2836.770 18.335 2836.785 ;
        RECT -4.800 2836.470 18.335 2836.770 ;
        RECT -4.800 2836.020 2.400 2836.470 ;
        RECT 18.005 2836.455 18.335 2836.470 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 16.630 2549.560 16.950 2549.620 ;
        RECT 27.210 2549.560 27.530 2549.620 ;
        RECT 16.630 2549.420 27.530 2549.560 ;
        RECT 16.630 2549.360 16.950 2549.420 ;
        RECT 27.210 2549.360 27.530 2549.420 ;
        RECT 27.210 1773.340 27.530 1773.400 ;
        RECT 692.370 1773.340 692.690 1773.400 ;
        RECT 27.210 1773.200 692.690 1773.340 ;
        RECT 27.210 1773.140 27.530 1773.200 ;
        RECT 692.370 1773.140 692.690 1773.200 ;
      LAYER via ;
        RECT 16.660 2549.360 16.920 2549.620 ;
        RECT 27.240 2549.360 27.500 2549.620 ;
        RECT 27.240 1773.140 27.500 1773.400 ;
        RECT 692.400 1773.140 692.660 1773.400 ;
      LAYER met2 ;
        RECT 16.650 2549.475 16.930 2549.845 ;
        RECT 16.660 2549.330 16.920 2549.475 ;
        RECT 27.240 2549.330 27.500 2549.650 ;
        RECT 27.300 1773.430 27.440 2549.330 ;
        RECT 27.240 1773.110 27.500 1773.430 ;
        RECT 692.400 1773.110 692.660 1773.430 ;
        RECT 692.460 1771.245 692.600 1773.110 ;
        RECT 692.390 1770.875 692.670 1771.245 ;
      LAYER via2 ;
        RECT 16.650 2549.520 16.930 2549.800 ;
        RECT 692.390 1770.920 692.670 1771.200 ;
      LAYER met3 ;
        RECT -4.800 2549.810 2.400 2550.260 ;
        RECT 16.625 2549.810 16.955 2549.825 ;
        RECT -4.800 2549.510 16.955 2549.810 ;
        RECT -4.800 2549.060 2.400 2549.510 ;
        RECT 16.625 2549.495 16.955 2549.510 ;
        RECT 692.365 1771.210 692.695 1771.225 ;
        RECT 715.810 1771.210 719.810 1771.215 ;
        RECT 692.365 1770.910 719.810 1771.210 ;
        RECT 692.365 1770.895 692.695 1770.910 ;
        RECT 715.810 1770.615 719.810 1770.910 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.950 2367.235 19.230 2367.605 ;
        RECT 1766.490 2367.235 1766.770 2367.605 ;
        RECT 19.020 2262.205 19.160 2367.235 ;
        RECT 18.950 2261.835 19.230 2262.205 ;
        RECT 1766.560 2152.045 1766.700 2367.235 ;
        RECT 1766.490 2151.675 1766.770 2152.045 ;
      LAYER via2 ;
        RECT 18.950 2367.280 19.230 2367.560 ;
        RECT 1766.490 2367.280 1766.770 2367.560 ;
        RECT 18.950 2261.880 19.230 2262.160 ;
        RECT 1766.490 2151.720 1766.770 2152.000 ;
      LAYER met3 ;
        RECT 18.925 2367.570 19.255 2367.585 ;
        RECT 1766.465 2367.570 1766.795 2367.585 ;
        RECT 18.925 2367.270 1766.795 2367.570 ;
        RECT 18.925 2367.255 19.255 2367.270 ;
        RECT 1766.465 2367.255 1766.795 2367.270 ;
        RECT -4.800 2262.170 2.400 2262.620 ;
        RECT 18.925 2262.170 19.255 2262.185 ;
        RECT -4.800 2261.870 19.255 2262.170 ;
        RECT -4.800 2261.420 2.400 2261.870 ;
        RECT 18.925 2261.855 19.255 2261.870 ;
        RECT 1755.835 2152.010 1759.835 2152.015 ;
        RECT 1766.465 2152.010 1766.795 2152.025 ;
        RECT 1755.835 2151.710 1766.795 2152.010 ;
        RECT 1755.835 2151.415 1759.835 2151.710 ;
        RECT 1766.465 2151.695 1766.795 2151.710 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 19.390 1318.420 19.710 1318.480 ;
        RECT 943.990 1318.420 944.310 1318.480 ;
        RECT 19.390 1318.280 944.310 1318.420 ;
        RECT 19.390 1318.220 19.710 1318.280 ;
        RECT 943.990 1318.220 944.310 1318.280 ;
      LAYER via ;
        RECT 19.420 1318.220 19.680 1318.480 ;
        RECT 944.020 1318.220 944.280 1318.480 ;
      LAYER met2 ;
        RECT 19.410 1974.875 19.690 1975.245 ;
        RECT 19.480 1318.510 19.620 1974.875 ;
        RECT 944.060 1323.135 944.340 1327.135 ;
        RECT 944.080 1318.510 944.220 1323.135 ;
        RECT 19.420 1318.190 19.680 1318.510 ;
        RECT 944.020 1318.190 944.280 1318.510 ;
      LAYER via2 ;
        RECT 19.410 1974.920 19.690 1975.200 ;
      LAYER met3 ;
        RECT -4.800 1975.210 2.400 1975.660 ;
        RECT 19.385 1975.210 19.715 1975.225 ;
        RECT -4.800 1974.910 19.715 1975.210 ;
        RECT -4.800 1974.460 2.400 1974.910 ;
        RECT 19.385 1974.895 19.715 1974.910 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 718.130 2152.100 718.450 2152.160 ;
        RECT 719.510 2152.100 719.830 2152.160 ;
        RECT 718.130 2151.960 719.830 2152.100 ;
        RECT 718.130 2151.900 718.450 2151.960 ;
        RECT 719.510 2151.900 719.830 2151.960 ;
        RECT 1070.950 553.420 1071.270 553.480 ;
        RECT 1110.510 553.420 1110.830 553.480 ;
        RECT 1070.950 553.280 1110.830 553.420 ;
        RECT 1070.950 553.220 1071.270 553.280 ;
        RECT 1110.510 553.220 1110.830 553.280 ;
        RECT 1750.370 553.420 1750.690 553.480 ;
        RECT 1755.890 553.420 1756.210 553.480 ;
        RECT 1750.370 553.280 1756.210 553.420 ;
        RECT 1750.370 553.220 1750.690 553.280 ;
        RECT 1755.890 553.220 1756.210 553.280 ;
        RECT 1993.710 553.420 1994.030 553.480 ;
        RECT 2028.210 553.420 2028.530 553.480 ;
        RECT 1993.710 553.280 2028.530 553.420 ;
        RECT 1993.710 553.220 1994.030 553.280 ;
        RECT 2028.210 553.220 2028.530 553.280 ;
        RECT 2283.510 553.420 2283.830 553.480 ;
        RECT 2318.010 553.420 2318.330 553.480 ;
        RECT 2283.510 553.280 2318.330 553.420 ;
        RECT 2283.510 553.220 2283.830 553.280 ;
        RECT 2318.010 553.220 2318.330 553.280 ;
        RECT 1220.910 553.080 1221.230 553.140 ;
        RECT 1255.410 553.080 1255.730 553.140 ;
        RECT 1220.910 552.940 1255.730 553.080 ;
        RECT 1220.910 552.880 1221.230 552.940 ;
        RECT 1255.410 552.880 1255.730 552.940 ;
        RECT 1796.370 553.080 1796.690 553.140 ;
        RECT 1835.010 553.080 1835.330 553.140 ;
        RECT 1796.370 552.940 1835.330 553.080 ;
        RECT 1796.370 552.880 1796.690 552.940 ;
        RECT 1835.010 552.880 1835.330 552.940 ;
        RECT 1607.310 552.740 1607.630 552.800 ;
        RECT 1641.810 552.740 1642.130 552.800 ;
        RECT 1607.310 552.600 1642.130 552.740 ;
        RECT 1607.310 552.540 1607.630 552.600 ;
        RECT 1641.810 552.540 1642.130 552.600 ;
      LAYER via ;
        RECT 718.160 2151.900 718.420 2152.160 ;
        RECT 719.540 2151.900 719.800 2152.160 ;
        RECT 1070.980 553.220 1071.240 553.480 ;
        RECT 1110.540 553.220 1110.800 553.480 ;
        RECT 1750.400 553.220 1750.660 553.480 ;
        RECT 1755.920 553.220 1756.180 553.480 ;
        RECT 1993.740 553.220 1994.000 553.480 ;
        RECT 2028.240 553.220 2028.500 553.480 ;
        RECT 2283.540 553.220 2283.800 553.480 ;
        RECT 2318.040 553.220 2318.300 553.480 ;
        RECT 1220.940 552.880 1221.200 553.140 ;
        RECT 1255.440 552.880 1255.700 553.140 ;
        RECT 1796.400 552.880 1796.660 553.140 ;
        RECT 1835.040 552.880 1835.300 553.140 ;
        RECT 1607.340 552.540 1607.600 552.800 ;
        RECT 1641.840 552.540 1642.100 552.800 ;
      LAYER met2 ;
        RECT 718.150 2221.715 718.430 2222.085 ;
        RECT 718.220 2152.190 718.360 2221.715 ;
        RECT 718.160 2151.870 718.420 2152.190 ;
        RECT 719.540 2151.870 719.800 2152.190 ;
        RECT 719.070 2100.250 719.350 2100.365 ;
        RECT 719.600 2100.250 719.740 2151.870 ;
        RECT 719.070 2100.110 719.740 2100.250 ;
        RECT 719.070 2099.995 719.350 2100.110 ;
        RECT 713.090 1857.235 713.370 1857.605 ;
        RECT 713.160 1817.485 713.300 1857.235 ;
        RECT 713.090 1817.115 713.370 1817.485 ;
        RECT 710.330 1661.395 710.610 1661.765 ;
        RECT 710.400 1631.165 710.540 1661.395 ;
        RECT 710.330 1630.795 710.610 1631.165 ;
        RECT 717.230 1542.395 717.510 1542.765 ;
        RECT 717.300 1518.285 717.440 1542.395 ;
        RECT 717.230 1517.915 717.510 1518.285 ;
        RECT 729.190 1322.755 729.470 1323.125 ;
        RECT 729.260 1180.325 729.400 1322.755 ;
        RECT 729.190 1179.955 729.470 1180.325 ;
        RECT 726.430 631.195 726.710 631.565 ;
        RECT 726.500 552.685 726.640 631.195 ;
        RECT 965.630 555.035 965.910 555.405 ;
        RECT 965.700 554.045 965.840 555.035 ;
        RECT 1973.030 554.355 1973.310 554.725 ;
        RECT 965.630 553.675 965.910 554.045 ;
        RECT 1110.530 553.675 1110.810 554.045 ;
        RECT 1414.130 553.930 1414.410 554.045 ;
        RECT 1690.130 553.930 1690.410 554.045 ;
        RECT 1414.130 553.790 1415.260 553.930 ;
        RECT 1414.130 553.675 1414.410 553.790 ;
        RECT 1110.600 553.510 1110.740 553.675 ;
        RECT 1070.980 553.190 1071.240 553.510 ;
        RECT 1110.540 553.190 1110.800 553.510 ;
        RECT 1071.040 552.685 1071.180 553.190 ;
        RECT 1220.930 552.995 1221.210 553.365 ;
        RECT 1220.940 552.850 1221.200 552.995 ;
        RECT 1255.440 552.850 1255.700 553.170 ;
        RECT 1255.500 552.685 1255.640 552.850 ;
        RECT 1415.120 552.685 1415.260 553.790 ;
        RECT 1689.740 553.790 1690.410 553.930 ;
        RECT 1607.330 552.995 1607.610 553.365 ;
        RECT 1607.400 552.830 1607.540 552.995 ;
        RECT 726.430 552.315 726.710 552.685 ;
        RECT 1070.970 552.315 1071.250 552.685 ;
        RECT 1255.430 552.315 1255.710 552.685 ;
        RECT 1415.050 552.315 1415.330 552.685 ;
        RECT 1607.340 552.510 1607.600 552.830 ;
        RECT 1641.840 552.685 1642.100 552.830 ;
        RECT 1689.740 552.685 1689.880 553.790 ;
        RECT 1690.130 553.675 1690.410 553.790 ;
        RECT 1755.910 553.675 1756.190 554.045 ;
        RECT 1796.390 553.675 1796.670 554.045 ;
        RECT 1897.130 553.675 1897.410 554.045 ;
        RECT 1755.980 553.510 1756.120 553.675 ;
        RECT 1750.400 553.365 1750.660 553.510 ;
        RECT 1750.390 552.995 1750.670 553.365 ;
        RECT 1755.920 553.190 1756.180 553.510 ;
        RECT 1796.460 553.170 1796.600 553.675 ;
        RECT 1897.200 553.250 1897.340 553.675 ;
        RECT 1898.050 553.250 1898.330 553.365 ;
        RECT 1796.400 552.850 1796.660 553.170 ;
        RECT 1835.040 552.850 1835.300 553.170 ;
        RECT 1897.200 553.110 1898.330 553.250 ;
        RECT 1898.050 552.995 1898.330 553.110 ;
        RECT 1835.100 552.685 1835.240 552.850 ;
        RECT 1973.100 552.685 1973.240 554.355 ;
        RECT 2028.230 553.675 2028.510 554.045 ;
        RECT 2138.170 553.675 2138.450 554.045 ;
        RECT 2207.630 553.675 2207.910 554.045 ;
        RECT 2318.030 553.675 2318.310 554.045 ;
        RECT 2607.370 553.675 2607.650 554.045 ;
        RECT 2608.290 553.675 2608.570 554.045 ;
        RECT 2028.300 553.510 2028.440 553.675 ;
        RECT 1993.740 553.365 1994.000 553.510 ;
        RECT 1993.730 552.995 1994.010 553.365 ;
        RECT 2028.240 553.190 2028.500 553.510 ;
        RECT 2138.240 553.250 2138.380 553.675 ;
        RECT 2139.550 553.250 2139.830 553.365 ;
        RECT 2138.240 553.110 2139.830 553.250 ;
        RECT 2139.550 552.995 2139.830 553.110 ;
        RECT 1641.830 552.315 1642.110 552.685 ;
        RECT 1689.670 552.315 1689.950 552.685 ;
        RECT 1835.030 552.315 1835.310 552.685 ;
        RECT 1973.030 552.315 1973.310 552.685 ;
        RECT 2207.700 552.005 2207.840 553.675 ;
        RECT 2318.100 553.510 2318.240 553.675 ;
        RECT 2283.540 553.365 2283.800 553.510 ;
        RECT 2283.530 552.995 2283.810 553.365 ;
        RECT 2318.040 553.190 2318.300 553.510 ;
        RECT 2207.630 551.635 2207.910 552.005 ;
        RECT 2607.440 551.325 2607.580 553.675 ;
        RECT 2608.360 551.325 2608.500 553.675 ;
        RECT 2607.370 550.955 2607.650 551.325 ;
        RECT 2608.290 550.955 2608.570 551.325 ;
      LAYER via2 ;
        RECT 718.150 2221.760 718.430 2222.040 ;
        RECT 719.070 2100.040 719.350 2100.320 ;
        RECT 713.090 1857.280 713.370 1857.560 ;
        RECT 713.090 1817.160 713.370 1817.440 ;
        RECT 710.330 1661.440 710.610 1661.720 ;
        RECT 710.330 1630.840 710.610 1631.120 ;
        RECT 717.230 1542.440 717.510 1542.720 ;
        RECT 717.230 1517.960 717.510 1518.240 ;
        RECT 729.190 1322.800 729.470 1323.080 ;
        RECT 729.190 1180.000 729.470 1180.280 ;
        RECT 726.430 631.240 726.710 631.520 ;
        RECT 965.630 555.080 965.910 555.360 ;
        RECT 1973.030 554.400 1973.310 554.680 ;
        RECT 965.630 553.720 965.910 554.000 ;
        RECT 1110.530 553.720 1110.810 554.000 ;
        RECT 1414.130 553.720 1414.410 554.000 ;
        RECT 1220.930 553.040 1221.210 553.320 ;
        RECT 1607.330 553.040 1607.610 553.320 ;
        RECT 726.430 552.360 726.710 552.640 ;
        RECT 1070.970 552.360 1071.250 552.640 ;
        RECT 1255.430 552.360 1255.710 552.640 ;
        RECT 1415.050 552.360 1415.330 552.640 ;
        RECT 1690.130 553.720 1690.410 554.000 ;
        RECT 1755.910 553.720 1756.190 554.000 ;
        RECT 1796.390 553.720 1796.670 554.000 ;
        RECT 1897.130 553.720 1897.410 554.000 ;
        RECT 1750.390 553.040 1750.670 553.320 ;
        RECT 1898.050 553.040 1898.330 553.320 ;
        RECT 2028.230 553.720 2028.510 554.000 ;
        RECT 2138.170 553.720 2138.450 554.000 ;
        RECT 2207.630 553.720 2207.910 554.000 ;
        RECT 2318.030 553.720 2318.310 554.000 ;
        RECT 2607.370 553.720 2607.650 554.000 ;
        RECT 2608.290 553.720 2608.570 554.000 ;
        RECT 1993.730 553.040 1994.010 553.320 ;
        RECT 2139.550 553.040 2139.830 553.320 ;
        RECT 1641.830 552.360 1642.110 552.640 ;
        RECT 1689.670 552.360 1689.950 552.640 ;
        RECT 1835.030 552.360 1835.310 552.640 ;
        RECT 1973.030 552.360 1973.310 552.640 ;
        RECT 2283.530 553.040 2283.810 553.320 ;
        RECT 2207.630 551.680 2207.910 551.960 ;
        RECT 2607.370 551.000 2607.650 551.280 ;
        RECT 2608.290 551.000 2608.570 551.280 ;
      LAYER met3 ;
        RECT 715.810 2360.855 719.810 2361.455 ;
        RECT 718.830 2358.740 719.130 2360.855 ;
        RECT 718.790 2358.420 719.170 2358.740 ;
        RECT 718.125 2222.050 718.455 2222.065 ;
        RECT 719.020 2222.050 719.400 2222.060 ;
        RECT 718.125 2221.750 719.400 2222.050 ;
        RECT 718.125 2221.735 718.455 2221.750 ;
        RECT 719.020 2221.740 719.400 2221.750 ;
        RECT 719.045 2100.340 719.375 2100.345 ;
        RECT 718.790 2100.330 719.375 2100.340 ;
        RECT 718.590 2100.030 719.375 2100.330 ;
        RECT 718.790 2100.020 719.375 2100.030 ;
        RECT 719.045 2100.015 719.375 2100.020 ;
        RECT 714.190 2040.490 714.570 2040.500 ;
        RECT 718.790 2040.490 719.170 2040.500 ;
        RECT 714.190 2040.190 719.170 2040.490 ;
        RECT 714.190 2040.180 714.570 2040.190 ;
        RECT 718.790 2040.180 719.170 2040.190 ;
        RECT 712.350 1964.330 712.730 1964.340 ;
        RECT 714.190 1964.330 714.570 1964.340 ;
        RECT 712.350 1964.030 714.570 1964.330 ;
        RECT 712.350 1964.020 712.730 1964.030 ;
        RECT 714.190 1964.020 714.570 1964.030 ;
        RECT 712.350 1904.490 712.730 1904.500 ;
        RECT 717.870 1904.490 718.250 1904.500 ;
        RECT 712.350 1904.190 718.250 1904.490 ;
        RECT 712.350 1904.180 712.730 1904.190 ;
        RECT 717.870 1904.180 718.250 1904.190 ;
        RECT 713.065 1857.570 713.395 1857.585 ;
        RECT 718.790 1857.570 719.170 1857.580 ;
        RECT 713.065 1857.270 719.170 1857.570 ;
        RECT 713.065 1857.255 713.395 1857.270 ;
        RECT 718.790 1857.260 719.170 1857.270 ;
        RECT 713.065 1817.450 713.395 1817.465 ;
        RECT 718.790 1817.450 719.170 1817.460 ;
        RECT 713.065 1817.150 719.170 1817.450 ;
        RECT 713.065 1817.135 713.395 1817.150 ;
        RECT 718.790 1817.140 719.170 1817.150 ;
        RECT 712.350 1783.450 712.730 1783.460 ;
        RECT 718.790 1783.450 719.170 1783.460 ;
        RECT 712.350 1783.150 719.170 1783.450 ;
        RECT 712.350 1783.140 712.730 1783.150 ;
        RECT 718.790 1783.140 719.170 1783.150 ;
        RECT 712.350 1732.450 712.730 1732.460 ;
        RECT 711.470 1732.150 712.730 1732.450 ;
        RECT 711.470 1731.090 711.770 1732.150 ;
        RECT 712.350 1732.140 712.730 1732.150 ;
        RECT 714.190 1731.090 714.570 1731.100 ;
        RECT 711.470 1730.790 714.570 1731.090 ;
        RECT 714.190 1730.780 714.570 1730.790 ;
        RECT 714.190 1693.690 714.570 1693.700 ;
        RECT 717.870 1693.690 718.250 1693.700 ;
        RECT 714.190 1693.390 718.250 1693.690 ;
        RECT 714.190 1693.380 714.570 1693.390 ;
        RECT 717.870 1693.380 718.250 1693.390 ;
        RECT 710.305 1661.730 710.635 1661.745 ;
        RECT 717.870 1661.730 718.250 1661.740 ;
        RECT 710.305 1661.430 718.250 1661.730 ;
        RECT 710.305 1661.415 710.635 1661.430 ;
        RECT 717.870 1661.420 718.250 1661.430 ;
        RECT 710.305 1631.130 710.635 1631.145 ;
        RECT 718.790 1631.130 719.170 1631.140 ;
        RECT 710.305 1630.830 719.170 1631.130 ;
        RECT 710.305 1630.815 710.635 1630.830 ;
        RECT 718.790 1630.820 719.170 1630.830 ;
        RECT 717.205 1542.730 717.535 1542.745 ;
        RECT 718.790 1542.730 719.170 1542.740 ;
        RECT 717.205 1542.430 719.170 1542.730 ;
        RECT 717.205 1542.415 717.535 1542.430 ;
        RECT 718.790 1542.420 719.170 1542.430 ;
        RECT 717.205 1518.250 717.535 1518.265 ;
        RECT 718.790 1518.250 719.170 1518.260 ;
        RECT 717.205 1517.950 719.170 1518.250 ;
        RECT 717.205 1517.935 717.535 1517.950 ;
        RECT 718.790 1517.940 719.170 1517.950 ;
        RECT 727.070 1323.090 727.450 1323.100 ;
        RECT 729.165 1323.090 729.495 1323.105 ;
        RECT 727.070 1322.790 729.495 1323.090 ;
        RECT 727.070 1322.780 727.450 1322.790 ;
        RECT 729.165 1322.775 729.495 1322.790 ;
        RECT 729.165 1180.300 729.495 1180.305 ;
        RECT 728.910 1180.290 729.495 1180.300 ;
        RECT 728.910 1179.990 729.720 1180.290 ;
        RECT 728.910 1179.980 729.495 1179.990 ;
        RECT 729.165 1179.975 729.495 1179.980 ;
        RECT 726.150 1055.850 726.530 1055.860 ;
        RECT 727.990 1055.850 728.370 1055.860 ;
        RECT 726.150 1055.550 728.370 1055.850 ;
        RECT 726.150 1055.540 726.530 1055.550 ;
        RECT 727.990 1055.540 728.370 1055.550 ;
        RECT 726.150 994.340 726.530 994.660 ;
        RECT 726.190 993.970 726.490 994.340 ;
        RECT 727.070 993.970 727.450 993.980 ;
        RECT 726.190 993.670 727.450 993.970 ;
        RECT 727.070 993.660 727.450 993.670 ;
        RECT 727.070 879.730 727.450 879.740 ;
        RECT 726.190 879.430 727.450 879.730 ;
        RECT 726.190 879.060 726.490 879.430 ;
        RECT 727.070 879.420 727.450 879.430 ;
        RECT 726.150 878.740 726.530 879.060 ;
        RECT 726.150 799.860 726.530 800.180 ;
        RECT 726.190 799.490 726.490 799.860 ;
        RECT 727.990 799.490 728.370 799.500 ;
        RECT 726.190 799.190 728.370 799.490 ;
        RECT 727.990 799.180 728.370 799.190 ;
        RECT 725.230 631.530 725.610 631.540 ;
        RECT 726.405 631.530 726.735 631.545 ;
        RECT 725.230 631.230 726.735 631.530 ;
        RECT 725.230 631.220 725.610 631.230 ;
        RECT 726.405 631.215 726.735 631.230 ;
        RECT 2917.600 557.410 2924.800 557.860 ;
        RECT 2916.710 557.110 2924.800 557.410 ;
        RECT 917.510 555.370 917.890 555.380 ;
        RECT 965.605 555.370 965.935 555.385 ;
        RECT 917.510 555.070 965.935 555.370 ;
        RECT 917.510 555.060 917.890 555.070 ;
        RECT 965.605 555.055 965.935 555.070 ;
        RECT 1544.030 554.690 1544.410 554.700 ;
        RECT 1510.030 554.390 1544.410 554.690 ;
        RECT 1924.910 554.690 1925.290 554.700 ;
        RECT 1973.005 554.690 1973.335 554.705 ;
        RECT 965.605 554.010 965.935 554.025 ;
        RECT 1110.505 554.010 1110.835 554.025 ;
        RECT 1414.105 554.010 1414.435 554.025 ;
        RECT 844.870 553.710 870.010 554.010 ;
        RECT 844.870 553.330 845.170 553.710 ;
        RECT 797.030 553.160 834.130 553.330 ;
        RECT 835.670 553.160 845.170 553.330 ;
        RECT 797.030 553.030 845.170 553.160 ;
        RECT 869.710 553.330 870.010 553.710 ;
        RECT 965.605 553.710 1028.250 554.010 ;
        RECT 965.605 553.695 965.935 553.710 ;
        RECT 917.510 553.330 917.890 553.340 ;
        RECT 869.710 553.030 917.890 553.330 ;
        RECT 726.405 552.650 726.735 552.665 ;
        RECT 797.030 552.650 797.330 553.030 ;
        RECT 833.830 552.860 835.970 553.030 ;
        RECT 917.510 553.020 917.890 553.030 ;
        RECT 726.405 552.350 797.330 552.650 ;
        RECT 1027.950 552.650 1028.250 553.710 ;
        RECT 1110.505 553.710 1124.850 554.010 ;
        RECT 1110.505 553.695 1110.835 553.710 ;
        RECT 1070.945 552.650 1071.275 552.665 ;
        RECT 1027.950 552.350 1071.275 552.650 ;
        RECT 1124.550 552.650 1124.850 553.710 ;
        RECT 1280.030 553.710 1328.170 554.010 ;
        RECT 1220.905 553.330 1221.235 553.345 ;
        RECT 1173.310 553.030 1221.235 553.330 ;
        RECT 1173.310 552.650 1173.610 553.030 ;
        RECT 1220.905 553.015 1221.235 553.030 ;
        RECT 1124.550 552.350 1173.610 552.650 ;
        RECT 1255.405 552.650 1255.735 552.665 ;
        RECT 1280.030 552.650 1280.330 553.710 ;
        RECT 1327.870 553.330 1328.170 553.710 ;
        RECT 1352.710 553.710 1414.435 554.010 ;
        RECT 1352.710 553.330 1353.010 553.710 ;
        RECT 1414.105 553.695 1414.435 553.710 ;
        RECT 1510.030 553.330 1510.330 554.390 ;
        RECT 1544.030 554.380 1544.410 554.390 ;
        RECT 1703.230 554.220 1705.370 554.520 ;
        RECT 1924.910 554.390 1973.335 554.690 ;
        RECT 1924.910 554.380 1925.290 554.390 ;
        RECT 1973.005 554.375 1973.335 554.390 ;
        RECT 1690.105 554.010 1690.435 554.025 ;
        RECT 1703.230 554.010 1703.530 554.220 ;
        RECT 1690.105 553.710 1703.530 554.010 ;
        RECT 1705.070 554.010 1705.370 554.220 ;
        RECT 1755.885 554.010 1756.215 554.025 ;
        RECT 1796.365 554.010 1796.695 554.025 ;
        RECT 1897.105 554.010 1897.435 554.025 ;
        RECT 1705.070 553.710 1714.570 554.010 ;
        RECT 1690.105 553.695 1690.435 553.710 ;
        RECT 1607.305 553.330 1607.635 553.345 ;
        RECT 1327.870 553.030 1353.010 553.330 ;
        RECT 1463.110 553.030 1510.330 553.330 ;
        RECT 1559.710 553.030 1607.635 553.330 ;
        RECT 1714.270 553.330 1714.570 553.710 ;
        RECT 1755.885 553.710 1796.695 554.010 ;
        RECT 1755.885 553.695 1756.215 553.710 ;
        RECT 1796.365 553.695 1796.695 553.710 ;
        RECT 1849.510 553.710 1897.435 554.010 ;
        RECT 1750.365 553.330 1750.695 553.345 ;
        RECT 1714.270 553.030 1750.695 553.330 ;
        RECT 1255.405 552.350 1280.330 552.650 ;
        RECT 1415.025 552.650 1415.355 552.665 ;
        RECT 1463.110 552.650 1463.410 553.030 ;
        RECT 1415.025 552.350 1463.410 552.650 ;
        RECT 1544.950 552.650 1545.330 552.660 ;
        RECT 1559.710 552.650 1560.010 553.030 ;
        RECT 1607.305 553.015 1607.635 553.030 ;
        RECT 1750.365 553.015 1750.695 553.030 ;
        RECT 1544.950 552.350 1560.010 552.650 ;
        RECT 1641.805 552.650 1642.135 552.665 ;
        RECT 1689.645 552.650 1689.975 552.665 ;
        RECT 1641.805 552.350 1689.975 552.650 ;
        RECT 726.405 552.335 726.735 552.350 ;
        RECT 1070.945 552.335 1071.275 552.350 ;
        RECT 1255.405 552.335 1255.735 552.350 ;
        RECT 1415.025 552.335 1415.355 552.350 ;
        RECT 1544.950 552.340 1545.330 552.350 ;
        RECT 1641.805 552.335 1642.135 552.350 ;
        RECT 1689.645 552.335 1689.975 552.350 ;
        RECT 1835.005 552.650 1835.335 552.665 ;
        RECT 1849.510 552.650 1849.810 553.710 ;
        RECT 1897.105 553.695 1897.435 553.710 ;
        RECT 2028.205 554.010 2028.535 554.025 ;
        RECT 2138.145 554.010 2138.475 554.025 ;
        RECT 2028.205 553.710 2138.475 554.010 ;
        RECT 2028.205 553.695 2028.535 553.710 ;
        RECT 2138.145 553.695 2138.475 553.710 ;
        RECT 2207.605 554.010 2207.935 554.025 ;
        RECT 2318.005 554.010 2318.335 554.025 ;
        RECT 2607.345 554.010 2607.675 554.025 ;
        RECT 2608.265 554.010 2608.595 554.025 ;
        RECT 2207.605 553.710 2236.210 554.010 ;
        RECT 2207.605 553.695 2207.935 553.710 ;
        RECT 1898.025 553.330 1898.355 553.345 ;
        RECT 1924.910 553.330 1925.290 553.340 ;
        RECT 1993.705 553.330 1994.035 553.345 ;
        RECT 1898.025 553.030 1925.290 553.330 ;
        RECT 1898.025 553.015 1898.355 553.030 ;
        RECT 1924.910 553.020 1925.290 553.030 ;
        RECT 1980.150 553.030 1994.035 553.330 ;
        RECT 1835.005 552.350 1849.810 552.650 ;
        RECT 1973.005 552.650 1973.335 552.665 ;
        RECT 1980.150 552.650 1980.450 553.030 ;
        RECT 1993.705 553.015 1994.035 553.030 ;
        RECT 2139.525 553.330 2139.855 553.345 ;
        RECT 2173.310 553.330 2173.690 553.340 ;
        RECT 2139.525 553.030 2173.690 553.330 ;
        RECT 2235.910 553.330 2236.210 553.710 ;
        RECT 2318.005 553.710 2380.650 554.010 ;
        RECT 2318.005 553.695 2318.335 553.710 ;
        RECT 2283.505 553.330 2283.835 553.345 ;
        RECT 2235.910 553.030 2283.835 553.330 ;
        RECT 2380.350 553.330 2380.650 553.710 ;
        RECT 2524.790 553.710 2546.250 554.010 ;
        RECT 2524.790 553.330 2525.090 553.710 ;
        RECT 2380.350 553.030 2428.490 553.330 ;
        RECT 2139.525 553.015 2139.855 553.030 ;
        RECT 2173.310 553.020 2173.690 553.030 ;
        RECT 2283.505 553.015 2283.835 553.030 ;
        RECT 1973.005 552.350 1980.450 552.650 ;
        RECT 2428.190 552.650 2428.490 553.030 ;
        RECT 2476.950 553.030 2525.090 553.330 ;
        RECT 2545.950 553.330 2546.250 553.710 ;
        RECT 2607.345 553.710 2608.595 554.010 ;
        RECT 2607.345 553.695 2607.675 553.710 ;
        RECT 2608.265 553.695 2608.595 553.710 ;
        RECT 2656.310 554.010 2656.690 554.020 ;
        RECT 2656.310 553.710 2739.450 554.010 ;
        RECT 2656.310 553.700 2656.690 553.710 ;
        RECT 2559.710 553.330 2560.090 553.340 ;
        RECT 2545.950 553.030 2560.090 553.330 ;
        RECT 2739.150 553.330 2739.450 553.710 ;
        RECT 2787.910 553.710 2836.050 554.010 ;
        RECT 2739.150 553.030 2787.290 553.330 ;
        RECT 2476.950 552.650 2477.250 553.030 ;
        RECT 2559.710 553.020 2560.090 553.030 ;
        RECT 2428.190 552.350 2477.250 552.650 ;
        RECT 2786.990 552.650 2787.290 553.030 ;
        RECT 2787.910 552.650 2788.210 553.710 ;
        RECT 2835.750 553.330 2836.050 553.710 ;
        RECT 2916.710 553.330 2917.010 557.110 ;
        RECT 2917.600 556.660 2924.800 557.110 ;
        RECT 2835.750 553.030 2883.890 553.330 ;
        RECT 2786.990 552.350 2788.210 552.650 ;
        RECT 2883.590 552.650 2883.890 553.030 ;
        RECT 2884.510 553.030 2917.010 553.330 ;
        RECT 2884.510 552.650 2884.810 553.030 ;
        RECT 2883.590 552.350 2884.810 552.650 ;
        RECT 1835.005 552.335 1835.335 552.350 ;
        RECT 1973.005 552.335 1973.335 552.350 ;
        RECT 2173.310 551.970 2173.690 551.980 ;
        RECT 2207.605 551.970 2207.935 551.985 ;
        RECT 2173.310 551.670 2207.935 551.970 ;
        RECT 2173.310 551.660 2173.690 551.670 ;
        RECT 2207.605 551.655 2207.935 551.670 ;
        RECT 2559.710 551.290 2560.090 551.300 ;
        RECT 2607.345 551.290 2607.675 551.305 ;
        RECT 2559.710 550.990 2607.675 551.290 ;
        RECT 2559.710 550.980 2560.090 550.990 ;
        RECT 2607.345 550.975 2607.675 550.990 ;
        RECT 2608.265 551.290 2608.595 551.305 ;
        RECT 2656.310 551.290 2656.690 551.300 ;
        RECT 2608.265 550.990 2656.690 551.290 ;
        RECT 2608.265 550.975 2608.595 550.990 ;
        RECT 2656.310 550.980 2656.690 550.990 ;
      LAYER via3 ;
        RECT 718.820 2358.420 719.140 2358.740 ;
        RECT 719.050 2221.740 719.370 2222.060 ;
        RECT 718.820 2100.020 719.140 2100.340 ;
        RECT 714.220 2040.180 714.540 2040.500 ;
        RECT 718.820 2040.180 719.140 2040.500 ;
        RECT 712.380 1964.020 712.700 1964.340 ;
        RECT 714.220 1964.020 714.540 1964.340 ;
        RECT 712.380 1904.180 712.700 1904.500 ;
        RECT 717.900 1904.180 718.220 1904.500 ;
        RECT 718.820 1857.260 719.140 1857.580 ;
        RECT 718.820 1817.140 719.140 1817.460 ;
        RECT 712.380 1783.140 712.700 1783.460 ;
        RECT 718.820 1783.140 719.140 1783.460 ;
        RECT 712.380 1732.140 712.700 1732.460 ;
        RECT 714.220 1730.780 714.540 1731.100 ;
        RECT 714.220 1693.380 714.540 1693.700 ;
        RECT 717.900 1693.380 718.220 1693.700 ;
        RECT 717.900 1661.420 718.220 1661.740 ;
        RECT 718.820 1630.820 719.140 1631.140 ;
        RECT 718.820 1542.420 719.140 1542.740 ;
        RECT 718.820 1517.940 719.140 1518.260 ;
        RECT 727.100 1322.780 727.420 1323.100 ;
        RECT 728.940 1179.980 729.260 1180.300 ;
        RECT 726.180 1055.540 726.500 1055.860 ;
        RECT 728.020 1055.540 728.340 1055.860 ;
        RECT 726.180 994.340 726.500 994.660 ;
        RECT 727.100 993.660 727.420 993.980 ;
        RECT 727.100 879.420 727.420 879.740 ;
        RECT 726.180 878.740 726.500 879.060 ;
        RECT 726.180 799.860 726.500 800.180 ;
        RECT 728.020 799.180 728.340 799.500 ;
        RECT 725.260 631.220 725.580 631.540 ;
        RECT 917.540 555.060 917.860 555.380 ;
        RECT 917.540 553.020 917.860 553.340 ;
        RECT 1544.060 554.380 1544.380 554.700 ;
        RECT 1924.940 554.380 1925.260 554.700 ;
        RECT 1544.980 552.340 1545.300 552.660 ;
        RECT 1924.940 553.020 1925.260 553.340 ;
        RECT 2173.340 553.020 2173.660 553.340 ;
        RECT 2656.340 553.700 2656.660 554.020 ;
        RECT 2559.740 553.020 2560.060 553.340 ;
        RECT 2173.340 551.660 2173.660 551.980 ;
        RECT 2559.740 550.980 2560.060 551.300 ;
        RECT 2656.340 550.980 2656.660 551.300 ;
      LAYER met4 ;
        RECT 718.815 2358.415 719.145 2358.745 ;
        RECT 718.830 2327.450 719.130 2358.415 ;
        RECT 718.830 2327.150 720.970 2327.450 ;
        RECT 720.670 2307.050 720.970 2327.150 ;
        RECT 720.670 2306.750 724.650 2307.050 ;
        RECT 724.350 2290.050 724.650 2306.750 ;
        RECT 720.670 2289.750 724.650 2290.050 ;
        RECT 719.045 2222.050 719.375 2222.065 ;
        RECT 720.670 2222.050 720.970 2289.750 ;
        RECT 719.045 2221.750 720.970 2222.050 ;
        RECT 719.045 2221.735 719.375 2221.750 ;
        RECT 718.815 2100.015 719.145 2100.345 ;
        RECT 718.830 2089.450 719.130 2100.015 ;
        RECT 718.830 2089.150 720.970 2089.450 ;
        RECT 720.670 2071.770 720.970 2089.150 ;
        RECT 719.750 2071.470 720.970 2071.770 ;
        RECT 719.750 2052.050 720.050 2071.470 ;
        RECT 718.830 2051.750 720.050 2052.050 ;
        RECT 718.830 2040.505 719.130 2051.750 ;
        RECT 714.215 2040.175 714.545 2040.505 ;
        RECT 718.815 2040.175 719.145 2040.505 ;
        RECT 714.230 1964.345 714.530 2040.175 ;
        RECT 712.375 1964.015 712.705 1964.345 ;
        RECT 714.215 1964.015 714.545 1964.345 ;
        RECT 712.390 1904.505 712.690 1964.015 ;
        RECT 717.910 1904.870 723.730 1905.170 ;
        RECT 717.910 1904.505 718.210 1904.870 ;
        RECT 712.375 1904.175 712.705 1904.505 ;
        RECT 717.895 1904.175 718.225 1904.505 ;
        RECT 718.815 1857.570 719.145 1857.585 ;
        RECT 723.430 1857.570 723.730 1904.870 ;
        RECT 718.815 1857.270 723.730 1857.570 ;
        RECT 718.815 1857.255 719.145 1857.270 ;
        RECT 718.815 1817.450 719.145 1817.465 ;
        RECT 718.815 1817.150 720.050 1817.450 ;
        RECT 718.815 1817.135 719.145 1817.150 ;
        RECT 712.375 1783.135 712.705 1783.465 ;
        RECT 718.815 1783.450 719.145 1783.465 ;
        RECT 719.750 1783.450 720.050 1817.150 ;
        RECT 718.815 1783.150 720.050 1783.450 ;
        RECT 718.815 1783.135 719.145 1783.150 ;
        RECT 712.390 1732.465 712.690 1783.135 ;
        RECT 712.375 1732.135 712.705 1732.465 ;
        RECT 714.215 1730.775 714.545 1731.105 ;
        RECT 714.230 1693.705 714.530 1730.775 ;
        RECT 714.215 1693.375 714.545 1693.705 ;
        RECT 717.895 1693.375 718.225 1693.705 ;
        RECT 717.910 1661.745 718.210 1693.375 ;
        RECT 717.895 1661.415 718.225 1661.745 ;
        RECT 718.815 1631.130 719.145 1631.145 ;
        RECT 718.815 1630.830 723.730 1631.130 ;
        RECT 718.815 1630.815 719.145 1630.830 ;
        RECT 723.430 1593.050 723.730 1630.830 ;
        RECT 721.590 1592.750 723.730 1593.050 ;
        RECT 721.590 1576.050 721.890 1592.750 ;
        RECT 721.590 1575.750 727.410 1576.050 ;
        RECT 727.110 1548.850 727.410 1575.750 ;
        RECT 718.830 1548.550 727.410 1548.850 ;
        RECT 718.830 1542.745 719.130 1548.550 ;
        RECT 718.815 1542.415 719.145 1542.745 ;
        RECT 718.815 1518.250 719.145 1518.265 ;
        RECT 718.815 1517.950 725.570 1518.250 ;
        RECT 718.815 1517.935 719.145 1517.950 ;
        RECT 725.270 1501.250 725.570 1517.950 ;
        RECT 722.510 1500.950 725.570 1501.250 ;
        RECT 722.510 1484.250 722.810 1500.950 ;
        RECT 722.510 1483.950 726.490 1484.250 ;
        RECT 726.190 1419.650 726.490 1483.950 ;
        RECT 725.270 1419.350 726.490 1419.650 ;
        RECT 725.270 1386.090 725.570 1419.350 ;
        RECT 724.830 1384.910 726.010 1386.090 ;
        RECT 723.910 1378.110 725.090 1379.290 ;
        RECT 724.350 1355.730 724.650 1378.110 ;
        RECT 724.350 1355.430 725.570 1355.730 ;
        RECT 725.270 1355.050 725.570 1355.430 ;
        RECT 725.270 1354.750 727.410 1355.050 ;
        RECT 727.110 1323.105 727.410 1354.750 ;
        RECT 727.095 1322.775 727.425 1323.105 ;
        RECT 728.935 1179.975 729.265 1180.305 ;
        RECT 728.950 1113.650 729.250 1179.975 ;
        RECT 728.030 1113.350 729.250 1113.650 ;
        RECT 728.030 1055.865 728.330 1113.350 ;
        RECT 726.175 1055.535 726.505 1055.865 ;
        RECT 728.015 1055.535 728.345 1055.865 ;
        RECT 726.190 994.665 726.490 1055.535 ;
        RECT 726.175 994.335 726.505 994.665 ;
        RECT 727.095 993.655 727.425 993.985 ;
        RECT 727.110 879.745 727.410 993.655 ;
        RECT 727.095 879.415 727.425 879.745 ;
        RECT 726.175 878.735 726.505 879.065 ;
        RECT 726.190 800.185 726.490 878.735 ;
        RECT 726.175 799.855 726.505 800.185 ;
        RECT 728.015 799.175 728.345 799.505 ;
        RECT 728.030 729.450 728.330 799.175 ;
        RECT 727.110 729.150 728.330 729.450 ;
        RECT 727.110 678.450 727.410 729.150 ;
        RECT 725.270 678.150 727.410 678.450 ;
        RECT 725.270 631.545 725.570 678.150 ;
        RECT 725.255 631.215 725.585 631.545 ;
        RECT 917.535 555.055 917.865 555.385 ;
        RECT 917.550 553.345 917.850 555.055 ;
        RECT 1544.055 554.375 1544.385 554.705 ;
        RECT 1924.935 554.375 1925.265 554.705 ;
        RECT 917.535 553.015 917.865 553.345 ;
        RECT 1544.070 552.650 1544.370 554.375 ;
        RECT 1924.950 553.345 1925.250 554.375 ;
        RECT 2656.335 553.695 2656.665 554.025 ;
        RECT 1924.935 553.015 1925.265 553.345 ;
        RECT 2173.335 553.015 2173.665 553.345 ;
        RECT 2559.735 553.015 2560.065 553.345 ;
        RECT 1544.975 552.650 1545.305 552.665 ;
        RECT 1544.070 552.350 1545.305 552.650 ;
        RECT 1544.975 552.335 1545.305 552.350 ;
        RECT 2173.350 551.985 2173.650 553.015 ;
        RECT 2173.335 551.655 2173.665 551.985 ;
        RECT 2559.750 551.305 2560.050 553.015 ;
        RECT 2656.350 551.305 2656.650 553.695 ;
        RECT 2559.735 550.975 2560.065 551.305 ;
        RECT 2656.335 550.975 2656.665 551.305 ;
      LAYER met5 ;
        RECT 723.700 1384.700 726.220 1386.300 ;
        RECT 723.700 1377.900 725.300 1384.700 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 13.870 1683.920 14.190 1683.980 ;
        RECT 25.830 1683.920 26.150 1683.980 ;
        RECT 13.870 1683.780 26.150 1683.920 ;
        RECT 13.870 1683.720 14.190 1683.780 ;
        RECT 25.830 1683.720 26.150 1683.780 ;
        RECT 25.830 1320.120 26.150 1320.180 ;
        RECT 1620.190 1320.120 1620.510 1320.180 ;
        RECT 25.830 1319.980 1620.510 1320.120 ;
        RECT 25.830 1319.920 26.150 1319.980 ;
        RECT 1620.190 1319.920 1620.510 1319.980 ;
      LAYER via ;
        RECT 13.900 1683.720 14.160 1683.980 ;
        RECT 25.860 1683.720 26.120 1683.980 ;
        RECT 25.860 1319.920 26.120 1320.180 ;
        RECT 1620.220 1319.920 1620.480 1320.180 ;
      LAYER met2 ;
        RECT 13.890 1687.235 14.170 1687.605 ;
        RECT 13.960 1684.010 14.100 1687.235 ;
        RECT 13.900 1683.690 14.160 1684.010 ;
        RECT 25.860 1683.690 26.120 1684.010 ;
        RECT 25.920 1320.210 26.060 1683.690 ;
        RECT 1620.260 1323.135 1620.540 1327.135 ;
        RECT 1620.280 1320.210 1620.420 1323.135 ;
        RECT 25.860 1319.890 26.120 1320.210 ;
        RECT 1620.220 1319.890 1620.480 1320.210 ;
      LAYER via2 ;
        RECT 13.890 1687.280 14.170 1687.560 ;
      LAYER met3 ;
        RECT -4.800 1687.570 2.400 1688.020 ;
        RECT 13.865 1687.570 14.195 1687.585 ;
        RECT -4.800 1687.270 14.195 1687.570 ;
        RECT -4.800 1686.820 2.400 1687.270 ;
        RECT 13.865 1687.255 14.195 1687.270 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 26.750 2382.620 27.070 2382.680 ;
        RECT 1161.110 2382.620 1161.430 2382.680 ;
        RECT 26.750 2382.480 1161.430 2382.620 ;
        RECT 26.750 2382.420 27.070 2382.480 ;
        RECT 1161.110 2382.420 1161.430 2382.480 ;
        RECT 13.870 1475.500 14.190 1475.560 ;
        RECT 26.750 1475.500 27.070 1475.560 ;
        RECT 13.870 1475.360 27.070 1475.500 ;
        RECT 13.870 1475.300 14.190 1475.360 ;
        RECT 26.750 1475.300 27.070 1475.360 ;
      LAYER via ;
        RECT 26.780 2382.420 27.040 2382.680 ;
        RECT 1161.140 2382.420 1161.400 2382.680 ;
        RECT 13.900 1475.300 14.160 1475.560 ;
        RECT 26.780 1475.300 27.040 1475.560 ;
      LAYER met2 ;
        RECT 26.780 2382.390 27.040 2382.710 ;
        RECT 1161.140 2382.390 1161.400 2382.710 ;
        RECT 26.840 1475.590 26.980 2382.390 ;
        RECT 1161.200 2377.880 1161.340 2382.390 ;
        RECT 1161.180 2373.880 1161.460 2377.880 ;
        RECT 13.900 1475.270 14.160 1475.590 ;
        RECT 26.780 1475.270 27.040 1475.590 ;
        RECT 13.960 1472.045 14.100 1475.270 ;
        RECT 13.890 1471.675 14.170 1472.045 ;
      LAYER via2 ;
        RECT 13.890 1471.720 14.170 1472.000 ;
      LAYER met3 ;
        RECT -4.800 1472.010 2.400 1472.460 ;
        RECT 13.865 1472.010 14.195 1472.025 ;
        RECT -4.800 1471.710 14.195 1472.010 ;
        RECT -4.800 1471.260 2.400 1471.710 ;
        RECT 13.865 1471.695 14.195 1471.710 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 24.910 1401.040 25.230 1401.100 ;
        RECT 706.630 1401.040 706.950 1401.100 ;
        RECT 24.910 1400.900 706.950 1401.040 ;
        RECT 24.910 1400.840 25.230 1400.900 ;
        RECT 706.630 1400.840 706.950 1400.900 ;
        RECT 13.870 1258.920 14.190 1258.980 ;
        RECT 24.910 1258.920 25.230 1258.980 ;
        RECT 13.870 1258.780 25.230 1258.920 ;
        RECT 13.870 1258.720 14.190 1258.780 ;
        RECT 24.910 1258.720 25.230 1258.780 ;
      LAYER via ;
        RECT 24.940 1400.840 25.200 1401.100 ;
        RECT 706.660 1400.840 706.920 1401.100 ;
        RECT 13.900 1258.720 14.160 1258.980 ;
        RECT 24.940 1258.720 25.200 1258.980 ;
      LAYER met2 ;
        RECT 706.650 1403.675 706.930 1404.045 ;
        RECT 706.720 1401.130 706.860 1403.675 ;
        RECT 24.940 1400.810 25.200 1401.130 ;
        RECT 706.660 1400.810 706.920 1401.130 ;
        RECT 25.000 1259.010 25.140 1400.810 ;
        RECT 13.900 1258.690 14.160 1259.010 ;
        RECT 24.940 1258.690 25.200 1259.010 ;
        RECT 13.960 1256.485 14.100 1258.690 ;
        RECT 13.890 1256.115 14.170 1256.485 ;
      LAYER via2 ;
        RECT 706.650 1403.720 706.930 1404.000 ;
        RECT 13.890 1256.160 14.170 1256.440 ;
      LAYER met3 ;
        RECT 706.625 1404.010 706.955 1404.025 ;
        RECT 715.810 1404.010 719.810 1404.015 ;
        RECT 706.625 1403.710 719.810 1404.010 ;
        RECT 706.625 1403.695 706.955 1403.710 ;
        RECT 715.810 1403.415 719.810 1403.710 ;
        RECT -4.800 1256.450 2.400 1256.900 ;
        RECT 13.865 1256.450 14.195 1256.465 ;
        RECT -4.800 1256.150 14.195 1256.450 ;
        RECT -4.800 1255.700 2.400 1256.150 ;
        RECT 13.865 1256.135 14.195 1256.150 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 26.290 2381.940 26.610 2382.000 ;
        RECT 1207.110 2381.940 1207.430 2382.000 ;
        RECT 26.290 2381.800 1207.430 2381.940 ;
        RECT 26.290 2381.740 26.610 2381.800 ;
        RECT 1207.110 2381.740 1207.430 2381.800 ;
        RECT 13.870 1041.320 14.190 1041.380 ;
        RECT 26.290 1041.320 26.610 1041.380 ;
        RECT 13.870 1041.180 26.610 1041.320 ;
        RECT 13.870 1041.120 14.190 1041.180 ;
        RECT 26.290 1041.120 26.610 1041.180 ;
      LAYER via ;
        RECT 26.320 2381.740 26.580 2382.000 ;
        RECT 1207.140 2381.740 1207.400 2382.000 ;
        RECT 13.900 1041.120 14.160 1041.380 ;
        RECT 26.320 1041.120 26.580 1041.380 ;
      LAYER met2 ;
        RECT 26.320 2381.710 26.580 2382.030 ;
        RECT 1207.140 2381.710 1207.400 2382.030 ;
        RECT 26.380 1041.410 26.520 2381.710 ;
        RECT 1207.200 2377.880 1207.340 2381.710 ;
        RECT 1207.180 2373.880 1207.460 2377.880 ;
        RECT 13.900 1041.090 14.160 1041.410 ;
        RECT 26.320 1041.090 26.580 1041.410 ;
        RECT 13.960 1040.925 14.100 1041.090 ;
        RECT 13.890 1040.555 14.170 1040.925 ;
      LAYER via2 ;
        RECT 13.890 1040.600 14.170 1040.880 ;
      LAYER met3 ;
        RECT -4.800 1040.890 2.400 1041.340 ;
        RECT 13.865 1040.890 14.195 1040.905 ;
        RECT -4.800 1040.590 14.195 1040.890 ;
        RECT -4.800 1040.140 2.400 1040.590 ;
        RECT 13.865 1040.575 14.195 1040.590 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 24.450 2382.960 24.770 2383.020 ;
        RECT 1138.110 2382.960 1138.430 2383.020 ;
        RECT 24.450 2382.820 1138.430 2382.960 ;
        RECT 24.450 2382.760 24.770 2382.820 ;
        RECT 1138.110 2382.760 1138.430 2382.820 ;
        RECT 13.870 826.780 14.190 826.840 ;
        RECT 24.450 826.780 24.770 826.840 ;
        RECT 13.870 826.640 24.770 826.780 ;
        RECT 13.870 826.580 14.190 826.640 ;
        RECT 24.450 826.580 24.770 826.640 ;
      LAYER via ;
        RECT 24.480 2382.760 24.740 2383.020 ;
        RECT 1138.140 2382.760 1138.400 2383.020 ;
        RECT 13.900 826.580 14.160 826.840 ;
        RECT 24.480 826.580 24.740 826.840 ;
      LAYER met2 ;
        RECT 24.480 2382.730 24.740 2383.050 ;
        RECT 1138.140 2382.730 1138.400 2383.050 ;
        RECT 24.540 826.870 24.680 2382.730 ;
        RECT 1138.200 2377.880 1138.340 2382.730 ;
        RECT 1138.180 2373.880 1138.460 2377.880 ;
        RECT 13.900 826.550 14.160 826.870 ;
        RECT 24.480 826.550 24.740 826.870 ;
        RECT 13.960 825.365 14.100 826.550 ;
        RECT 13.890 824.995 14.170 825.365 ;
      LAYER via2 ;
        RECT 13.890 825.040 14.170 825.320 ;
      LAYER met3 ;
        RECT -4.800 825.330 2.400 825.780 ;
        RECT 13.865 825.330 14.195 825.345 ;
        RECT -4.800 825.030 14.195 825.330 ;
        RECT -4.800 824.580 2.400 825.030 ;
        RECT 13.865 825.015 14.195 825.030 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.550 613.940 17.870 614.000 ;
        RECT 1187.330 613.940 1187.650 614.000 ;
        RECT 17.550 613.800 1187.650 613.940 ;
        RECT 17.550 613.740 17.870 613.800 ;
        RECT 1187.330 613.740 1187.650 613.800 ;
      LAYER via ;
        RECT 17.580 613.740 17.840 614.000 ;
        RECT 1187.360 613.740 1187.620 614.000 ;
      LAYER met2 ;
        RECT 1192.460 1323.690 1192.740 1327.135 ;
        RECT 1187.420 1323.550 1192.740 1323.690 ;
        RECT 1187.420 614.030 1187.560 1323.550 ;
        RECT 1192.460 1323.135 1192.740 1323.550 ;
        RECT 17.580 613.710 17.840 614.030 ;
        RECT 1187.360 613.710 1187.620 614.030 ;
        RECT 17.640 610.485 17.780 613.710 ;
        RECT 17.570 610.115 17.850 610.485 ;
      LAYER via2 ;
        RECT 17.570 610.160 17.850 610.440 ;
      LAYER met3 ;
        RECT -4.800 610.450 2.400 610.900 ;
        RECT 17.545 610.450 17.875 610.465 ;
        RECT -4.800 610.150 17.875 610.450 ;
        RECT -4.800 609.700 2.400 610.150 ;
        RECT 17.545 610.135 17.875 610.150 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 16.650 399.995 16.930 400.365 ;
        RECT 16.720 394.925 16.860 399.995 ;
        RECT 16.650 394.555 16.930 394.925 ;
      LAYER via2 ;
        RECT 16.650 400.040 16.930 400.320 ;
        RECT 16.650 394.600 16.930 394.880 ;
      LAYER met3 ;
        RECT 1755.835 2177.850 1759.835 2177.855 ;
        RECT 1780.470 2177.850 1780.850 2177.860 ;
        RECT 1755.835 2177.550 1780.850 2177.850 ;
        RECT 1755.835 2177.255 1759.835 2177.550 ;
        RECT 1780.470 2177.540 1780.850 2177.550 ;
        RECT 16.625 400.330 16.955 400.345 ;
        RECT 1780.470 400.330 1780.850 400.340 ;
        RECT 16.625 400.030 1780.850 400.330 ;
        RECT 16.625 400.015 16.955 400.030 ;
        RECT 1780.470 400.020 1780.850 400.030 ;
        RECT -4.800 394.890 2.400 395.340 ;
        RECT 16.625 394.890 16.955 394.905 ;
        RECT -4.800 394.590 16.955 394.890 ;
        RECT -4.800 394.140 2.400 394.590 ;
        RECT 16.625 394.575 16.955 394.590 ;
      LAYER via3 ;
        RECT 1780.500 2177.540 1780.820 2177.860 ;
        RECT 1780.500 400.020 1780.820 400.340 ;
      LAYER met4 ;
        RECT 1780.495 2177.535 1780.825 2177.865 ;
        RECT 1780.510 400.345 1780.810 2177.535 ;
        RECT 1780.495 400.015 1780.825 400.345 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 23.990 2380.580 24.310 2380.640 ;
        RECT 1704.830 2380.580 1705.150 2380.640 ;
        RECT 23.990 2380.440 1705.150 2380.580 ;
        RECT 23.990 2380.380 24.310 2380.440 ;
        RECT 1704.830 2380.380 1705.150 2380.440 ;
        RECT 13.870 179.420 14.190 179.480 ;
        RECT 23.990 179.420 24.310 179.480 ;
        RECT 13.870 179.280 24.310 179.420 ;
        RECT 13.870 179.220 14.190 179.280 ;
        RECT 23.990 179.220 24.310 179.280 ;
      LAYER via ;
        RECT 24.020 2380.380 24.280 2380.640 ;
        RECT 1704.860 2380.380 1705.120 2380.640 ;
        RECT 13.900 179.220 14.160 179.480 ;
        RECT 24.020 179.220 24.280 179.480 ;
      LAYER met2 ;
        RECT 24.020 2380.350 24.280 2380.670 ;
        RECT 1704.860 2380.350 1705.120 2380.670 ;
        RECT 24.080 179.510 24.220 2380.350 ;
        RECT 1704.920 2377.880 1705.060 2380.350 ;
        RECT 1704.900 2373.880 1705.180 2377.880 ;
        RECT 13.900 179.365 14.160 179.510 ;
        RECT 13.890 178.995 14.170 179.365 ;
        RECT 24.020 179.190 24.280 179.510 ;
      LAYER via2 ;
        RECT 13.890 179.040 14.170 179.320 ;
      LAYER met3 ;
        RECT -4.800 179.330 2.400 179.780 ;
        RECT 13.865 179.330 14.195 179.345 ;
        RECT -4.800 179.030 14.195 179.330 ;
        RECT -4.800 178.580 2.400 179.030 ;
        RECT 13.865 179.015 14.195 179.030 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1772.910 1911.380 1773.230 1911.440 ;
        RECT 1777.970 1911.380 1778.290 1911.440 ;
        RECT 1772.910 1911.240 1778.290 1911.380 ;
        RECT 1772.910 1911.180 1773.230 1911.240 ;
        RECT 1777.970 1911.180 1778.290 1911.240 ;
        RECT 1777.970 793.460 1778.290 793.520 ;
        RECT 2900.370 793.460 2900.690 793.520 ;
        RECT 1777.970 793.320 2900.690 793.460 ;
        RECT 1777.970 793.260 1778.290 793.320 ;
        RECT 2900.370 793.260 2900.690 793.320 ;
      LAYER via ;
        RECT 1772.940 1911.180 1773.200 1911.440 ;
        RECT 1778.000 1911.180 1778.260 1911.440 ;
        RECT 1778.000 793.260 1778.260 793.520 ;
        RECT 2900.400 793.260 2900.660 793.520 ;
      LAYER met2 ;
        RECT 1772.930 1912.315 1773.210 1912.685 ;
        RECT 1773.000 1911.470 1773.140 1912.315 ;
        RECT 1772.940 1911.150 1773.200 1911.470 ;
        RECT 1778.000 1911.150 1778.260 1911.470 ;
        RECT 1778.060 793.550 1778.200 1911.150 ;
        RECT 1778.000 793.230 1778.260 793.550 ;
        RECT 2900.400 793.230 2900.660 793.550 ;
        RECT 2900.460 792.045 2900.600 793.230 ;
        RECT 2900.390 791.675 2900.670 792.045 ;
      LAYER via2 ;
        RECT 1772.930 1912.360 1773.210 1912.640 ;
        RECT 2900.390 791.720 2900.670 792.000 ;
      LAYER met3 ;
        RECT 1755.835 1912.650 1759.835 1912.655 ;
        RECT 1772.905 1912.650 1773.235 1912.665 ;
        RECT 1755.835 1912.350 1773.235 1912.650 ;
        RECT 1755.835 1912.055 1759.835 1912.350 ;
        RECT 1772.905 1912.335 1773.235 1912.350 ;
        RECT 2900.365 792.010 2900.695 792.025 ;
        RECT 2917.600 792.010 2924.800 792.460 ;
        RECT 2900.365 791.710 2924.800 792.010 ;
        RECT 2900.365 791.695 2900.695 791.710 ;
        RECT 2917.600 791.260 2924.800 791.710 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1103.610 1028.060 1103.930 1028.120 ;
        RECT 2900.370 1028.060 2900.690 1028.120 ;
        RECT 1103.610 1027.920 2900.690 1028.060 ;
        RECT 1103.610 1027.860 1103.930 1027.920 ;
        RECT 2900.370 1027.860 2900.690 1027.920 ;
      LAYER via ;
        RECT 1103.640 1027.860 1103.900 1028.120 ;
        RECT 2900.400 1027.860 2900.660 1028.120 ;
      LAYER met2 ;
        RECT 1100.460 1323.690 1100.740 1327.135 ;
        RECT 1100.460 1323.550 1103.840 1323.690 ;
        RECT 1100.460 1323.135 1100.740 1323.550 ;
        RECT 1103.700 1028.150 1103.840 1323.550 ;
        RECT 1103.640 1027.830 1103.900 1028.150 ;
        RECT 2900.400 1027.830 2900.660 1028.150 ;
        RECT 2900.460 1026.645 2900.600 1027.830 ;
        RECT 2900.390 1026.275 2900.670 1026.645 ;
      LAYER via2 ;
        RECT 2900.390 1026.320 2900.670 1026.600 ;
      LAYER met3 ;
        RECT 2900.365 1026.610 2900.695 1026.625 ;
        RECT 2917.600 1026.610 2924.800 1027.060 ;
        RECT 2900.365 1026.310 2924.800 1026.610 ;
        RECT 2900.365 1026.295 2900.695 1026.310 ;
        RECT 2917.600 1025.860 2924.800 1026.310 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 868.550 1262.660 868.870 1262.720 ;
        RECT 2900.370 1262.660 2900.690 1262.720 ;
        RECT 868.550 1262.520 2900.690 1262.660 ;
        RECT 868.550 1262.460 868.870 1262.520 ;
        RECT 2900.370 1262.460 2900.690 1262.520 ;
      LAYER via ;
        RECT 868.580 1262.460 868.840 1262.720 ;
        RECT 2900.400 1262.460 2900.660 1262.720 ;
      LAYER met2 ;
        RECT 868.620 1323.135 868.900 1327.135 ;
        RECT 868.640 1262.750 868.780 1323.135 ;
        RECT 868.580 1262.430 868.840 1262.750 ;
        RECT 2900.400 1262.430 2900.660 1262.750 ;
        RECT 2900.460 1261.245 2900.600 1262.430 ;
        RECT 2900.390 1260.875 2900.670 1261.245 ;
      LAYER via2 ;
        RECT 2900.390 1260.920 2900.670 1261.200 ;
      LAYER met3 ;
        RECT 2900.365 1261.210 2900.695 1261.225 ;
        RECT 2917.600 1261.210 2924.800 1261.660 ;
        RECT 2900.365 1260.910 2924.800 1261.210 ;
        RECT 2900.365 1260.895 2900.695 1260.910 ;
        RECT 2917.600 1260.460 2924.800 1260.910 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1754.585 2242.725 1754.755 2296.615 ;
        RECT 1754.585 2214.845 1754.755 2240.175 ;
        RECT 1754.585 1994.525 1754.755 2048.415 ;
      LAYER mcon ;
        RECT 1754.585 2296.445 1754.755 2296.615 ;
        RECT 1754.585 2240.005 1754.755 2240.175 ;
        RECT 1754.585 2048.245 1754.755 2048.415 ;
      LAYER met1 ;
        RECT 1754.510 2342.500 1754.830 2342.560 ;
        RECT 1756.350 2342.500 1756.670 2342.560 ;
        RECT 1754.510 2342.360 1756.670 2342.500 ;
        RECT 1754.510 2342.300 1754.830 2342.360 ;
        RECT 1756.350 2342.300 1756.670 2342.360 ;
        RECT 1754.510 2320.200 1754.830 2320.460 ;
        RECT 1754.600 2319.780 1754.740 2320.200 ;
        RECT 1754.510 2319.520 1754.830 2319.780 ;
        RECT 1754.510 2296.600 1754.830 2296.660 ;
        RECT 1754.315 2296.460 1754.830 2296.600 ;
        RECT 1754.510 2296.400 1754.830 2296.460 ;
        RECT 1754.510 2242.880 1754.830 2242.940 ;
        RECT 1754.315 2242.740 1754.830 2242.880 ;
        RECT 1754.510 2242.680 1754.830 2242.740 ;
        RECT 1754.510 2240.160 1754.830 2240.220 ;
        RECT 1754.315 2240.020 1754.830 2240.160 ;
        RECT 1754.510 2239.960 1754.830 2240.020 ;
        RECT 1754.510 2215.000 1754.830 2215.060 ;
        RECT 1754.315 2214.860 1754.830 2215.000 ;
        RECT 1754.510 2214.800 1754.830 2214.860 ;
        RECT 1754.510 2048.400 1754.830 2048.460 ;
        RECT 1754.315 2048.260 1754.830 2048.400 ;
        RECT 1754.510 2048.200 1754.830 2048.260 ;
        RECT 1754.510 1994.680 1754.830 1994.740 ;
        RECT 1754.315 1994.540 1754.830 1994.680 ;
        RECT 1754.510 1994.480 1754.830 1994.540 ;
        RECT 1754.970 1845.420 1755.290 1845.480 ;
        RECT 1779.810 1845.420 1780.130 1845.480 ;
        RECT 1754.970 1845.280 1780.130 1845.420 ;
        RECT 1754.970 1845.220 1755.290 1845.280 ;
        RECT 1779.810 1845.220 1780.130 1845.280 ;
        RECT 1779.810 1497.260 1780.130 1497.320 ;
        RECT 2900.830 1497.260 2901.150 1497.320 ;
        RECT 1779.810 1497.120 2901.150 1497.260 ;
        RECT 1779.810 1497.060 1780.130 1497.120 ;
        RECT 2900.830 1497.060 2901.150 1497.120 ;
      LAYER via ;
        RECT 1754.540 2342.300 1754.800 2342.560 ;
        RECT 1756.380 2342.300 1756.640 2342.560 ;
        RECT 1754.540 2320.200 1754.800 2320.460 ;
        RECT 1754.540 2319.520 1754.800 2319.780 ;
        RECT 1754.540 2296.400 1754.800 2296.660 ;
        RECT 1754.540 2242.680 1754.800 2242.940 ;
        RECT 1754.540 2239.960 1754.800 2240.220 ;
        RECT 1754.540 2214.800 1754.800 2215.060 ;
        RECT 1754.540 2048.200 1754.800 2048.460 ;
        RECT 1754.540 1994.480 1754.800 1994.740 ;
        RECT 1755.000 1845.220 1755.260 1845.480 ;
        RECT 1779.840 1845.220 1780.100 1845.480 ;
        RECT 1779.840 1497.060 1780.100 1497.320 ;
        RECT 2900.860 1497.060 2901.120 1497.320 ;
      LAYER met2 ;
        RECT 1756.420 2373.880 1756.700 2377.880 ;
        RECT 1756.440 2342.590 1756.580 2373.880 ;
        RECT 1754.540 2342.270 1754.800 2342.590 ;
        RECT 1756.380 2342.270 1756.640 2342.590 ;
        RECT 1754.600 2320.490 1754.740 2342.270 ;
        RECT 1754.540 2320.170 1754.800 2320.490 ;
        RECT 1754.540 2319.490 1754.800 2319.810 ;
        RECT 1754.600 2296.690 1754.740 2319.490 ;
        RECT 1754.540 2296.370 1754.800 2296.690 ;
        RECT 1754.540 2242.650 1754.800 2242.970 ;
        RECT 1754.600 2240.250 1754.740 2242.650 ;
        RECT 1754.540 2239.930 1754.800 2240.250 ;
        RECT 1754.540 2214.770 1754.800 2215.090 ;
        RECT 1754.600 2048.490 1754.740 2214.770 ;
        RECT 1754.540 2048.170 1754.800 2048.490 ;
        RECT 1754.540 1994.450 1754.800 1994.770 ;
        RECT 1754.600 1873.130 1754.740 1994.450 ;
        RECT 1754.600 1872.990 1755.200 1873.130 ;
        RECT 1755.060 1845.510 1755.200 1872.990 ;
        RECT 1755.000 1845.190 1755.260 1845.510 ;
        RECT 1779.840 1845.190 1780.100 1845.510 ;
        RECT 1779.900 1497.350 1780.040 1845.190 ;
        RECT 1779.840 1497.030 1780.100 1497.350 ;
        RECT 2900.860 1497.030 2901.120 1497.350 ;
        RECT 2900.920 1495.845 2901.060 1497.030 ;
        RECT 2900.850 1495.475 2901.130 1495.845 ;
      LAYER via2 ;
        RECT 2900.850 1495.520 2901.130 1495.800 ;
      LAYER met3 ;
        RECT 2900.825 1495.810 2901.155 1495.825 ;
        RECT 2917.600 1495.810 2924.800 1496.260 ;
        RECT 2900.825 1495.510 2924.800 1495.810 ;
        RECT 2900.825 1495.495 2901.155 1495.510 ;
        RECT 2917.600 1495.060 2924.800 1495.510 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1311.070 2387.380 1311.390 2387.440 ;
        RECT 1778.890 2387.380 1779.210 2387.440 ;
        RECT 1311.070 2387.240 1779.210 2387.380 ;
        RECT 1311.070 2387.180 1311.390 2387.240 ;
        RECT 1778.890 2387.180 1779.210 2387.240 ;
        RECT 1778.890 1731.860 1779.210 1731.920 ;
        RECT 2900.830 1731.860 2901.150 1731.920 ;
        RECT 1778.890 1731.720 2901.150 1731.860 ;
        RECT 1778.890 1731.660 1779.210 1731.720 ;
        RECT 2900.830 1731.660 2901.150 1731.720 ;
      LAYER via ;
        RECT 1311.100 2387.180 1311.360 2387.440 ;
        RECT 1778.920 2387.180 1779.180 2387.440 ;
        RECT 1778.920 1731.660 1779.180 1731.920 ;
        RECT 2900.860 1731.660 2901.120 1731.920 ;
      LAYER met2 ;
        RECT 1311.100 2387.150 1311.360 2387.470 ;
        RECT 1778.920 2387.150 1779.180 2387.470 ;
        RECT 1311.160 2377.880 1311.300 2387.150 ;
        RECT 1311.140 2373.880 1311.420 2377.880 ;
        RECT 1778.980 1731.950 1779.120 2387.150 ;
        RECT 1778.920 1731.630 1779.180 1731.950 ;
        RECT 2900.860 1731.630 2901.120 1731.950 ;
        RECT 2900.920 1730.445 2901.060 1731.630 ;
        RECT 2900.850 1730.075 2901.130 1730.445 ;
      LAYER via2 ;
        RECT 2900.850 1730.120 2901.130 1730.400 ;
      LAYER met3 ;
        RECT 2900.825 1730.410 2901.155 1730.425 ;
        RECT 2917.600 1730.410 2924.800 1730.860 ;
        RECT 2900.825 1730.110 2924.800 1730.410 ;
        RECT 2900.825 1730.095 2901.155 1730.110 ;
        RECT 2917.600 1729.660 2924.800 1730.110 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 837.270 2383.980 837.590 2384.040 ;
        RECT 1777.970 2383.980 1778.290 2384.040 ;
        RECT 837.270 2383.840 1778.290 2383.980 ;
        RECT 837.270 2383.780 837.590 2383.840 ;
        RECT 1777.970 2383.780 1778.290 2383.840 ;
        RECT 1777.970 1966.460 1778.290 1966.520 ;
        RECT 2900.830 1966.460 2901.150 1966.520 ;
        RECT 1777.970 1966.320 2901.150 1966.460 ;
        RECT 1777.970 1966.260 1778.290 1966.320 ;
        RECT 2900.830 1966.260 2901.150 1966.320 ;
      LAYER via ;
        RECT 837.300 2383.780 837.560 2384.040 ;
        RECT 1778.000 2383.780 1778.260 2384.040 ;
        RECT 1778.000 1966.260 1778.260 1966.520 ;
        RECT 2900.860 1966.260 2901.120 1966.520 ;
      LAYER met2 ;
        RECT 837.300 2383.750 837.560 2384.070 ;
        RECT 1778.000 2383.750 1778.260 2384.070 ;
        RECT 837.360 2377.880 837.500 2383.750 ;
        RECT 837.340 2373.880 837.620 2377.880 ;
        RECT 1778.060 1966.550 1778.200 2383.750 ;
        RECT 1778.000 1966.230 1778.260 1966.550 ;
        RECT 2900.860 1966.230 2901.120 1966.550 ;
        RECT 2900.920 1965.045 2901.060 1966.230 ;
        RECT 2900.850 1964.675 2901.130 1965.045 ;
      LAYER via2 ;
        RECT 2900.850 1964.720 2901.130 1965.000 ;
      LAYER met3 ;
        RECT 2900.825 1965.010 2901.155 1965.025 ;
        RECT 2917.600 1965.010 2924.800 1965.460 ;
        RECT 2900.825 1964.710 2924.800 1965.010 ;
        RECT 2900.825 1964.695 2901.155 1964.710 ;
        RECT 2917.600 1964.260 2924.800 1964.710 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 964.230 2384.660 964.550 2384.720 ;
        RECT 1762.790 2384.660 1763.110 2384.720 ;
        RECT 964.230 2384.520 1763.110 2384.660 ;
        RECT 964.230 2384.460 964.550 2384.520 ;
        RECT 1762.790 2384.460 1763.110 2384.520 ;
        RECT 1762.790 2201.060 1763.110 2201.120 ;
        RECT 2898.530 2201.060 2898.850 2201.120 ;
        RECT 1762.790 2200.920 2898.850 2201.060 ;
        RECT 1762.790 2200.860 1763.110 2200.920 ;
        RECT 2898.530 2200.860 2898.850 2200.920 ;
      LAYER via ;
        RECT 964.260 2384.460 964.520 2384.720 ;
        RECT 1762.820 2384.460 1763.080 2384.720 ;
        RECT 1762.820 2200.860 1763.080 2201.120 ;
        RECT 2898.560 2200.860 2898.820 2201.120 ;
      LAYER met2 ;
        RECT 964.260 2384.430 964.520 2384.750 ;
        RECT 1762.820 2384.430 1763.080 2384.750 ;
        RECT 964.320 2377.880 964.460 2384.430 ;
        RECT 964.300 2373.880 964.580 2377.880 ;
        RECT 1762.880 2201.150 1763.020 2384.430 ;
        RECT 1762.820 2200.830 1763.080 2201.150 ;
        RECT 2898.560 2200.830 2898.820 2201.150 ;
        RECT 2898.620 2199.645 2898.760 2200.830 ;
        RECT 2898.550 2199.275 2898.830 2199.645 ;
      LAYER via2 ;
        RECT 2898.550 2199.320 2898.830 2199.600 ;
      LAYER met3 ;
        RECT 2898.525 2199.610 2898.855 2199.625 ;
        RECT 2917.600 2199.610 2924.800 2200.060 ;
        RECT 2898.525 2199.310 2924.800 2199.610 ;
        RECT 2898.525 2199.295 2898.855 2199.310 ;
        RECT 2917.600 2198.860 2924.800 2199.310 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1772.910 1900.500 1773.230 1900.560 ;
        RECT 1791.310 1900.500 1791.630 1900.560 ;
        RECT 1772.910 1900.360 1791.630 1900.500 ;
        RECT 1772.910 1900.300 1773.230 1900.360 ;
        RECT 1791.310 1900.300 1791.630 1900.360 ;
        RECT 1791.310 206.960 1791.630 207.020 ;
        RECT 2900.830 206.960 2901.150 207.020 ;
        RECT 1791.310 206.820 2901.150 206.960 ;
        RECT 1791.310 206.760 1791.630 206.820 ;
        RECT 2900.830 206.760 2901.150 206.820 ;
      LAYER via ;
        RECT 1772.940 1900.300 1773.200 1900.560 ;
        RECT 1791.340 1900.300 1791.600 1900.560 ;
        RECT 1791.340 206.760 1791.600 207.020 ;
        RECT 2900.860 206.760 2901.120 207.020 ;
      LAYER met2 ;
        RECT 1772.930 1904.155 1773.210 1904.525 ;
        RECT 1773.000 1900.590 1773.140 1904.155 ;
        RECT 1772.940 1900.270 1773.200 1900.590 ;
        RECT 1791.340 1900.270 1791.600 1900.590 ;
        RECT 1791.400 207.050 1791.540 1900.270 ;
        RECT 1791.340 206.730 1791.600 207.050 ;
        RECT 2900.860 206.730 2901.120 207.050 ;
        RECT 2900.920 205.205 2901.060 206.730 ;
        RECT 2900.850 204.835 2901.130 205.205 ;
      LAYER via2 ;
        RECT 1772.930 1904.200 1773.210 1904.480 ;
        RECT 2900.850 204.880 2901.130 205.160 ;
      LAYER met3 ;
        RECT 1755.835 1904.490 1759.835 1904.495 ;
        RECT 1772.905 1904.490 1773.235 1904.505 ;
        RECT 1755.835 1904.190 1773.235 1904.490 ;
        RECT 1755.835 1903.895 1759.835 1904.190 ;
        RECT 1772.905 1904.175 1773.235 1904.190 ;
        RECT 2900.825 205.170 2901.155 205.185 ;
        RECT 2917.600 205.170 2924.800 205.620 ;
        RECT 2900.825 204.870 2924.800 205.170 ;
        RECT 2900.825 204.855 2901.155 204.870 ;
        RECT 2917.600 204.420 2924.800 204.870 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1770.150 2546.500 1770.470 2546.560 ;
        RECT 2898.990 2546.500 2899.310 2546.560 ;
        RECT 1770.150 2546.360 2899.310 2546.500 ;
        RECT 1770.150 2546.300 1770.470 2546.360 ;
        RECT 2898.990 2546.300 2899.310 2546.360 ;
      LAYER via ;
        RECT 1770.180 2546.300 1770.440 2546.560 ;
        RECT 2899.020 2546.300 2899.280 2546.560 ;
      LAYER met2 ;
        RECT 2899.010 2551.515 2899.290 2551.885 ;
        RECT 2899.080 2546.590 2899.220 2551.515 ;
        RECT 1770.180 2546.270 1770.440 2546.590 ;
        RECT 2899.020 2546.270 2899.280 2546.590 ;
        RECT 1770.240 2271.725 1770.380 2546.270 ;
        RECT 1770.170 2271.355 1770.450 2271.725 ;
      LAYER via2 ;
        RECT 2899.010 2551.560 2899.290 2551.840 ;
        RECT 1770.170 2271.400 1770.450 2271.680 ;
      LAYER met3 ;
        RECT 2898.985 2551.850 2899.315 2551.865 ;
        RECT 2917.600 2551.850 2924.800 2552.300 ;
        RECT 2898.985 2551.550 2924.800 2551.850 ;
        RECT 2898.985 2551.535 2899.315 2551.550 ;
        RECT 2917.600 2551.100 2924.800 2551.550 ;
        RECT 1755.835 2271.690 1759.835 2271.695 ;
        RECT 1770.145 2271.690 1770.475 2271.705 ;
        RECT 1755.835 2271.390 1770.475 2271.690 ;
        RECT 1755.835 2271.095 1759.835 2271.390 ;
        RECT 1770.145 2271.375 1770.475 2271.390 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1777.510 2781.100 1777.830 2781.160 ;
        RECT 2900.830 2781.100 2901.150 2781.160 ;
        RECT 1777.510 2780.960 2901.150 2781.100 ;
        RECT 1777.510 2780.900 1777.830 2780.960 ;
        RECT 2900.830 2780.900 2901.150 2780.960 ;
        RECT 1767.390 1784.900 1767.710 1784.960 ;
        RECT 1777.510 1784.900 1777.830 1784.960 ;
        RECT 1767.390 1784.760 1777.830 1784.900 ;
        RECT 1767.390 1784.700 1767.710 1784.760 ;
        RECT 1777.510 1784.700 1777.830 1784.760 ;
      LAYER via ;
        RECT 1777.540 2780.900 1777.800 2781.160 ;
        RECT 2900.860 2780.900 2901.120 2781.160 ;
        RECT 1767.420 1784.700 1767.680 1784.960 ;
        RECT 1777.540 1784.700 1777.800 1784.960 ;
      LAYER met2 ;
        RECT 2900.850 2786.115 2901.130 2786.485 ;
        RECT 2900.920 2781.190 2901.060 2786.115 ;
        RECT 1777.540 2780.870 1777.800 2781.190 ;
        RECT 2900.860 2780.870 2901.120 2781.190 ;
        RECT 1777.600 1784.990 1777.740 2780.870 ;
        RECT 1767.420 1784.845 1767.680 1784.990 ;
        RECT 1767.410 1784.475 1767.690 1784.845 ;
        RECT 1777.540 1784.670 1777.800 1784.990 ;
      LAYER via2 ;
        RECT 2900.850 2786.160 2901.130 2786.440 ;
        RECT 1767.410 1784.520 1767.690 1784.800 ;
      LAYER met3 ;
        RECT 2900.825 2786.450 2901.155 2786.465 ;
        RECT 2917.600 2786.450 2924.800 2786.900 ;
        RECT 2900.825 2786.150 2924.800 2786.450 ;
        RECT 2900.825 2786.135 2901.155 2786.150 ;
        RECT 2917.600 2785.700 2924.800 2786.150 ;
        RECT 1755.835 1784.810 1759.835 1784.815 ;
        RECT 1767.385 1784.810 1767.715 1784.825 ;
        RECT 1755.835 1784.510 1767.715 1784.810 ;
        RECT 1755.835 1784.215 1759.835 1784.510 ;
        RECT 1767.385 1784.495 1767.715 1784.510 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 712.610 3015.700 712.930 3015.760 ;
        RECT 2900.830 3015.700 2901.150 3015.760 ;
        RECT 712.610 3015.560 2901.150 3015.700 ;
        RECT 712.610 3015.500 712.930 3015.560 ;
        RECT 2900.830 3015.500 2901.150 3015.560 ;
      LAYER via ;
        RECT 712.640 3015.500 712.900 3015.760 ;
        RECT 2900.860 3015.500 2901.120 3015.760 ;
      LAYER met2 ;
        RECT 2900.850 3020.715 2901.130 3021.085 ;
        RECT 2900.920 3015.790 2901.060 3020.715 ;
        RECT 712.640 3015.470 712.900 3015.790 ;
        RECT 2900.860 3015.470 2901.120 3015.790 ;
        RECT 712.700 1601.245 712.840 3015.470 ;
        RECT 712.630 1600.875 712.910 1601.245 ;
      LAYER via2 ;
        RECT 2900.850 3020.760 2901.130 3021.040 ;
        RECT 712.630 1600.920 712.910 1601.200 ;
      LAYER met3 ;
        RECT 2900.825 3021.050 2901.155 3021.065 ;
        RECT 2917.600 3021.050 2924.800 3021.500 ;
        RECT 2900.825 3020.750 2924.800 3021.050 ;
        RECT 2900.825 3020.735 2901.155 3020.750 ;
        RECT 2917.600 3020.300 2924.800 3020.750 ;
        RECT 712.605 1601.210 712.935 1601.225 ;
        RECT 715.810 1601.210 719.810 1601.215 ;
        RECT 712.605 1600.910 719.810 1601.210 ;
        RECT 712.605 1600.895 712.935 1600.910 ;
        RECT 715.810 1600.615 719.810 1600.910 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 979.410 3250.300 979.730 3250.360 ;
        RECT 2900.830 3250.300 2901.150 3250.360 ;
        RECT 979.410 3250.160 2901.150 3250.300 ;
        RECT 979.410 3250.100 979.730 3250.160 ;
        RECT 2900.830 3250.100 2901.150 3250.160 ;
      LAYER via ;
        RECT 979.440 3250.100 979.700 3250.360 ;
        RECT 2900.860 3250.100 2901.120 3250.360 ;
      LAYER met2 ;
        RECT 2900.850 3255.315 2901.130 3255.685 ;
        RECT 2900.920 3250.390 2901.060 3255.315 ;
        RECT 979.440 3250.070 979.700 3250.390 ;
        RECT 2900.860 3250.070 2901.120 3250.390 ;
        RECT 976.260 2377.010 976.540 2377.880 ;
        RECT 979.500 2377.010 979.640 3250.070 ;
        RECT 976.260 2376.870 979.640 2377.010 ;
        RECT 976.260 2373.880 976.540 2376.870 ;
      LAYER via2 ;
        RECT 2900.850 3255.360 2901.130 3255.640 ;
      LAYER met3 ;
        RECT 2900.825 3255.650 2901.155 3255.665 ;
        RECT 2917.600 3255.650 2924.800 3256.100 ;
        RECT 2900.825 3255.350 2924.800 3255.650 ;
        RECT 2900.825 3255.335 2901.155 3255.350 ;
        RECT 2917.600 3254.900 2924.800 3255.350 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2415.070 3486.260 2415.390 3486.320 ;
        RECT 2435.310 3486.260 2435.630 3486.320 ;
        RECT 2415.070 3486.120 2435.630 3486.260 ;
        RECT 2415.070 3486.060 2415.390 3486.120 ;
        RECT 2435.310 3486.060 2435.630 3486.120 ;
      LAYER via ;
        RECT 2415.100 3486.060 2415.360 3486.320 ;
        RECT 2435.340 3486.060 2435.600 3486.320 ;
      LAYER met2 ;
        RECT 2415.100 3486.205 2415.360 3486.350 ;
        RECT 2415.090 3485.835 2415.370 3486.205 ;
        RECT 2435.340 3486.030 2435.600 3486.350 ;
        RECT 2435.400 3484.845 2435.540 3486.030 ;
        RECT 2435.330 3484.475 2435.610 3484.845 ;
        RECT 903.580 1323.135 903.860 1327.135 ;
        RECT 903.600 1319.725 903.740 1323.135 ;
        RECT 903.530 1319.355 903.810 1319.725 ;
      LAYER via2 ;
        RECT 2415.090 3485.880 2415.370 3486.160 ;
        RECT 2435.330 3484.520 2435.610 3484.800 ;
        RECT 903.530 1319.400 903.810 1319.680 ;
      LAYER met3 ;
        RECT 2917.600 3490.250 2924.800 3490.700 ;
        RECT 2916.710 3489.950 2924.800 3490.250 ;
        RECT 2415.065 3486.170 2415.395 3486.185 ;
        RECT 1918.510 3485.870 1966.650 3486.170 ;
        RECT 1778.630 3484.810 1779.010 3484.820 ;
        RECT 1918.510 3484.810 1918.810 3485.870 ;
        RECT 1966.350 3485.490 1966.650 3485.870 ;
        RECT 2015.110 3485.870 2063.250 3486.170 ;
        RECT 1966.350 3485.190 2014.490 3485.490 ;
        RECT 1778.630 3484.510 1918.810 3484.810 ;
        RECT 2014.190 3484.810 2014.490 3485.190 ;
        RECT 2015.110 3484.810 2015.410 3485.870 ;
        RECT 2062.950 3485.490 2063.250 3485.870 ;
        RECT 2111.710 3485.870 2159.850 3486.170 ;
        RECT 2062.950 3485.190 2111.090 3485.490 ;
        RECT 2014.190 3484.510 2015.410 3484.810 ;
        RECT 2110.790 3484.810 2111.090 3485.190 ;
        RECT 2111.710 3484.810 2112.010 3485.870 ;
        RECT 2159.550 3485.490 2159.850 3485.870 ;
        RECT 2208.310 3485.870 2256.450 3486.170 ;
        RECT 2159.550 3485.190 2207.690 3485.490 ;
        RECT 2110.790 3484.510 2112.010 3484.810 ;
        RECT 2207.390 3484.810 2207.690 3485.190 ;
        RECT 2208.310 3484.810 2208.610 3485.870 ;
        RECT 2256.150 3485.490 2256.450 3485.870 ;
        RECT 2304.910 3485.870 2353.050 3486.170 ;
        RECT 2256.150 3485.190 2304.290 3485.490 ;
        RECT 2207.390 3484.510 2208.610 3484.810 ;
        RECT 2303.990 3484.810 2304.290 3485.190 ;
        RECT 2304.910 3484.810 2305.210 3485.870 ;
        RECT 2352.750 3485.490 2353.050 3485.870 ;
        RECT 2401.510 3485.870 2415.395 3486.170 ;
        RECT 2352.750 3485.190 2400.890 3485.490 ;
        RECT 2303.990 3484.510 2305.210 3484.810 ;
        RECT 2400.590 3484.810 2400.890 3485.190 ;
        RECT 2401.510 3484.810 2401.810 3485.870 ;
        RECT 2415.065 3485.855 2415.395 3485.870 ;
        RECT 2463.110 3486.170 2463.490 3486.180 ;
        RECT 2463.110 3485.870 2546.250 3486.170 ;
        RECT 2463.110 3485.860 2463.490 3485.870 ;
        RECT 2545.950 3485.490 2546.250 3485.870 ;
        RECT 2594.710 3485.870 2642.850 3486.170 ;
        RECT 2545.950 3485.190 2594.090 3485.490 ;
        RECT 2400.590 3484.510 2401.810 3484.810 ;
        RECT 2435.305 3484.810 2435.635 3484.825 ;
        RECT 2463.110 3484.810 2463.490 3484.820 ;
        RECT 2435.305 3484.510 2463.490 3484.810 ;
        RECT 2593.790 3484.810 2594.090 3485.190 ;
        RECT 2594.710 3484.810 2595.010 3485.870 ;
        RECT 2642.550 3485.490 2642.850 3485.870 ;
        RECT 2691.310 3485.870 2739.450 3486.170 ;
        RECT 2642.550 3485.190 2690.690 3485.490 ;
        RECT 2593.790 3484.510 2595.010 3484.810 ;
        RECT 2690.390 3484.810 2690.690 3485.190 ;
        RECT 2691.310 3484.810 2691.610 3485.870 ;
        RECT 2739.150 3485.490 2739.450 3485.870 ;
        RECT 2787.910 3485.870 2836.050 3486.170 ;
        RECT 2739.150 3485.190 2787.290 3485.490 ;
        RECT 2690.390 3484.510 2691.610 3484.810 ;
        RECT 2786.990 3484.810 2787.290 3485.190 ;
        RECT 2787.910 3484.810 2788.210 3485.870 ;
        RECT 2835.750 3485.490 2836.050 3485.870 ;
        RECT 2916.710 3485.490 2917.010 3489.950 ;
        RECT 2917.600 3489.500 2924.800 3489.950 ;
        RECT 2835.750 3485.190 2883.890 3485.490 ;
        RECT 2786.990 3484.510 2788.210 3484.810 ;
        RECT 2883.590 3484.810 2883.890 3485.190 ;
        RECT 2884.510 3485.190 2917.010 3485.490 ;
        RECT 2884.510 3484.810 2884.810 3485.190 ;
        RECT 2883.590 3484.510 2884.810 3484.810 ;
        RECT 1778.630 3484.500 1779.010 3484.510 ;
        RECT 2435.305 3484.495 2435.635 3484.510 ;
        RECT 2463.110 3484.500 2463.490 3484.510 ;
        RECT 1778.630 1396.530 1779.010 1396.540 ;
        RECT 1778.630 1396.230 1779.890 1396.530 ;
        RECT 1778.630 1396.220 1779.010 1396.230 ;
        RECT 1778.630 1394.490 1779.010 1394.500 ;
        RECT 1779.590 1394.490 1779.890 1396.230 ;
        RECT 1778.630 1394.190 1779.890 1394.490 ;
        RECT 1778.630 1394.180 1779.010 1394.190 ;
        RECT 903.505 1319.690 903.835 1319.705 ;
        RECT 1778.630 1319.690 1779.010 1319.700 ;
        RECT 903.505 1319.390 1779.010 1319.690 ;
        RECT 903.505 1319.375 903.835 1319.390 ;
        RECT 1778.630 1319.380 1779.010 1319.390 ;
      LAYER via3 ;
        RECT 1778.660 3484.500 1778.980 3484.820 ;
        RECT 2463.140 3485.860 2463.460 3486.180 ;
        RECT 2463.140 3484.500 2463.460 3484.820 ;
        RECT 1778.660 1396.220 1778.980 1396.540 ;
        RECT 1778.660 1394.180 1778.980 1394.500 ;
        RECT 1778.660 1319.380 1778.980 1319.700 ;
      LAYER met4 ;
        RECT 2463.135 3485.855 2463.465 3486.185 ;
        RECT 2463.150 3484.825 2463.450 3485.855 ;
        RECT 1778.655 3484.495 1778.985 3484.825 ;
        RECT 2463.135 3484.495 2463.465 3484.825 ;
        RECT 1778.670 1396.545 1778.970 3484.495 ;
        RECT 1778.655 1396.215 1778.985 1396.545 ;
        RECT 1778.655 1394.175 1778.985 1394.505 ;
        RECT 1778.670 1319.705 1778.970 1394.175 ;
        RECT 1778.655 1319.375 1778.985 1319.705 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1768.310 1400.700 1768.630 1400.760 ;
        RECT 2635.870 1400.700 2636.190 1400.760 ;
        RECT 1768.310 1400.560 2636.190 1400.700 ;
        RECT 1768.310 1400.500 1768.630 1400.560 ;
        RECT 2635.870 1400.500 2636.190 1400.560 ;
      LAYER via ;
        RECT 1768.340 1400.500 1768.600 1400.760 ;
        RECT 2635.900 1400.500 2636.160 1400.760 ;
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
        RECT 2635.960 1400.790 2636.100 3517.600 ;
        RECT 1768.340 1400.470 1768.600 1400.790 ;
        RECT 2635.900 1400.470 2636.160 1400.790 ;
        RECT 1768.400 1399.965 1768.540 1400.470 ;
        RECT 1768.330 1399.595 1768.610 1399.965 ;
      LAYER via2 ;
        RECT 1768.330 1399.640 1768.610 1399.920 ;
      LAYER met3 ;
        RECT 1755.835 1399.930 1759.835 1399.935 ;
        RECT 1768.305 1399.930 1768.635 1399.945 ;
        RECT 1755.835 1399.630 1768.635 1399.930 ;
        RECT 1755.835 1399.335 1759.835 1399.630 ;
        RECT 1768.305 1399.615 1768.635 1399.630 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 711.690 3502.240 712.010 3502.300 ;
        RECT 2311.570 3502.240 2311.890 3502.300 ;
        RECT 711.690 3502.100 2311.890 3502.240 ;
        RECT 711.690 3502.040 712.010 3502.100 ;
        RECT 2311.570 3502.040 2311.890 3502.100 ;
      LAYER via ;
        RECT 711.720 3502.040 711.980 3502.300 ;
        RECT 2311.600 3502.040 2311.860 3502.300 ;
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
        RECT 2311.660 3502.330 2311.800 3517.600 ;
        RECT 711.720 3502.010 711.980 3502.330 ;
        RECT 2311.600 3502.010 2311.860 3502.330 ;
        RECT 711.780 1541.405 711.920 3502.010 ;
        RECT 711.710 1541.035 711.990 1541.405 ;
      LAYER via2 ;
        RECT 711.710 1541.080 711.990 1541.360 ;
      LAYER met3 ;
        RECT 711.685 1541.370 712.015 1541.385 ;
        RECT 715.810 1541.370 719.810 1541.375 ;
        RECT 711.685 1541.070 719.810 1541.370 ;
        RECT 711.685 1541.055 712.015 1541.070 ;
        RECT 715.810 1540.775 719.810 1541.070 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1790.390 3502.920 1790.710 3502.980 ;
        RECT 1987.270 3502.920 1987.590 3502.980 ;
        RECT 1790.390 3502.780 1987.590 3502.920 ;
        RECT 1790.390 3502.720 1790.710 3502.780 ;
        RECT 1987.270 3502.720 1987.590 3502.780 ;
        RECT 1772.910 1771.980 1773.230 1772.040 ;
        RECT 1790.390 1771.980 1790.710 1772.040 ;
        RECT 1772.910 1771.840 1790.710 1771.980 ;
        RECT 1772.910 1771.780 1773.230 1771.840 ;
        RECT 1790.390 1771.780 1790.710 1771.840 ;
      LAYER via ;
        RECT 1790.420 3502.720 1790.680 3502.980 ;
        RECT 1987.300 3502.720 1987.560 3502.980 ;
        RECT 1772.940 1771.780 1773.200 1772.040 ;
        RECT 1790.420 1771.780 1790.680 1772.040 ;
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
        RECT 1987.360 3503.010 1987.500 3517.600 ;
        RECT 1790.420 3502.690 1790.680 3503.010 ;
        RECT 1987.300 3502.690 1987.560 3503.010 ;
        RECT 1790.480 1772.070 1790.620 3502.690 ;
        RECT 1772.940 1771.750 1773.200 1772.070 ;
        RECT 1790.420 1771.750 1790.680 1772.070 ;
        RECT 1773.000 1767.165 1773.140 1771.750 ;
        RECT 1772.930 1766.795 1773.210 1767.165 ;
      LAYER via2 ;
        RECT 1772.930 1766.840 1773.210 1767.120 ;
      LAYER met3 ;
        RECT 1755.835 1767.130 1759.835 1767.135 ;
        RECT 1772.905 1767.130 1773.235 1767.145 ;
        RECT 1755.835 1766.830 1773.235 1767.130 ;
        RECT 1755.835 1766.535 1759.835 1766.830 ;
        RECT 1772.905 1766.815 1773.235 1766.830 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1662.510 3502.920 1662.830 3502.980 ;
        RECT 1776.130 3502.920 1776.450 3502.980 ;
        RECT 1662.510 3502.780 1776.450 3502.920 ;
        RECT 1662.510 3502.720 1662.830 3502.780 ;
        RECT 1776.130 3502.720 1776.450 3502.780 ;
        RECT 1464.710 1317.740 1465.030 1317.800 ;
        RECT 1776.130 1317.740 1776.450 1317.800 ;
        RECT 1464.710 1317.600 1776.450 1317.740 ;
        RECT 1464.710 1317.540 1465.030 1317.600 ;
        RECT 1776.130 1317.540 1776.450 1317.600 ;
      LAYER via ;
        RECT 1662.540 3502.720 1662.800 3502.980 ;
        RECT 1776.160 3502.720 1776.420 3502.980 ;
        RECT 1464.740 1317.540 1465.000 1317.800 ;
        RECT 1776.160 1317.540 1776.420 1317.800 ;
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
        RECT 1662.600 3503.010 1662.740 3517.600 ;
        RECT 1662.540 3502.690 1662.800 3503.010 ;
        RECT 1776.160 3502.690 1776.420 3503.010 ;
        RECT 1464.780 1323.135 1465.060 1327.135 ;
        RECT 1464.800 1317.830 1464.940 1323.135 ;
        RECT 1776.220 1317.830 1776.360 3502.690 ;
        RECT 1464.740 1317.510 1465.000 1317.830 ;
        RECT 1776.160 1317.510 1776.420 1317.830 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 727.865 1325.745 728.035 1327.615 ;
      LAYER mcon ;
        RECT 727.865 1327.445 728.035 1327.615 ;
      LAYER met1 ;
        RECT 693.750 3504.280 694.070 3504.340 ;
        RECT 1338.210 3504.280 1338.530 3504.340 ;
        RECT 693.750 3504.140 1338.530 3504.280 ;
        RECT 693.750 3504.080 694.070 3504.140 ;
        RECT 1338.210 3504.080 1338.530 3504.140 ;
        RECT 727.805 1327.600 728.095 1327.645 ;
        RECT 727.805 1327.460 856.360 1327.600 ;
        RECT 727.805 1327.415 728.095 1327.460 ;
        RECT 856.220 1326.640 856.360 1327.460 ;
        RECT 856.130 1326.380 856.450 1326.640 ;
        RECT 693.750 1325.900 694.070 1325.960 ;
        RECT 727.805 1325.900 728.095 1325.945 ;
        RECT 693.750 1325.760 728.095 1325.900 ;
        RECT 693.750 1325.700 694.070 1325.760 ;
        RECT 727.805 1325.715 728.095 1325.760 ;
      LAYER via ;
        RECT 693.780 3504.080 694.040 3504.340 ;
        RECT 1338.240 3504.080 1338.500 3504.340 ;
        RECT 856.160 1326.380 856.420 1326.640 ;
        RECT 693.780 1325.700 694.040 1325.960 ;
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
        RECT 1338.300 3504.370 1338.440 3517.600 ;
        RECT 693.780 3504.050 694.040 3504.370 ;
        RECT 1338.240 3504.050 1338.500 3504.370 ;
        RECT 693.840 1393.845 693.980 3504.050 ;
        RECT 693.770 1393.475 694.050 1393.845 ;
        RECT 693.770 1390.755 694.050 1391.125 ;
        RECT 693.840 1325.990 693.980 1390.755 ;
        RECT 856.160 1326.410 856.420 1326.670 ;
        RECT 856.660 1326.410 856.940 1327.135 ;
        RECT 856.160 1326.350 856.940 1326.410 ;
        RECT 856.220 1326.270 856.940 1326.350 ;
        RECT 693.780 1325.670 694.040 1325.990 ;
        RECT 856.660 1323.135 856.940 1326.270 ;
      LAYER via2 ;
        RECT 693.770 1393.520 694.050 1393.800 ;
        RECT 693.770 1390.800 694.050 1391.080 ;
      LAYER met3 ;
        RECT 693.745 1393.810 694.075 1393.825 ;
        RECT 693.745 1393.495 694.290 1393.810 ;
        RECT 693.990 1391.105 694.290 1393.495 ;
        RECT 693.745 1390.790 694.290 1391.105 ;
        RECT 693.745 1390.775 694.075 1390.790 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2283.510 436.120 2283.830 436.180 ;
        RECT 2318.010 436.120 2318.330 436.180 ;
        RECT 2283.510 435.980 2318.330 436.120 ;
        RECT 2283.510 435.920 2283.830 435.980 ;
        RECT 2318.010 435.920 2318.330 435.980 ;
        RECT 2089.390 435.780 2089.710 435.840 ;
        RECT 2124.810 435.780 2125.130 435.840 ;
        RECT 2089.390 435.640 2125.130 435.780 ;
        RECT 2089.390 435.580 2089.710 435.640 ;
        RECT 2124.810 435.580 2125.130 435.640 ;
      LAYER via ;
        RECT 2283.540 435.920 2283.800 436.180 ;
        RECT 2318.040 435.920 2318.300 436.180 ;
        RECT 2089.420 435.580 2089.680 435.840 ;
        RECT 2124.840 435.580 2125.100 435.840 ;
      LAYER met2 ;
        RECT 1016.690 2382.875 1016.970 2383.245 ;
        RECT 1016.760 2377.880 1016.900 2382.875 ;
        RECT 1016.740 2373.880 1017.020 2377.880 ;
        RECT 2221.430 438.755 2221.710 439.125 ;
        RECT 2149.210 437.395 2149.490 437.765 ;
        RECT 1931.630 436.715 1931.910 437.085 ;
        RECT 1931.700 435.725 1931.840 436.715 ;
        RECT 2124.830 436.035 2125.110 436.405 ;
        RECT 2124.900 435.870 2125.040 436.035 ;
        RECT 2089.420 435.725 2089.680 435.870 ;
        RECT 1931.630 435.355 1931.910 435.725 ;
        RECT 2089.410 435.355 2089.690 435.725 ;
        RECT 2124.840 435.550 2125.100 435.870 ;
        RECT 2149.280 435.045 2149.420 437.395 ;
        RECT 2221.500 437.085 2221.640 438.755 ;
        RECT 2221.430 436.715 2221.710 437.085 ;
        RECT 2283.540 435.890 2283.800 436.210 ;
        RECT 2318.030 436.035 2318.310 436.405 ;
        RECT 2627.610 436.035 2627.890 436.405 ;
        RECT 2318.040 435.890 2318.300 436.035 ;
        RECT 2283.600 435.725 2283.740 435.890 ;
        RECT 2283.530 435.355 2283.810 435.725 ;
        RECT 2627.680 435.045 2627.820 436.035 ;
        RECT 2149.210 434.675 2149.490 435.045 ;
        RECT 2627.610 434.675 2627.890 435.045 ;
      LAYER via2 ;
        RECT 1016.690 2382.920 1016.970 2383.200 ;
        RECT 2221.430 438.800 2221.710 439.080 ;
        RECT 2149.210 437.440 2149.490 437.720 ;
        RECT 1931.630 436.760 1931.910 437.040 ;
        RECT 2124.830 436.080 2125.110 436.360 ;
        RECT 1931.630 435.400 1931.910 435.680 ;
        RECT 2089.410 435.400 2089.690 435.680 ;
        RECT 2221.430 436.760 2221.710 437.040 ;
        RECT 2318.030 436.080 2318.310 436.360 ;
        RECT 2627.610 436.080 2627.890 436.360 ;
        RECT 2283.530 435.400 2283.810 435.680 ;
        RECT 2149.210 434.720 2149.490 435.000 ;
        RECT 2627.610 434.720 2627.890 435.000 ;
      LAYER met3 ;
        RECT 1016.665 2383.210 1016.995 2383.225 ;
        RECT 1779.550 2383.210 1779.930 2383.220 ;
        RECT 1016.665 2382.910 1779.930 2383.210 ;
        RECT 1016.665 2382.895 1016.995 2382.910 ;
        RECT 1779.550 2382.900 1779.930 2382.910 ;
        RECT 1779.550 1335.330 1779.930 1335.340 ;
        RECT 1779.550 1335.030 1780.810 1335.330 ;
        RECT 1779.550 1335.020 1779.930 1335.030 ;
        RECT 1779.550 1331.930 1779.930 1331.940 ;
        RECT 1780.510 1331.930 1780.810 1335.030 ;
        RECT 1779.550 1331.630 1780.810 1331.930 ;
        RECT 1779.550 1331.620 1779.930 1331.630 ;
        RECT 2917.600 439.770 2924.800 440.220 ;
        RECT 2916.710 439.470 2924.800 439.770 ;
        RECT 2173.310 439.090 2173.690 439.100 ;
        RECT 2221.405 439.090 2221.735 439.105 ;
        RECT 2173.310 438.790 2221.735 439.090 ;
        RECT 2173.310 438.780 2173.690 438.790 ;
        RECT 2221.405 438.775 2221.735 438.790 ;
        RECT 2149.185 437.730 2149.515 437.745 ;
        RECT 2173.310 437.730 2173.690 437.740 ;
        RECT 2149.185 437.430 2173.690 437.730 ;
        RECT 2149.185 437.415 2149.515 437.430 ;
        RECT 2173.310 437.420 2173.690 437.430 ;
        RECT 1883.510 437.050 1883.890 437.060 ;
        RECT 1931.605 437.050 1931.935 437.065 ;
        RECT 1883.510 436.750 1931.935 437.050 ;
        RECT 1883.510 436.740 1883.890 436.750 ;
        RECT 1931.605 436.735 1931.935 436.750 ;
        RECT 2221.405 437.050 2221.735 437.065 ;
        RECT 2221.405 436.750 2236.210 437.050 ;
        RECT 2221.405 436.735 2221.735 436.750 ;
        RECT 2124.805 436.370 2125.135 436.385 ;
        RECT 2125.470 436.370 2125.850 436.380 ;
        RECT 1800.750 436.070 1849.810 436.370 ;
        RECT 1779.550 435.010 1779.930 435.020 ;
        RECT 1800.750 435.010 1801.050 436.070 ;
        RECT 1779.550 434.710 1801.050 435.010 ;
        RECT 1849.510 435.010 1849.810 436.070 ;
        RECT 2015.110 436.070 2043.010 436.370 ;
        RECT 1931.605 435.690 1931.935 435.705 ;
        RECT 1931.605 435.390 2014.490 435.690 ;
        RECT 1931.605 435.375 1931.935 435.390 ;
        RECT 1883.510 435.010 1883.890 435.020 ;
        RECT 1849.510 434.710 1883.890 435.010 ;
        RECT 2014.190 435.010 2014.490 435.390 ;
        RECT 2015.110 435.010 2015.410 436.070 ;
        RECT 2042.710 435.690 2043.010 436.070 ;
        RECT 2124.805 436.070 2125.850 436.370 ;
        RECT 2124.805 436.055 2125.135 436.070 ;
        RECT 2125.470 436.060 2125.850 436.070 ;
        RECT 2089.385 435.690 2089.715 435.705 ;
        RECT 2042.710 435.390 2089.715 435.690 ;
        RECT 2235.910 435.690 2236.210 436.750 ;
        RECT 2318.005 436.370 2318.335 436.385 ;
        RECT 2627.585 436.370 2627.915 436.385 ;
        RECT 2318.005 436.070 2380.650 436.370 ;
        RECT 2318.005 436.055 2318.335 436.070 ;
        RECT 2283.505 435.690 2283.835 435.705 ;
        RECT 2235.910 435.390 2283.835 435.690 ;
        RECT 2380.350 435.690 2380.650 436.070 ;
        RECT 2524.790 436.070 2546.250 436.370 ;
        RECT 2524.790 435.690 2525.090 436.070 ;
        RECT 2380.350 435.390 2428.490 435.690 ;
        RECT 2089.385 435.375 2089.715 435.390 ;
        RECT 2283.505 435.375 2283.835 435.390 ;
        RECT 2014.190 434.710 2015.410 435.010 ;
        RECT 2125.470 435.010 2125.850 435.020 ;
        RECT 2149.185 435.010 2149.515 435.025 ;
        RECT 2125.470 434.710 2149.515 435.010 ;
        RECT 2428.190 435.010 2428.490 435.390 ;
        RECT 2476.950 435.390 2525.090 435.690 ;
        RECT 2545.950 435.690 2546.250 436.070 ;
        RECT 2594.710 436.070 2627.915 436.370 ;
        RECT 2545.950 435.390 2594.090 435.690 ;
        RECT 2476.950 435.010 2477.250 435.390 ;
        RECT 2428.190 434.710 2477.250 435.010 ;
        RECT 2593.790 435.010 2594.090 435.390 ;
        RECT 2594.710 435.010 2595.010 436.070 ;
        RECT 2627.585 436.055 2627.915 436.070 ;
        RECT 2656.310 436.370 2656.690 436.380 ;
        RECT 2656.310 436.070 2739.450 436.370 ;
        RECT 2656.310 436.060 2656.690 436.070 ;
        RECT 2739.150 435.690 2739.450 436.070 ;
        RECT 2787.910 436.070 2836.050 436.370 ;
        RECT 2739.150 435.390 2787.290 435.690 ;
        RECT 2593.790 434.710 2595.010 435.010 ;
        RECT 2627.585 435.010 2627.915 435.025 ;
        RECT 2656.310 435.010 2656.690 435.020 ;
        RECT 2627.585 434.710 2656.690 435.010 ;
        RECT 2786.990 435.010 2787.290 435.390 ;
        RECT 2787.910 435.010 2788.210 436.070 ;
        RECT 2835.750 435.690 2836.050 436.070 ;
        RECT 2916.710 435.690 2917.010 439.470 ;
        RECT 2917.600 439.020 2924.800 439.470 ;
        RECT 2835.750 435.390 2883.890 435.690 ;
        RECT 2786.990 434.710 2788.210 435.010 ;
        RECT 2883.590 435.010 2883.890 435.390 ;
        RECT 2884.510 435.390 2917.010 435.690 ;
        RECT 2884.510 435.010 2884.810 435.390 ;
        RECT 2883.590 434.710 2884.810 435.010 ;
        RECT 1779.550 434.700 1779.930 434.710 ;
        RECT 1883.510 434.700 1883.890 434.710 ;
        RECT 2125.470 434.700 2125.850 434.710 ;
        RECT 2149.185 434.695 2149.515 434.710 ;
        RECT 2627.585 434.695 2627.915 434.710 ;
        RECT 2656.310 434.700 2656.690 434.710 ;
      LAYER via3 ;
        RECT 1779.580 2382.900 1779.900 2383.220 ;
        RECT 1779.580 1335.020 1779.900 1335.340 ;
        RECT 1779.580 1331.620 1779.900 1331.940 ;
        RECT 2173.340 438.780 2173.660 439.100 ;
        RECT 2173.340 437.420 2173.660 437.740 ;
        RECT 1883.540 436.740 1883.860 437.060 ;
        RECT 1779.580 434.700 1779.900 435.020 ;
        RECT 1883.540 434.700 1883.860 435.020 ;
        RECT 2125.500 436.060 2125.820 436.380 ;
        RECT 2125.500 434.700 2125.820 435.020 ;
        RECT 2656.340 436.060 2656.660 436.380 ;
        RECT 2656.340 434.700 2656.660 435.020 ;
      LAYER met4 ;
        RECT 1779.575 2382.895 1779.905 2383.225 ;
        RECT 1779.590 1335.345 1779.890 2382.895 ;
        RECT 1779.575 1335.015 1779.905 1335.345 ;
        RECT 1779.575 1331.615 1779.905 1331.945 ;
        RECT 1779.590 435.025 1779.890 1331.615 ;
        RECT 2173.335 438.775 2173.665 439.105 ;
        RECT 2173.350 437.745 2173.650 438.775 ;
        RECT 2173.335 437.415 2173.665 437.745 ;
        RECT 1883.535 436.735 1883.865 437.065 ;
        RECT 1883.550 435.025 1883.850 436.735 ;
        RECT 2125.495 436.055 2125.825 436.385 ;
        RECT 2656.335 436.055 2656.665 436.385 ;
        RECT 2125.510 435.025 2125.810 436.055 ;
        RECT 2656.350 435.025 2656.650 436.055 ;
        RECT 1779.575 434.695 1779.905 435.025 ;
        RECT 1883.535 434.695 1883.865 435.025 ;
        RECT 2125.495 434.695 2125.825 435.025 ;
        RECT 2656.335 434.695 2656.665 435.025 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1753.665 3429.665 1753.835 3443.775 ;
        RECT 1754.125 3139.645 1754.295 3175.515 ;
        RECT 1751.825 2642.905 1751.995 2691.015 ;
        RECT 1753.205 2429.725 1753.375 2463.215 ;
        RECT 1755.965 2373.625 1756.135 2414.935 ;
      LAYER mcon ;
        RECT 1753.665 3443.605 1753.835 3443.775 ;
        RECT 1754.125 3175.345 1754.295 3175.515 ;
        RECT 1751.825 2690.845 1751.995 2691.015 ;
        RECT 1753.205 2463.045 1753.375 2463.215 ;
        RECT 1755.965 2414.765 1756.135 2414.935 ;
      LAYER met1 ;
        RECT 1013.910 3503.940 1014.230 3504.000 ;
        RECT 1753.590 3503.940 1753.910 3504.000 ;
        RECT 1013.910 3503.800 1753.910 3503.940 ;
        RECT 1013.910 3503.740 1014.230 3503.800 ;
        RECT 1753.590 3503.740 1753.910 3503.800 ;
        RECT 1753.590 3443.760 1753.910 3443.820 ;
        RECT 1753.395 3443.620 1753.910 3443.760 ;
        RECT 1753.590 3443.560 1753.910 3443.620 ;
        RECT 1753.590 3429.820 1753.910 3429.880 ;
        RECT 1753.395 3429.680 1753.910 3429.820 ;
        RECT 1753.590 3429.620 1753.910 3429.680 ;
        RECT 1752.670 3429.140 1752.990 3429.200 ;
        RECT 1753.590 3429.140 1753.910 3429.200 ;
        RECT 1752.670 3429.000 1753.910 3429.140 ;
        RECT 1752.670 3428.940 1752.990 3429.000 ;
        RECT 1753.590 3428.940 1753.910 3429.000 ;
        RECT 1752.670 3340.400 1752.990 3340.460 ;
        RECT 1754.510 3340.400 1754.830 3340.460 ;
        RECT 1752.670 3340.260 1754.830 3340.400 ;
        RECT 1752.670 3340.200 1752.990 3340.260 ;
        RECT 1754.510 3340.200 1754.830 3340.260 ;
        RECT 1754.510 3284.980 1754.830 3285.040 ;
        RECT 1752.760 3284.840 1754.830 3284.980 ;
        RECT 1752.760 3284.700 1752.900 3284.840 ;
        RECT 1754.510 3284.780 1754.830 3284.840 ;
        RECT 1752.670 3284.440 1752.990 3284.700 ;
        RECT 1752.670 3202.020 1752.990 3202.080 ;
        RECT 1753.590 3202.020 1753.910 3202.080 ;
        RECT 1752.670 3201.880 1753.910 3202.020 ;
        RECT 1752.670 3201.820 1752.990 3201.880 ;
        RECT 1753.590 3201.820 1753.910 3201.880 ;
        RECT 1752.670 3175.500 1752.990 3175.560 ;
        RECT 1754.065 3175.500 1754.355 3175.545 ;
        RECT 1752.670 3175.360 1754.355 3175.500 ;
        RECT 1752.670 3175.300 1752.990 3175.360 ;
        RECT 1754.065 3175.315 1754.355 3175.360 ;
        RECT 1754.050 3139.800 1754.370 3139.860 ;
        RECT 1753.855 3139.660 1754.370 3139.800 ;
        RECT 1754.050 3139.600 1754.370 3139.660 ;
        RECT 1752.670 3105.460 1752.990 3105.520 ;
        RECT 1754.050 3105.460 1754.370 3105.520 ;
        RECT 1752.670 3105.320 1754.370 3105.460 ;
        RECT 1752.670 3105.260 1752.990 3105.320 ;
        RECT 1754.050 3105.260 1754.370 3105.320 ;
        RECT 1752.670 3056.640 1752.990 3056.900 ;
        RECT 1752.760 3056.500 1752.900 3056.640 ;
        RECT 1753.590 3056.500 1753.910 3056.560 ;
        RECT 1752.760 3056.360 1753.910 3056.500 ;
        RECT 1753.590 3056.300 1753.910 3056.360 ;
        RECT 1753.590 2995.300 1753.910 2995.360 ;
        RECT 1752.760 2995.160 1753.910 2995.300 ;
        RECT 1752.760 2995.020 1752.900 2995.160 ;
        RECT 1753.590 2995.100 1753.910 2995.160 ;
        RECT 1752.670 2994.760 1752.990 2995.020 ;
        RECT 1752.670 2989.520 1752.990 2989.580 ;
        RECT 1754.050 2989.520 1754.370 2989.580 ;
        RECT 1752.670 2989.380 1754.370 2989.520 ;
        RECT 1752.670 2989.320 1752.990 2989.380 ;
        RECT 1754.050 2989.320 1754.370 2989.380 ;
        RECT 1754.050 2946.140 1754.370 2946.400 ;
        RECT 1751.750 2946.000 1752.070 2946.060 ;
        RECT 1754.140 2946.000 1754.280 2946.140 ;
        RECT 1751.750 2945.860 1754.280 2946.000 ;
        RECT 1751.750 2945.800 1752.070 2945.860 ;
        RECT 1751.750 2876.300 1752.070 2876.360 ;
        RECT 1754.510 2876.300 1754.830 2876.360 ;
        RECT 1751.750 2876.160 1754.830 2876.300 ;
        RECT 1751.750 2876.100 1752.070 2876.160 ;
        RECT 1754.510 2876.100 1754.830 2876.160 ;
        RECT 1753.130 2715.140 1753.450 2715.200 ;
        RECT 1754.050 2715.140 1754.370 2715.200 ;
        RECT 1753.130 2715.000 1754.370 2715.140 ;
        RECT 1753.130 2714.940 1753.450 2715.000 ;
        RECT 1754.050 2714.940 1754.370 2715.000 ;
        RECT 1751.765 2691.000 1752.055 2691.045 ;
        RECT 1753.130 2691.000 1753.450 2691.060 ;
        RECT 1751.765 2690.860 1753.450 2691.000 ;
        RECT 1751.765 2690.815 1752.055 2690.860 ;
        RECT 1753.130 2690.800 1753.450 2690.860 ;
        RECT 1751.750 2643.060 1752.070 2643.120 ;
        RECT 1751.555 2642.920 1752.070 2643.060 ;
        RECT 1751.750 2642.860 1752.070 2642.920 ;
        RECT 1751.750 2594.780 1752.070 2594.840 ;
        RECT 1752.670 2594.780 1752.990 2594.840 ;
        RECT 1751.750 2594.640 1752.990 2594.780 ;
        RECT 1751.750 2594.580 1752.070 2594.640 ;
        RECT 1752.670 2594.580 1752.990 2594.640 ;
        RECT 1752.670 2476.940 1752.990 2477.200 ;
        RECT 1752.760 2476.460 1752.900 2476.940 ;
        RECT 1753.130 2476.460 1753.450 2476.520 ;
        RECT 1752.760 2476.320 1753.450 2476.460 ;
        RECT 1753.130 2476.260 1753.450 2476.320 ;
        RECT 1753.130 2463.200 1753.450 2463.260 ;
        RECT 1752.935 2463.060 1753.450 2463.200 ;
        RECT 1753.130 2463.000 1753.450 2463.060 ;
        RECT 1753.145 2429.880 1753.435 2429.925 ;
        RECT 1753.590 2429.880 1753.910 2429.940 ;
        RECT 1753.145 2429.740 1753.910 2429.880 ;
        RECT 1753.145 2429.695 1753.435 2429.740 ;
        RECT 1753.590 2429.680 1753.910 2429.740 ;
        RECT 1753.590 2414.920 1753.910 2414.980 ;
        RECT 1755.905 2414.920 1756.195 2414.965 ;
        RECT 1753.590 2414.780 1756.195 2414.920 ;
        RECT 1753.590 2414.720 1753.910 2414.780 ;
        RECT 1755.905 2414.735 1756.195 2414.780 ;
        RECT 1754.970 2373.780 1755.290 2373.840 ;
        RECT 1755.905 2373.780 1756.195 2373.825 ;
        RECT 1754.970 2373.640 1756.195 2373.780 ;
        RECT 1754.970 2373.580 1755.290 2373.640 ;
        RECT 1755.905 2373.595 1756.195 2373.640 ;
        RECT 1754.970 2256.140 1755.290 2256.200 ;
        RECT 1756.810 2256.140 1757.130 2256.200 ;
        RECT 1754.970 2256.000 1757.130 2256.140 ;
        RECT 1754.970 2255.940 1755.290 2256.000 ;
        RECT 1756.810 2255.940 1757.130 2256.000 ;
      LAYER via ;
        RECT 1013.940 3503.740 1014.200 3504.000 ;
        RECT 1753.620 3503.740 1753.880 3504.000 ;
        RECT 1753.620 3443.560 1753.880 3443.820 ;
        RECT 1753.620 3429.620 1753.880 3429.880 ;
        RECT 1752.700 3428.940 1752.960 3429.200 ;
        RECT 1753.620 3428.940 1753.880 3429.200 ;
        RECT 1752.700 3340.200 1752.960 3340.460 ;
        RECT 1754.540 3340.200 1754.800 3340.460 ;
        RECT 1754.540 3284.780 1754.800 3285.040 ;
        RECT 1752.700 3284.440 1752.960 3284.700 ;
        RECT 1752.700 3201.820 1752.960 3202.080 ;
        RECT 1753.620 3201.820 1753.880 3202.080 ;
        RECT 1752.700 3175.300 1752.960 3175.560 ;
        RECT 1754.080 3139.600 1754.340 3139.860 ;
        RECT 1752.700 3105.260 1752.960 3105.520 ;
        RECT 1754.080 3105.260 1754.340 3105.520 ;
        RECT 1752.700 3056.640 1752.960 3056.900 ;
        RECT 1753.620 3056.300 1753.880 3056.560 ;
        RECT 1753.620 2995.100 1753.880 2995.360 ;
        RECT 1752.700 2994.760 1752.960 2995.020 ;
        RECT 1752.700 2989.320 1752.960 2989.580 ;
        RECT 1754.080 2989.320 1754.340 2989.580 ;
        RECT 1754.080 2946.140 1754.340 2946.400 ;
        RECT 1751.780 2945.800 1752.040 2946.060 ;
        RECT 1751.780 2876.100 1752.040 2876.360 ;
        RECT 1754.540 2876.100 1754.800 2876.360 ;
        RECT 1753.160 2714.940 1753.420 2715.200 ;
        RECT 1754.080 2714.940 1754.340 2715.200 ;
        RECT 1753.160 2690.800 1753.420 2691.060 ;
        RECT 1751.780 2642.860 1752.040 2643.120 ;
        RECT 1751.780 2594.580 1752.040 2594.840 ;
        RECT 1752.700 2594.580 1752.960 2594.840 ;
        RECT 1752.700 2476.940 1752.960 2477.200 ;
        RECT 1753.160 2476.260 1753.420 2476.520 ;
        RECT 1753.160 2463.000 1753.420 2463.260 ;
        RECT 1753.620 2429.680 1753.880 2429.940 ;
        RECT 1753.620 2414.720 1753.880 2414.980 ;
        RECT 1755.000 2373.580 1755.260 2373.840 ;
        RECT 1755.000 2255.940 1755.260 2256.200 ;
        RECT 1756.840 2255.940 1757.100 2256.200 ;
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
        RECT 1014.000 3504.030 1014.140 3517.600 ;
        RECT 1013.940 3503.710 1014.200 3504.030 ;
        RECT 1753.620 3503.710 1753.880 3504.030 ;
        RECT 1753.680 3443.850 1753.820 3503.710 ;
        RECT 1753.620 3443.530 1753.880 3443.850 ;
        RECT 1753.620 3429.590 1753.880 3429.910 ;
        RECT 1753.680 3429.230 1753.820 3429.590 ;
        RECT 1752.700 3428.910 1752.960 3429.230 ;
        RECT 1753.620 3428.910 1753.880 3429.230 ;
        RECT 1752.760 3340.490 1752.900 3428.910 ;
        RECT 1752.700 3340.170 1752.960 3340.490 ;
        RECT 1754.540 3340.170 1754.800 3340.490 ;
        RECT 1754.600 3285.070 1754.740 3340.170 ;
        RECT 1754.540 3284.750 1754.800 3285.070 ;
        RECT 1752.700 3284.410 1752.960 3284.730 ;
        RECT 1752.760 3249.450 1752.900 3284.410 ;
        RECT 1752.760 3249.310 1753.820 3249.450 ;
        RECT 1753.680 3202.110 1753.820 3249.310 ;
        RECT 1752.700 3201.790 1752.960 3202.110 ;
        RECT 1753.620 3201.790 1753.880 3202.110 ;
        RECT 1752.760 3175.590 1752.900 3201.790 ;
        RECT 1752.700 3175.270 1752.960 3175.590 ;
        RECT 1754.080 3139.570 1754.340 3139.890 ;
        RECT 1754.140 3105.550 1754.280 3139.570 ;
        RECT 1752.700 3105.230 1752.960 3105.550 ;
        RECT 1754.080 3105.230 1754.340 3105.550 ;
        RECT 1752.760 3056.930 1752.900 3105.230 ;
        RECT 1752.700 3056.610 1752.960 3056.930 ;
        RECT 1753.620 3056.270 1753.880 3056.590 ;
        RECT 1753.680 2995.390 1753.820 3056.270 ;
        RECT 1753.620 2995.070 1753.880 2995.390 ;
        RECT 1752.700 2994.730 1752.960 2995.050 ;
        RECT 1752.760 2989.610 1752.900 2994.730 ;
        RECT 1752.700 2989.290 1752.960 2989.610 ;
        RECT 1754.080 2989.290 1754.340 2989.610 ;
        RECT 1754.140 2946.430 1754.280 2989.290 ;
        RECT 1754.080 2946.110 1754.340 2946.430 ;
        RECT 1751.780 2945.770 1752.040 2946.090 ;
        RECT 1751.840 2939.485 1751.980 2945.770 ;
        RECT 1750.850 2939.115 1751.130 2939.485 ;
        RECT 1751.770 2939.115 1752.050 2939.485 ;
        RECT 1750.920 2896.530 1751.060 2939.115 ;
        RECT 1750.920 2896.390 1751.980 2896.530 ;
        RECT 1751.840 2876.390 1751.980 2896.390 ;
        RECT 1751.780 2876.070 1752.040 2876.390 ;
        RECT 1754.540 2876.070 1754.800 2876.390 ;
        RECT 1754.600 2802.690 1754.740 2876.070 ;
        RECT 1754.140 2802.550 1754.740 2802.690 ;
        RECT 1754.140 2767.330 1754.280 2802.550 ;
        RECT 1754.140 2767.190 1754.740 2767.330 ;
        RECT 1754.600 2766.650 1754.740 2767.190 ;
        RECT 1754.140 2766.510 1754.740 2766.650 ;
        RECT 1754.140 2715.230 1754.280 2766.510 ;
        RECT 1753.160 2714.910 1753.420 2715.230 ;
        RECT 1754.080 2714.910 1754.340 2715.230 ;
        RECT 1753.220 2691.090 1753.360 2714.910 ;
        RECT 1753.160 2690.770 1753.420 2691.090 ;
        RECT 1751.780 2642.830 1752.040 2643.150 ;
        RECT 1751.840 2594.870 1751.980 2642.830 ;
        RECT 1751.780 2594.550 1752.040 2594.870 ;
        RECT 1752.700 2594.550 1752.960 2594.870 ;
        RECT 1752.760 2477.230 1752.900 2594.550 ;
        RECT 1752.700 2476.910 1752.960 2477.230 ;
        RECT 1753.160 2476.230 1753.420 2476.550 ;
        RECT 1753.220 2463.290 1753.360 2476.230 ;
        RECT 1753.160 2462.970 1753.420 2463.290 ;
        RECT 1753.620 2429.650 1753.880 2429.970 ;
        RECT 1753.680 2415.010 1753.820 2429.650 ;
        RECT 1753.620 2414.690 1753.880 2415.010 ;
        RECT 1755.000 2373.550 1755.260 2373.870 ;
        RECT 1755.060 2320.570 1755.200 2373.550 ;
        RECT 1755.060 2320.430 1755.660 2320.570 ;
        RECT 1755.520 2312.410 1755.660 2320.430 ;
        RECT 1755.060 2312.270 1755.660 2312.410 ;
        RECT 1755.060 2256.230 1755.200 2312.270 ;
        RECT 1755.000 2255.910 1755.260 2256.230 ;
        RECT 1756.840 2256.085 1757.100 2256.230 ;
        RECT 1756.830 2255.715 1757.110 2256.085 ;
      LAYER via2 ;
        RECT 1750.850 2939.160 1751.130 2939.440 ;
        RECT 1751.770 2939.160 1752.050 2939.440 ;
        RECT 1756.830 2255.760 1757.110 2256.040 ;
      LAYER met3 ;
        RECT 1750.825 2939.450 1751.155 2939.465 ;
        RECT 1751.745 2939.450 1752.075 2939.465 ;
        RECT 1750.825 2939.150 1752.075 2939.450 ;
        RECT 1750.825 2939.135 1751.155 2939.150 ;
        RECT 1751.745 2939.135 1752.075 2939.150 ;
        RECT 1756.805 2256.050 1757.135 2256.065 ;
        RECT 1756.590 2255.735 1757.135 2256.050 ;
        RECT 1756.590 2254.015 1756.890 2255.735 ;
        RECT 1755.835 2253.415 1759.835 2254.015 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 689.150 3503.600 689.470 3503.660 ;
        RECT 1455.970 3503.600 1456.290 3503.660 ;
        RECT 689.150 3503.460 1456.290 3503.600 ;
        RECT 689.150 3503.400 689.470 3503.460 ;
        RECT 1455.970 3503.400 1456.290 3503.460 ;
      LAYER via ;
        RECT 689.180 3503.400 689.440 3503.660 ;
        RECT 1456.000 3503.400 1456.260 3503.660 ;
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
        RECT 689.240 3503.690 689.380 3517.600 ;
        RECT 689.180 3503.370 689.440 3503.690 ;
        RECT 1456.000 3503.370 1456.260 3503.690 ;
        RECT 1456.060 2377.690 1456.200 3503.370 ;
        RECT 1456.500 2377.690 1456.780 2377.880 ;
        RECT 1456.060 2377.550 1456.780 2377.690 ;
        RECT 1456.500 2373.880 1456.780 2377.550 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1755.045 3278.025 1755.215 3332.595 ;
        RECT 1754.585 3235.525 1754.755 3277.515 ;
        RECT 1755.045 3133.185 1755.215 3180.955 ;
        RECT 1755.045 2898.245 1755.215 2946.355 ;
        RECT 1755.965 2698.325 1756.135 2704.955 ;
        RECT 1754.585 2297.125 1754.755 2343.195 ;
        RECT 1755.505 2283.865 1755.675 2297.295 ;
        RECT 1755.045 2035.665 1755.215 2044.335 ;
      LAYER mcon ;
        RECT 1755.045 3332.425 1755.215 3332.595 ;
        RECT 1754.585 3277.345 1754.755 3277.515 ;
        RECT 1755.045 3180.785 1755.215 3180.955 ;
        RECT 1755.045 2946.185 1755.215 2946.355 ;
        RECT 1755.965 2704.785 1756.135 2704.955 ;
        RECT 1754.585 2343.025 1754.755 2343.195 ;
        RECT 1755.505 2297.125 1755.675 2297.295 ;
        RECT 1755.045 2044.165 1755.215 2044.335 ;
      LAYER met1 ;
        RECT 364.850 3502.580 365.170 3502.640 ;
        RECT 1754.970 3502.580 1755.290 3502.640 ;
        RECT 364.850 3502.440 1755.290 3502.580 ;
        RECT 364.850 3502.380 365.170 3502.440 ;
        RECT 1754.970 3502.380 1755.290 3502.440 ;
        RECT 1754.970 3443.420 1755.290 3443.480 ;
        RECT 1754.600 3443.280 1755.290 3443.420 ;
        RECT 1754.600 3443.140 1754.740 3443.280 ;
        RECT 1754.970 3443.220 1755.290 3443.280 ;
        RECT 1754.510 3442.880 1754.830 3443.140 ;
        RECT 1754.050 3428.800 1754.370 3428.860 ;
        RECT 1754.510 3428.800 1754.830 3428.860 ;
        RECT 1754.050 3428.660 1754.830 3428.800 ;
        RECT 1754.050 3428.600 1754.370 3428.660 ;
        RECT 1754.510 3428.600 1754.830 3428.660 ;
        RECT 1754.970 3346.660 1755.290 3346.920 ;
        RECT 1755.060 3346.180 1755.200 3346.660 ;
        RECT 1755.430 3346.180 1755.750 3346.240 ;
        RECT 1755.060 3346.040 1755.750 3346.180 ;
        RECT 1755.430 3345.980 1755.750 3346.040 ;
        RECT 1754.985 3332.580 1755.275 3332.625 ;
        RECT 1755.430 3332.580 1755.750 3332.640 ;
        RECT 1754.985 3332.440 1755.750 3332.580 ;
        RECT 1754.985 3332.395 1755.275 3332.440 ;
        RECT 1755.430 3332.380 1755.750 3332.440 ;
        RECT 1754.970 3278.180 1755.290 3278.240 ;
        RECT 1754.775 3278.040 1755.290 3278.180 ;
        RECT 1754.970 3277.980 1755.290 3278.040 ;
        RECT 1754.510 3277.500 1754.830 3277.560 ;
        RECT 1754.315 3277.360 1754.830 3277.500 ;
        RECT 1754.510 3277.300 1754.830 3277.360 ;
        RECT 1754.525 3235.680 1754.815 3235.725 ;
        RECT 1754.970 3235.680 1755.290 3235.740 ;
        RECT 1754.525 3235.540 1755.290 3235.680 ;
        RECT 1754.525 3235.495 1754.815 3235.540 ;
        RECT 1754.970 3235.480 1755.290 3235.540 ;
        RECT 1754.970 3187.740 1755.290 3187.800 ;
        RECT 1755.430 3187.740 1755.750 3187.800 ;
        RECT 1754.970 3187.600 1755.750 3187.740 ;
        RECT 1754.970 3187.540 1755.290 3187.600 ;
        RECT 1755.430 3187.540 1755.750 3187.600 ;
        RECT 1754.985 3180.940 1755.275 3180.985 ;
        RECT 1755.430 3180.940 1755.750 3181.000 ;
        RECT 1754.985 3180.800 1755.750 3180.940 ;
        RECT 1754.985 3180.755 1755.275 3180.800 ;
        RECT 1755.430 3180.740 1755.750 3180.800 ;
        RECT 1754.970 3133.340 1755.290 3133.400 ;
        RECT 1754.775 3133.200 1755.290 3133.340 ;
        RECT 1754.970 3133.140 1755.290 3133.200 ;
        RECT 1753.590 3084.380 1753.910 3084.440 ;
        RECT 1755.430 3084.380 1755.750 3084.440 ;
        RECT 1753.590 3084.240 1755.750 3084.380 ;
        RECT 1753.590 3084.180 1753.910 3084.240 ;
        RECT 1755.430 3084.180 1755.750 3084.240 ;
        RECT 1754.970 2995.300 1755.290 2995.360 ;
        RECT 1755.430 2995.300 1755.750 2995.360 ;
        RECT 1754.970 2995.160 1755.750 2995.300 ;
        RECT 1754.970 2995.100 1755.290 2995.160 ;
        RECT 1755.430 2995.100 1755.750 2995.160 ;
        RECT 1754.970 2946.340 1755.290 2946.400 ;
        RECT 1754.775 2946.200 1755.290 2946.340 ;
        RECT 1754.970 2946.140 1755.290 2946.200 ;
        RECT 1754.510 2898.400 1754.830 2898.460 ;
        RECT 1754.985 2898.400 1755.275 2898.445 ;
        RECT 1754.510 2898.260 1755.275 2898.400 ;
        RECT 1754.510 2898.200 1754.830 2898.260 ;
        RECT 1754.985 2898.215 1755.275 2898.260 ;
        RECT 1754.970 2849.780 1755.290 2849.840 ;
        RECT 1755.890 2849.780 1756.210 2849.840 ;
        RECT 1754.970 2849.640 1756.210 2849.780 ;
        RECT 1754.970 2849.580 1755.290 2849.640 ;
        RECT 1755.890 2849.580 1756.210 2849.640 ;
        RECT 1754.970 2801.840 1755.290 2801.900 ;
        RECT 1755.890 2801.840 1756.210 2801.900 ;
        RECT 1754.970 2801.700 1756.210 2801.840 ;
        RECT 1754.970 2801.640 1755.290 2801.700 ;
        RECT 1755.890 2801.640 1756.210 2801.700 ;
        RECT 1754.970 2753.220 1755.290 2753.280 ;
        RECT 1755.890 2753.220 1756.210 2753.280 ;
        RECT 1754.970 2753.080 1756.210 2753.220 ;
        RECT 1754.970 2753.020 1755.290 2753.080 ;
        RECT 1755.890 2753.020 1756.210 2753.080 ;
        RECT 1755.890 2704.940 1756.210 2705.000 ;
        RECT 1755.695 2704.800 1756.210 2704.940 ;
        RECT 1755.890 2704.740 1756.210 2704.800 ;
        RECT 1755.890 2698.480 1756.210 2698.540 ;
        RECT 1755.695 2698.340 1756.210 2698.480 ;
        RECT 1755.890 2698.280 1756.210 2698.340 ;
        RECT 1754.510 2642.720 1754.830 2642.780 ;
        RECT 1755.430 2642.720 1755.750 2642.780 ;
        RECT 1754.510 2642.580 1755.750 2642.720 ;
        RECT 1754.510 2642.520 1754.830 2642.580 ;
        RECT 1755.430 2642.520 1755.750 2642.580 ;
        RECT 1754.970 2511.820 1755.290 2511.880 ;
        RECT 1755.430 2511.820 1755.750 2511.880 ;
        RECT 1754.970 2511.680 1755.750 2511.820 ;
        RECT 1754.970 2511.620 1755.290 2511.680 ;
        RECT 1755.430 2511.620 1755.750 2511.680 ;
        RECT 1754.510 2423.080 1754.830 2423.140 ;
        RECT 1756.350 2423.080 1756.670 2423.140 ;
        RECT 1754.510 2422.940 1756.670 2423.080 ;
        RECT 1754.510 2422.880 1754.830 2422.940 ;
        RECT 1756.350 2422.880 1756.670 2422.940 ;
        RECT 1754.510 2343.180 1754.830 2343.240 ;
        RECT 1754.315 2343.040 1754.830 2343.180 ;
        RECT 1754.510 2342.980 1754.830 2343.040 ;
        RECT 1754.525 2297.280 1754.815 2297.325 ;
        RECT 1755.445 2297.280 1755.735 2297.325 ;
        RECT 1754.525 2297.140 1755.735 2297.280 ;
        RECT 1754.525 2297.095 1754.815 2297.140 ;
        RECT 1755.445 2297.095 1755.735 2297.140 ;
        RECT 1754.510 2284.020 1754.830 2284.080 ;
        RECT 1755.445 2284.020 1755.735 2284.065 ;
        RECT 1754.510 2283.880 1755.735 2284.020 ;
        RECT 1754.510 2283.820 1754.830 2283.880 ;
        RECT 1755.445 2283.835 1755.735 2283.880 ;
        RECT 1754.510 2044.320 1754.830 2044.380 ;
        RECT 1754.985 2044.320 1755.275 2044.365 ;
        RECT 1754.510 2044.180 1755.275 2044.320 ;
        RECT 1754.510 2044.120 1754.830 2044.180 ;
        RECT 1754.985 2044.135 1755.275 2044.180 ;
        RECT 1754.510 2035.820 1754.830 2035.880 ;
        RECT 1754.985 2035.820 1755.275 2035.865 ;
        RECT 1754.510 2035.680 1755.275 2035.820 ;
        RECT 1754.510 2035.620 1754.830 2035.680 ;
        RECT 1754.985 2035.635 1755.275 2035.680 ;
        RECT 1754.970 1759.400 1755.290 1759.460 ;
        RECT 1757.730 1759.400 1758.050 1759.460 ;
        RECT 1754.970 1759.260 1758.050 1759.400 ;
        RECT 1754.970 1759.200 1755.290 1759.260 ;
        RECT 1757.730 1759.200 1758.050 1759.260 ;
      LAYER via ;
        RECT 364.880 3502.380 365.140 3502.640 ;
        RECT 1755.000 3502.380 1755.260 3502.640 ;
        RECT 1755.000 3443.220 1755.260 3443.480 ;
        RECT 1754.540 3442.880 1754.800 3443.140 ;
        RECT 1754.080 3428.600 1754.340 3428.860 ;
        RECT 1754.540 3428.600 1754.800 3428.860 ;
        RECT 1755.000 3346.660 1755.260 3346.920 ;
        RECT 1755.460 3345.980 1755.720 3346.240 ;
        RECT 1755.460 3332.380 1755.720 3332.640 ;
        RECT 1755.000 3277.980 1755.260 3278.240 ;
        RECT 1754.540 3277.300 1754.800 3277.560 ;
        RECT 1755.000 3235.480 1755.260 3235.740 ;
        RECT 1755.000 3187.540 1755.260 3187.800 ;
        RECT 1755.460 3187.540 1755.720 3187.800 ;
        RECT 1755.460 3180.740 1755.720 3181.000 ;
        RECT 1755.000 3133.140 1755.260 3133.400 ;
        RECT 1753.620 3084.180 1753.880 3084.440 ;
        RECT 1755.460 3084.180 1755.720 3084.440 ;
        RECT 1755.000 2995.100 1755.260 2995.360 ;
        RECT 1755.460 2995.100 1755.720 2995.360 ;
        RECT 1755.000 2946.140 1755.260 2946.400 ;
        RECT 1754.540 2898.200 1754.800 2898.460 ;
        RECT 1755.000 2849.580 1755.260 2849.840 ;
        RECT 1755.920 2849.580 1756.180 2849.840 ;
        RECT 1755.000 2801.640 1755.260 2801.900 ;
        RECT 1755.920 2801.640 1756.180 2801.900 ;
        RECT 1755.000 2753.020 1755.260 2753.280 ;
        RECT 1755.920 2753.020 1756.180 2753.280 ;
        RECT 1755.920 2704.740 1756.180 2705.000 ;
        RECT 1755.920 2698.280 1756.180 2698.540 ;
        RECT 1754.540 2642.520 1754.800 2642.780 ;
        RECT 1755.460 2642.520 1755.720 2642.780 ;
        RECT 1755.000 2511.620 1755.260 2511.880 ;
        RECT 1755.460 2511.620 1755.720 2511.880 ;
        RECT 1754.540 2422.880 1754.800 2423.140 ;
        RECT 1756.380 2422.880 1756.640 2423.140 ;
        RECT 1754.540 2342.980 1754.800 2343.240 ;
        RECT 1754.540 2283.820 1754.800 2284.080 ;
        RECT 1754.540 2044.120 1754.800 2044.380 ;
        RECT 1754.540 2035.620 1754.800 2035.880 ;
        RECT 1755.000 1759.200 1755.260 1759.460 ;
        RECT 1757.760 1759.200 1758.020 1759.460 ;
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
        RECT 364.940 3502.670 365.080 3517.600 ;
        RECT 364.880 3502.350 365.140 3502.670 ;
        RECT 1755.000 3502.350 1755.260 3502.670 ;
        RECT 1755.060 3443.510 1755.200 3502.350 ;
        RECT 1755.000 3443.190 1755.260 3443.510 ;
        RECT 1754.540 3442.850 1754.800 3443.170 ;
        RECT 1754.600 3428.890 1754.740 3442.850 ;
        RECT 1754.080 3428.570 1754.340 3428.890 ;
        RECT 1754.540 3428.570 1754.800 3428.890 ;
        RECT 1754.140 3381.370 1754.280 3428.570 ;
        RECT 1754.140 3381.230 1755.200 3381.370 ;
        RECT 1755.060 3346.950 1755.200 3381.230 ;
        RECT 1755.000 3346.630 1755.260 3346.950 ;
        RECT 1755.460 3345.950 1755.720 3346.270 ;
        RECT 1755.520 3332.670 1755.660 3345.950 ;
        RECT 1755.460 3332.350 1755.720 3332.670 ;
        RECT 1755.000 3278.010 1755.260 3278.270 ;
        RECT 1754.600 3277.950 1755.260 3278.010 ;
        RECT 1754.600 3277.870 1755.200 3277.950 ;
        RECT 1754.600 3277.590 1754.740 3277.870 ;
        RECT 1754.540 3277.270 1754.800 3277.590 ;
        RECT 1755.000 3235.450 1755.260 3235.770 ;
        RECT 1755.060 3187.830 1755.200 3235.450 ;
        RECT 1755.000 3187.510 1755.260 3187.830 ;
        RECT 1755.460 3187.510 1755.720 3187.830 ;
        RECT 1755.520 3181.030 1755.660 3187.510 ;
        RECT 1755.460 3180.710 1755.720 3181.030 ;
        RECT 1755.000 3133.110 1755.260 3133.430 ;
        RECT 1753.610 3132.235 1753.890 3132.605 ;
        RECT 1754.530 3132.490 1754.810 3132.605 ;
        RECT 1755.060 3132.490 1755.200 3133.110 ;
        RECT 1754.530 3132.350 1755.200 3132.490 ;
        RECT 1754.530 3132.235 1754.810 3132.350 ;
        RECT 1753.680 3084.470 1753.820 3132.235 ;
        RECT 1753.620 3084.150 1753.880 3084.470 ;
        RECT 1755.460 3084.150 1755.720 3084.470 ;
        RECT 1755.520 2995.390 1755.660 3084.150 ;
        RECT 1755.000 2995.070 1755.260 2995.390 ;
        RECT 1755.460 2995.070 1755.720 2995.390 ;
        RECT 1755.060 2946.430 1755.200 2995.070 ;
        RECT 1755.000 2946.110 1755.260 2946.430 ;
        RECT 1754.540 2898.400 1754.800 2898.490 ;
        RECT 1754.540 2898.260 1755.200 2898.400 ;
        RECT 1754.540 2898.170 1754.800 2898.260 ;
        RECT 1755.060 2898.005 1755.200 2898.260 ;
        RECT 1754.990 2897.635 1755.270 2898.005 ;
        RECT 1755.910 2897.635 1756.190 2898.005 ;
        RECT 1755.980 2849.870 1756.120 2897.635 ;
        RECT 1755.000 2849.725 1755.260 2849.870 ;
        RECT 1755.920 2849.725 1756.180 2849.870 ;
        RECT 1754.990 2849.355 1755.270 2849.725 ;
        RECT 1755.910 2849.355 1756.190 2849.725 ;
        RECT 1755.980 2801.930 1756.120 2849.355 ;
        RECT 1755.000 2801.610 1755.260 2801.930 ;
        RECT 1755.920 2801.610 1756.180 2801.930 ;
        RECT 1755.060 2801.445 1755.200 2801.610 ;
        RECT 1754.990 2801.075 1755.270 2801.445 ;
        RECT 1755.910 2801.075 1756.190 2801.445 ;
        RECT 1755.980 2753.310 1756.120 2801.075 ;
        RECT 1755.000 2753.165 1755.260 2753.310 ;
        RECT 1755.920 2753.165 1756.180 2753.310 ;
        RECT 1754.990 2752.795 1755.270 2753.165 ;
        RECT 1755.910 2752.795 1756.190 2753.165 ;
        RECT 1755.980 2705.030 1756.120 2752.795 ;
        RECT 1755.920 2704.710 1756.180 2705.030 ;
        RECT 1755.920 2698.250 1756.180 2698.570 ;
        RECT 1755.980 2659.890 1756.120 2698.250 ;
        RECT 1755.520 2659.750 1756.120 2659.890 ;
        RECT 1755.520 2642.810 1755.660 2659.750 ;
        RECT 1754.540 2642.490 1754.800 2642.810 ;
        RECT 1755.460 2642.490 1755.720 2642.810 ;
        RECT 1754.600 2622.320 1754.740 2642.490 ;
        RECT 1754.140 2622.180 1754.740 2622.320 ;
        RECT 1754.140 2553.245 1754.280 2622.180 ;
        RECT 1754.070 2552.875 1754.350 2553.245 ;
        RECT 1754.990 2552.875 1755.270 2553.245 ;
        RECT 1755.060 2525.930 1755.200 2552.875 ;
        RECT 1755.060 2525.790 1755.660 2525.930 ;
        RECT 1755.520 2511.910 1755.660 2525.790 ;
        RECT 1755.000 2511.765 1755.260 2511.910 ;
        RECT 1754.990 2511.395 1755.270 2511.765 ;
        RECT 1755.460 2511.590 1755.720 2511.910 ;
        RECT 1756.370 2511.395 1756.650 2511.765 ;
        RECT 1756.440 2423.170 1756.580 2511.395 ;
        RECT 1754.540 2422.850 1754.800 2423.170 ;
        RECT 1756.380 2422.850 1756.640 2423.170 ;
        RECT 1754.600 2343.270 1754.740 2422.850 ;
        RECT 1754.540 2342.950 1754.800 2343.270 ;
        RECT 1754.540 2284.020 1754.800 2284.110 ;
        RECT 1754.140 2283.880 1754.800 2284.020 ;
        RECT 1754.140 2264.810 1754.280 2283.880 ;
        RECT 1754.540 2283.790 1754.800 2283.880 ;
        RECT 1754.140 2264.670 1754.740 2264.810 ;
        RECT 1754.600 2261.410 1754.740 2264.670 ;
        RECT 1754.140 2261.270 1754.740 2261.410 ;
        RECT 1754.140 2239.650 1754.280 2261.270 ;
        RECT 1754.140 2239.510 1754.740 2239.650 ;
        RECT 1754.600 2238.290 1754.740 2239.510 ;
        RECT 1754.140 2238.150 1754.740 2238.290 ;
        RECT 1754.140 2149.890 1754.280 2238.150 ;
        RECT 1753.220 2149.750 1754.280 2149.890 ;
        RECT 1753.220 2136.970 1753.360 2149.750 ;
        RECT 1753.220 2136.830 1753.820 2136.970 ;
        RECT 1753.680 2100.930 1753.820 2136.830 ;
        RECT 1753.680 2100.790 1754.280 2100.930 ;
        RECT 1754.140 2044.490 1754.280 2100.790 ;
        RECT 1754.140 2044.410 1754.740 2044.490 ;
        RECT 1754.140 2044.350 1754.800 2044.410 ;
        RECT 1754.540 2044.090 1754.800 2044.350 ;
        RECT 1754.540 2035.650 1754.800 2035.910 ;
        RECT 1754.140 2035.590 1754.800 2035.650 ;
        RECT 1754.140 2035.510 1754.740 2035.590 ;
        RECT 1754.140 2028.170 1754.280 2035.510 ;
        RECT 1752.300 2028.030 1754.280 2028.170 ;
        RECT 1752.300 1993.490 1752.440 2028.030 ;
        RECT 1752.300 1993.350 1753.820 1993.490 ;
        RECT 1753.680 1949.290 1753.820 1993.350 ;
        RECT 1753.220 1949.150 1753.820 1949.290 ;
        RECT 1753.220 1945.210 1753.360 1949.150 ;
        RECT 1753.220 1945.070 1754.280 1945.210 ;
        RECT 1754.140 1894.210 1754.280 1945.070 ;
        RECT 1753.220 1894.070 1754.280 1894.210 ;
        RECT 1753.220 1807.850 1753.360 1894.070 ;
        RECT 1753.220 1807.710 1755.200 1807.850 ;
        RECT 1755.060 1759.490 1755.200 1807.710 ;
        RECT 1757.750 1759.995 1758.030 1760.365 ;
        RECT 1757.820 1759.490 1757.960 1759.995 ;
        RECT 1755.000 1759.170 1755.260 1759.490 ;
        RECT 1757.760 1759.170 1758.020 1759.490 ;
      LAYER via2 ;
        RECT 1753.610 3132.280 1753.890 3132.560 ;
        RECT 1754.530 3132.280 1754.810 3132.560 ;
        RECT 1754.990 2897.680 1755.270 2897.960 ;
        RECT 1755.910 2897.680 1756.190 2897.960 ;
        RECT 1754.990 2849.400 1755.270 2849.680 ;
        RECT 1755.910 2849.400 1756.190 2849.680 ;
        RECT 1754.990 2801.120 1755.270 2801.400 ;
        RECT 1755.910 2801.120 1756.190 2801.400 ;
        RECT 1754.990 2752.840 1755.270 2753.120 ;
        RECT 1755.910 2752.840 1756.190 2753.120 ;
        RECT 1754.070 2552.920 1754.350 2553.200 ;
        RECT 1754.990 2552.920 1755.270 2553.200 ;
        RECT 1754.990 2511.440 1755.270 2511.720 ;
        RECT 1756.370 2511.440 1756.650 2511.720 ;
        RECT 1757.750 1760.040 1758.030 1760.320 ;
      LAYER met3 ;
        RECT 1753.585 3132.570 1753.915 3132.585 ;
        RECT 1754.505 3132.570 1754.835 3132.585 ;
        RECT 1753.585 3132.270 1754.835 3132.570 ;
        RECT 1753.585 3132.255 1753.915 3132.270 ;
        RECT 1754.505 3132.255 1754.835 3132.270 ;
        RECT 1754.965 2897.970 1755.295 2897.985 ;
        RECT 1755.885 2897.970 1756.215 2897.985 ;
        RECT 1754.965 2897.670 1756.215 2897.970 ;
        RECT 1754.965 2897.655 1755.295 2897.670 ;
        RECT 1755.885 2897.655 1756.215 2897.670 ;
        RECT 1754.965 2849.690 1755.295 2849.705 ;
        RECT 1755.885 2849.690 1756.215 2849.705 ;
        RECT 1754.965 2849.390 1756.215 2849.690 ;
        RECT 1754.965 2849.375 1755.295 2849.390 ;
        RECT 1755.885 2849.375 1756.215 2849.390 ;
        RECT 1754.965 2801.410 1755.295 2801.425 ;
        RECT 1755.885 2801.410 1756.215 2801.425 ;
        RECT 1754.965 2801.110 1756.215 2801.410 ;
        RECT 1754.965 2801.095 1755.295 2801.110 ;
        RECT 1755.885 2801.095 1756.215 2801.110 ;
        RECT 1754.965 2753.130 1755.295 2753.145 ;
        RECT 1755.885 2753.130 1756.215 2753.145 ;
        RECT 1754.965 2752.830 1756.215 2753.130 ;
        RECT 1754.965 2752.815 1755.295 2752.830 ;
        RECT 1755.885 2752.815 1756.215 2752.830 ;
        RECT 1754.045 2553.210 1754.375 2553.225 ;
        RECT 1754.965 2553.210 1755.295 2553.225 ;
        RECT 1754.045 2552.910 1755.295 2553.210 ;
        RECT 1754.045 2552.895 1754.375 2552.910 ;
        RECT 1754.965 2552.895 1755.295 2552.910 ;
        RECT 1754.965 2511.730 1755.295 2511.745 ;
        RECT 1756.345 2511.730 1756.675 2511.745 ;
        RECT 1754.965 2511.430 1756.675 2511.730 ;
        RECT 1754.965 2511.415 1755.295 2511.430 ;
        RECT 1756.345 2511.415 1756.675 2511.430 ;
        RECT 1757.725 1760.330 1758.055 1760.345 ;
        RECT 1757.510 1760.015 1758.055 1760.330 ;
        RECT 1757.510 1758.975 1757.810 1760.015 ;
        RECT 1755.835 1758.375 1759.835 1758.975 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 40.625 3429.325 40.795 3477.435 ;
        RECT 40.165 2898.585 40.335 2946.355 ;
        RECT 40.165 2704.785 40.335 2752.895 ;
        RECT 39.705 2221.985 39.875 2270.095 ;
        RECT 40.625 2077.145 40.795 2090.915 ;
        RECT 40.625 1980.245 40.795 2028.355 ;
      LAYER mcon ;
        RECT 40.625 3477.265 40.795 3477.435 ;
        RECT 40.165 2946.185 40.335 2946.355 ;
        RECT 40.165 2752.725 40.335 2752.895 ;
        RECT 39.705 2269.925 39.875 2270.095 ;
        RECT 40.625 2090.745 40.795 2090.915 ;
        RECT 40.625 2028.185 40.795 2028.355 ;
      LAYER met1 ;
        RECT 40.090 3491.360 40.410 3491.420 ;
        RECT 41.010 3491.360 41.330 3491.420 ;
        RECT 40.090 3491.220 41.330 3491.360 ;
        RECT 40.090 3491.160 40.410 3491.220 ;
        RECT 41.010 3491.160 41.330 3491.220 ;
        RECT 40.565 3477.420 40.855 3477.465 ;
        RECT 41.010 3477.420 41.330 3477.480 ;
        RECT 40.565 3477.280 41.330 3477.420 ;
        RECT 40.565 3477.235 40.855 3477.280 ;
        RECT 41.010 3477.220 41.330 3477.280 ;
        RECT 40.550 3429.480 40.870 3429.540 ;
        RECT 40.355 3429.340 40.870 3429.480 ;
        RECT 40.550 3429.280 40.870 3429.340 ;
        RECT 40.550 3395.140 40.870 3395.200 ;
        RECT 40.180 3395.000 40.870 3395.140 ;
        RECT 40.180 3394.860 40.320 3395.000 ;
        RECT 40.550 3394.940 40.870 3395.000 ;
        RECT 40.090 3394.600 40.410 3394.860 ;
        RECT 40.090 3367.600 40.410 3367.660 ;
        RECT 41.010 3367.600 41.330 3367.660 ;
        RECT 40.090 3367.460 41.330 3367.600 ;
        RECT 40.090 3367.400 40.410 3367.460 ;
        RECT 41.010 3367.400 41.330 3367.460 ;
        RECT 40.090 3270.700 40.410 3270.760 ;
        RECT 41.010 3270.700 41.330 3270.760 ;
        RECT 40.090 3270.560 41.330 3270.700 ;
        RECT 40.090 3270.500 40.410 3270.560 ;
        RECT 41.010 3270.500 41.330 3270.560 ;
        RECT 40.090 3174.140 40.410 3174.200 ;
        RECT 41.010 3174.140 41.330 3174.200 ;
        RECT 40.090 3174.000 41.330 3174.140 ;
        RECT 40.090 3173.940 40.410 3174.000 ;
        RECT 41.010 3173.940 41.330 3174.000 ;
        RECT 40.090 3077.580 40.410 3077.640 ;
        RECT 41.010 3077.580 41.330 3077.640 ;
        RECT 40.090 3077.440 41.330 3077.580 ;
        RECT 40.090 3077.380 40.410 3077.440 ;
        RECT 41.010 3077.380 41.330 3077.440 ;
        RECT 40.090 2981.020 40.410 2981.080 ;
        RECT 41.010 2981.020 41.330 2981.080 ;
        RECT 40.090 2980.880 41.330 2981.020 ;
        RECT 40.090 2980.820 40.410 2980.880 ;
        RECT 41.010 2980.820 41.330 2980.880 ;
        RECT 40.090 2946.340 40.410 2946.400 ;
        RECT 39.895 2946.200 40.410 2946.340 ;
        RECT 40.090 2946.140 40.410 2946.200 ;
        RECT 40.090 2898.740 40.410 2898.800 ;
        RECT 39.895 2898.600 40.410 2898.740 ;
        RECT 40.090 2898.540 40.410 2898.600 ;
        RECT 39.630 2898.060 39.950 2898.120 ;
        RECT 40.550 2898.060 40.870 2898.120 ;
        RECT 39.630 2897.920 40.870 2898.060 ;
        RECT 39.630 2897.860 39.950 2897.920 ;
        RECT 40.550 2897.860 40.870 2897.920 ;
        RECT 39.630 2814.760 39.950 2814.820 ;
        RECT 40.550 2814.760 40.870 2814.820 ;
        RECT 39.630 2814.620 40.870 2814.760 ;
        RECT 39.630 2814.560 39.950 2814.620 ;
        RECT 40.550 2814.560 40.870 2814.620 ;
        RECT 40.090 2752.880 40.410 2752.940 ;
        RECT 39.895 2752.740 40.410 2752.880 ;
        RECT 40.090 2752.680 40.410 2752.740 ;
        RECT 40.105 2704.940 40.395 2704.985 ;
        RECT 41.010 2704.940 41.330 2705.000 ;
        RECT 40.105 2704.800 41.330 2704.940 ;
        RECT 40.105 2704.755 40.395 2704.800 ;
        RECT 41.010 2704.740 41.330 2704.800 ;
        RECT 41.010 2608.380 41.330 2608.440 ;
        RECT 41.930 2608.380 42.250 2608.440 ;
        RECT 41.010 2608.240 42.250 2608.380 ;
        RECT 41.010 2608.180 41.330 2608.240 ;
        RECT 41.930 2608.180 42.250 2608.240 ;
        RECT 41.010 2511.820 41.330 2511.880 ;
        RECT 41.930 2511.820 42.250 2511.880 ;
        RECT 41.010 2511.680 42.250 2511.820 ;
        RECT 41.010 2511.620 41.330 2511.680 ;
        RECT 41.930 2511.620 42.250 2511.680 ;
        RECT 40.090 2429.000 40.410 2429.260 ;
        RECT 40.180 2428.520 40.320 2429.000 ;
        RECT 40.550 2428.520 40.870 2428.580 ;
        RECT 40.180 2428.380 40.870 2428.520 ;
        RECT 40.550 2428.320 40.870 2428.380 ;
        RECT 39.170 2414.920 39.490 2414.980 ;
        RECT 40.550 2414.920 40.870 2414.980 ;
        RECT 39.170 2414.780 40.870 2414.920 ;
        RECT 39.170 2414.720 39.490 2414.780 ;
        RECT 40.550 2414.720 40.870 2414.780 ;
        RECT 40.090 2332.100 40.410 2332.360 ;
        RECT 40.180 2331.960 40.320 2332.100 ;
        RECT 41.010 2331.960 41.330 2332.020 ;
        RECT 40.180 2331.820 41.330 2331.960 ;
        RECT 41.010 2331.760 41.330 2331.820 ;
        RECT 39.645 2270.080 39.935 2270.125 ;
        RECT 40.090 2270.080 40.410 2270.140 ;
        RECT 39.645 2269.940 40.410 2270.080 ;
        RECT 39.645 2269.895 39.935 2269.940 ;
        RECT 40.090 2269.880 40.410 2269.940 ;
        RECT 39.630 2222.140 39.950 2222.200 ;
        RECT 39.435 2222.000 39.950 2222.140 ;
        RECT 39.630 2221.940 39.950 2222.000 ;
        RECT 40.550 2138.980 40.870 2139.240 ;
        RECT 40.640 2138.840 40.780 2138.980 ;
        RECT 41.010 2138.840 41.330 2138.900 ;
        RECT 40.640 2138.700 41.330 2138.840 ;
        RECT 41.010 2138.640 41.330 2138.700 ;
        RECT 40.550 2090.900 40.870 2090.960 ;
        RECT 40.355 2090.760 40.870 2090.900 ;
        RECT 40.550 2090.700 40.870 2090.760 ;
        RECT 40.550 2077.300 40.870 2077.360 ;
        RECT 40.355 2077.160 40.870 2077.300 ;
        RECT 40.550 2077.100 40.870 2077.160 ;
        RECT 40.550 2042.420 40.870 2042.680 ;
        RECT 40.640 2041.940 40.780 2042.420 ;
        RECT 41.010 2041.940 41.330 2042.000 ;
        RECT 40.640 2041.800 41.330 2041.940 ;
        RECT 41.010 2041.740 41.330 2041.800 ;
        RECT 40.565 2028.340 40.855 2028.385 ;
        RECT 41.010 2028.340 41.330 2028.400 ;
        RECT 40.565 2028.200 41.330 2028.340 ;
        RECT 40.565 2028.155 40.855 2028.200 ;
        RECT 41.010 2028.140 41.330 2028.200 ;
        RECT 40.550 1980.400 40.870 1980.460 ;
        RECT 40.355 1980.260 40.870 1980.400 ;
        RECT 40.550 1980.200 40.870 1980.260 ;
        RECT 40.550 1945.860 40.870 1946.120 ;
        RECT 40.640 1945.440 40.780 1945.860 ;
        RECT 40.550 1945.180 40.870 1945.440 ;
        RECT 40.550 1897.920 40.870 1898.180 ;
        RECT 40.640 1897.500 40.780 1897.920 ;
        RECT 40.550 1897.240 40.870 1897.500 ;
        RECT 39.630 1821.960 39.950 1822.020 ;
        RECT 41.010 1821.960 41.330 1822.020 ;
        RECT 39.630 1821.820 41.330 1821.960 ;
        RECT 39.630 1821.760 39.950 1821.820 ;
        RECT 41.010 1821.760 41.330 1821.820 ;
        RECT 39.630 1773.000 39.950 1773.060 ;
        RECT 41.010 1773.000 41.330 1773.060 ;
        RECT 39.630 1772.860 41.330 1773.000 ;
        RECT 39.630 1772.800 39.950 1772.860 ;
        RECT 41.010 1772.800 41.330 1772.860 ;
        RECT 39.630 1725.400 39.950 1725.460 ;
        RECT 41.010 1725.400 41.330 1725.460 ;
        RECT 39.630 1725.260 41.330 1725.400 ;
        RECT 39.630 1725.200 39.950 1725.260 ;
        RECT 41.010 1725.200 41.330 1725.260 ;
        RECT 39.630 1676.440 39.950 1676.500 ;
        RECT 41.010 1676.440 41.330 1676.500 ;
        RECT 39.630 1676.300 41.330 1676.440 ;
        RECT 39.630 1676.240 39.950 1676.300 ;
        RECT 41.010 1676.240 41.330 1676.300 ;
        RECT 39.630 1628.500 39.950 1628.560 ;
        RECT 41.010 1628.500 41.330 1628.560 ;
        RECT 39.630 1628.360 41.330 1628.500 ;
        RECT 39.630 1628.300 39.950 1628.360 ;
        RECT 41.010 1628.300 41.330 1628.360 ;
        RECT 39.630 1579.880 39.950 1579.940 ;
        RECT 41.010 1579.880 41.330 1579.940 ;
        RECT 39.630 1579.740 41.330 1579.880 ;
        RECT 39.630 1579.680 39.950 1579.740 ;
        RECT 41.010 1579.680 41.330 1579.740 ;
        RECT 39.630 1531.940 39.950 1532.000 ;
        RECT 41.010 1531.940 41.330 1532.000 ;
        RECT 39.630 1531.800 41.330 1531.940 ;
        RECT 39.630 1531.740 39.950 1531.800 ;
        RECT 41.010 1531.740 41.330 1531.800 ;
        RECT 39.630 1483.320 39.950 1483.380 ;
        RECT 41.010 1483.320 41.330 1483.380 ;
        RECT 39.630 1483.180 41.330 1483.320 ;
        RECT 39.630 1483.120 39.950 1483.180 ;
        RECT 41.010 1483.120 41.330 1483.180 ;
        RECT 39.630 1435.380 39.950 1435.440 ;
        RECT 41.010 1435.380 41.330 1435.440 ;
        RECT 39.630 1435.240 41.330 1435.380 ;
        RECT 39.630 1435.180 39.950 1435.240 ;
        RECT 41.010 1435.180 41.330 1435.240 ;
        RECT 41.010 1393.560 41.330 1393.620 ;
        RECT 684.550 1393.560 684.870 1393.620 ;
        RECT 41.010 1393.420 684.870 1393.560 ;
        RECT 41.010 1393.360 41.330 1393.420 ;
        RECT 684.550 1393.360 684.870 1393.420 ;
      LAYER via ;
        RECT 40.120 3491.160 40.380 3491.420 ;
        RECT 41.040 3491.160 41.300 3491.420 ;
        RECT 41.040 3477.220 41.300 3477.480 ;
        RECT 40.580 3429.280 40.840 3429.540 ;
        RECT 40.580 3394.940 40.840 3395.200 ;
        RECT 40.120 3394.600 40.380 3394.860 ;
        RECT 40.120 3367.400 40.380 3367.660 ;
        RECT 41.040 3367.400 41.300 3367.660 ;
        RECT 40.120 3270.500 40.380 3270.760 ;
        RECT 41.040 3270.500 41.300 3270.760 ;
        RECT 40.120 3173.940 40.380 3174.200 ;
        RECT 41.040 3173.940 41.300 3174.200 ;
        RECT 40.120 3077.380 40.380 3077.640 ;
        RECT 41.040 3077.380 41.300 3077.640 ;
        RECT 40.120 2980.820 40.380 2981.080 ;
        RECT 41.040 2980.820 41.300 2981.080 ;
        RECT 40.120 2946.140 40.380 2946.400 ;
        RECT 40.120 2898.540 40.380 2898.800 ;
        RECT 39.660 2897.860 39.920 2898.120 ;
        RECT 40.580 2897.860 40.840 2898.120 ;
        RECT 39.660 2814.560 39.920 2814.820 ;
        RECT 40.580 2814.560 40.840 2814.820 ;
        RECT 40.120 2752.680 40.380 2752.940 ;
        RECT 41.040 2704.740 41.300 2705.000 ;
        RECT 41.040 2608.180 41.300 2608.440 ;
        RECT 41.960 2608.180 42.220 2608.440 ;
        RECT 41.040 2511.620 41.300 2511.880 ;
        RECT 41.960 2511.620 42.220 2511.880 ;
        RECT 40.120 2429.000 40.380 2429.260 ;
        RECT 40.580 2428.320 40.840 2428.580 ;
        RECT 39.200 2414.720 39.460 2414.980 ;
        RECT 40.580 2414.720 40.840 2414.980 ;
        RECT 40.120 2332.100 40.380 2332.360 ;
        RECT 41.040 2331.760 41.300 2332.020 ;
        RECT 40.120 2269.880 40.380 2270.140 ;
        RECT 39.660 2221.940 39.920 2222.200 ;
        RECT 40.580 2138.980 40.840 2139.240 ;
        RECT 41.040 2138.640 41.300 2138.900 ;
        RECT 40.580 2090.700 40.840 2090.960 ;
        RECT 40.580 2077.100 40.840 2077.360 ;
        RECT 40.580 2042.420 40.840 2042.680 ;
        RECT 41.040 2041.740 41.300 2042.000 ;
        RECT 41.040 2028.140 41.300 2028.400 ;
        RECT 40.580 1980.200 40.840 1980.460 ;
        RECT 40.580 1945.860 40.840 1946.120 ;
        RECT 40.580 1945.180 40.840 1945.440 ;
        RECT 40.580 1897.920 40.840 1898.180 ;
        RECT 40.580 1897.240 40.840 1897.500 ;
        RECT 39.660 1821.760 39.920 1822.020 ;
        RECT 41.040 1821.760 41.300 1822.020 ;
        RECT 39.660 1772.800 39.920 1773.060 ;
        RECT 41.040 1772.800 41.300 1773.060 ;
        RECT 39.660 1725.200 39.920 1725.460 ;
        RECT 41.040 1725.200 41.300 1725.460 ;
        RECT 39.660 1676.240 39.920 1676.500 ;
        RECT 41.040 1676.240 41.300 1676.500 ;
        RECT 39.660 1628.300 39.920 1628.560 ;
        RECT 41.040 1628.300 41.300 1628.560 ;
        RECT 39.660 1579.680 39.920 1579.940 ;
        RECT 41.040 1579.680 41.300 1579.940 ;
        RECT 39.660 1531.740 39.920 1532.000 ;
        RECT 41.040 1531.740 41.300 1532.000 ;
        RECT 39.660 1483.120 39.920 1483.380 ;
        RECT 41.040 1483.120 41.300 1483.380 ;
        RECT 39.660 1435.180 39.920 1435.440 ;
        RECT 41.040 1435.180 41.300 1435.440 ;
        RECT 41.040 1393.360 41.300 1393.620 ;
        RECT 684.580 1393.360 684.840 1393.620 ;
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
        RECT 40.640 3517.370 40.780 3517.600 ;
        RECT 40.180 3517.230 40.780 3517.370 ;
        RECT 40.180 3491.450 40.320 3517.230 ;
        RECT 40.120 3491.130 40.380 3491.450 ;
        RECT 41.040 3491.130 41.300 3491.450 ;
        RECT 41.100 3477.510 41.240 3491.130 ;
        RECT 41.040 3477.190 41.300 3477.510 ;
        RECT 40.580 3429.250 40.840 3429.570 ;
        RECT 40.640 3395.230 40.780 3429.250 ;
        RECT 40.580 3394.910 40.840 3395.230 ;
        RECT 40.120 3394.570 40.380 3394.890 ;
        RECT 40.180 3367.690 40.320 3394.570 ;
        RECT 40.120 3367.370 40.380 3367.690 ;
        RECT 41.040 3367.370 41.300 3367.690 ;
        RECT 41.100 3318.810 41.240 3367.370 ;
        RECT 40.180 3318.670 41.240 3318.810 ;
        RECT 40.180 3270.790 40.320 3318.670 ;
        RECT 40.120 3270.470 40.380 3270.790 ;
        RECT 41.040 3270.470 41.300 3270.790 ;
        RECT 41.100 3222.250 41.240 3270.470 ;
        RECT 40.180 3222.110 41.240 3222.250 ;
        RECT 40.180 3174.230 40.320 3222.110 ;
        RECT 40.120 3173.910 40.380 3174.230 ;
        RECT 41.040 3173.910 41.300 3174.230 ;
        RECT 41.100 3125.690 41.240 3173.910 ;
        RECT 40.180 3125.550 41.240 3125.690 ;
        RECT 40.180 3077.670 40.320 3125.550 ;
        RECT 40.120 3077.350 40.380 3077.670 ;
        RECT 41.040 3077.350 41.300 3077.670 ;
        RECT 41.100 3029.130 41.240 3077.350 ;
        RECT 40.180 3028.990 41.240 3029.130 ;
        RECT 40.180 2981.110 40.320 3028.990 ;
        RECT 40.120 2980.790 40.380 2981.110 ;
        RECT 41.040 2980.850 41.300 2981.110 ;
        RECT 40.640 2980.790 41.300 2980.850 ;
        RECT 40.640 2980.710 41.240 2980.790 ;
        RECT 40.640 2959.770 40.780 2980.710 ;
        RECT 40.180 2959.630 40.780 2959.770 ;
        RECT 40.180 2946.430 40.320 2959.630 ;
        RECT 40.120 2946.110 40.380 2946.430 ;
        RECT 40.120 2898.570 40.380 2898.830 ;
        RECT 39.720 2898.510 40.380 2898.570 ;
        RECT 39.720 2898.430 40.320 2898.510 ;
        RECT 39.720 2898.150 39.860 2898.430 ;
        RECT 39.660 2897.830 39.920 2898.150 ;
        RECT 40.580 2897.830 40.840 2898.150 ;
        RECT 40.640 2814.850 40.780 2897.830 ;
        RECT 39.660 2814.530 39.920 2814.850 ;
        RECT 40.580 2814.530 40.840 2814.850 ;
        RECT 39.720 2766.650 39.860 2814.530 ;
        RECT 39.720 2766.510 40.320 2766.650 ;
        RECT 40.180 2752.970 40.320 2766.510 ;
        RECT 40.120 2752.650 40.380 2752.970 ;
        RECT 41.040 2704.710 41.300 2705.030 ;
        RECT 41.100 2670.090 41.240 2704.710 ;
        RECT 40.640 2669.950 41.240 2670.090 ;
        RECT 40.640 2656.605 40.780 2669.950 ;
        RECT 40.570 2656.235 40.850 2656.605 ;
        RECT 41.950 2656.235 42.230 2656.605 ;
        RECT 42.020 2608.470 42.160 2656.235 ;
        RECT 41.040 2608.150 41.300 2608.470 ;
        RECT 41.960 2608.150 42.220 2608.470 ;
        RECT 41.100 2573.530 41.240 2608.150 ;
        RECT 40.640 2573.390 41.240 2573.530 ;
        RECT 40.640 2560.045 40.780 2573.390 ;
        RECT 40.570 2559.675 40.850 2560.045 ;
        RECT 41.950 2559.675 42.230 2560.045 ;
        RECT 42.020 2511.910 42.160 2559.675 ;
        RECT 41.040 2511.590 41.300 2511.910 ;
        RECT 41.960 2511.590 42.220 2511.910 ;
        RECT 41.100 2476.970 41.240 2511.590 ;
        RECT 40.180 2476.830 41.240 2476.970 ;
        RECT 40.180 2429.290 40.320 2476.830 ;
        RECT 40.120 2428.970 40.380 2429.290 ;
        RECT 40.580 2428.290 40.840 2428.610 ;
        RECT 40.640 2415.010 40.780 2428.290 ;
        RECT 39.200 2414.690 39.460 2415.010 ;
        RECT 40.580 2414.690 40.840 2415.010 ;
        RECT 39.260 2366.925 39.400 2414.690 ;
        RECT 39.190 2366.555 39.470 2366.925 ;
        RECT 40.110 2366.555 40.390 2366.925 ;
        RECT 40.180 2332.390 40.320 2366.555 ;
        RECT 40.120 2332.070 40.380 2332.390 ;
        RECT 41.040 2331.730 41.300 2332.050 ;
        RECT 41.100 2283.850 41.240 2331.730 ;
        RECT 40.180 2283.710 41.240 2283.850 ;
        RECT 40.180 2270.170 40.320 2283.710 ;
        RECT 40.120 2269.850 40.380 2270.170 ;
        RECT 39.660 2221.910 39.920 2222.230 ;
        RECT 39.720 2187.290 39.860 2221.910 ;
        RECT 39.720 2187.150 40.780 2187.290 ;
        RECT 40.640 2139.270 40.780 2187.150 ;
        RECT 40.580 2138.950 40.840 2139.270 ;
        RECT 41.040 2138.610 41.300 2138.930 ;
        RECT 41.100 2125.240 41.240 2138.610 ;
        RECT 40.640 2125.100 41.240 2125.240 ;
        RECT 40.640 2090.990 40.780 2125.100 ;
        RECT 40.580 2090.670 40.840 2090.990 ;
        RECT 40.580 2077.070 40.840 2077.390 ;
        RECT 40.640 2042.710 40.780 2077.070 ;
        RECT 40.580 2042.390 40.840 2042.710 ;
        RECT 41.040 2041.710 41.300 2042.030 ;
        RECT 41.100 2028.430 41.240 2041.710 ;
        RECT 41.040 2028.110 41.300 2028.430 ;
        RECT 40.580 1980.170 40.840 1980.490 ;
        RECT 40.640 1946.150 40.780 1980.170 ;
        RECT 40.580 1945.830 40.840 1946.150 ;
        RECT 40.580 1945.150 40.840 1945.470 ;
        RECT 40.640 1898.210 40.780 1945.150 ;
        RECT 40.580 1897.890 40.840 1898.210 ;
        RECT 40.580 1897.210 40.840 1897.530 ;
        RECT 40.640 1849.330 40.780 1897.210 ;
        RECT 39.720 1849.190 40.780 1849.330 ;
        RECT 39.720 1822.050 39.860 1849.190 ;
        RECT 39.660 1821.730 39.920 1822.050 ;
        RECT 41.040 1821.730 41.300 1822.050 ;
        RECT 41.100 1773.090 41.240 1821.730 ;
        RECT 39.660 1772.770 39.920 1773.090 ;
        RECT 41.040 1772.770 41.300 1773.090 ;
        RECT 39.720 1725.490 39.860 1772.770 ;
        RECT 39.660 1725.170 39.920 1725.490 ;
        RECT 41.040 1725.170 41.300 1725.490 ;
        RECT 41.100 1676.530 41.240 1725.170 ;
        RECT 39.660 1676.210 39.920 1676.530 ;
        RECT 41.040 1676.210 41.300 1676.530 ;
        RECT 39.720 1628.590 39.860 1676.210 ;
        RECT 39.660 1628.270 39.920 1628.590 ;
        RECT 41.040 1628.270 41.300 1628.590 ;
        RECT 41.100 1579.970 41.240 1628.270 ;
        RECT 39.660 1579.650 39.920 1579.970 ;
        RECT 41.040 1579.650 41.300 1579.970 ;
        RECT 39.720 1532.030 39.860 1579.650 ;
        RECT 39.660 1531.710 39.920 1532.030 ;
        RECT 41.040 1531.710 41.300 1532.030 ;
        RECT 41.100 1483.410 41.240 1531.710 ;
        RECT 39.660 1483.090 39.920 1483.410 ;
        RECT 41.040 1483.090 41.300 1483.410 ;
        RECT 39.720 1435.470 39.860 1483.090 ;
        RECT 39.660 1435.150 39.920 1435.470 ;
        RECT 41.040 1435.150 41.300 1435.470 ;
        RECT 41.100 1393.650 41.240 1435.150 ;
        RECT 41.040 1393.330 41.300 1393.650 ;
        RECT 684.580 1393.330 684.840 1393.650 ;
        RECT 684.640 1387.725 684.780 1393.330 ;
        RECT 684.570 1387.355 684.850 1387.725 ;
      LAYER via2 ;
        RECT 40.570 2656.280 40.850 2656.560 ;
        RECT 41.950 2656.280 42.230 2656.560 ;
        RECT 40.570 2559.720 40.850 2560.000 ;
        RECT 41.950 2559.720 42.230 2560.000 ;
        RECT 39.190 2366.600 39.470 2366.880 ;
        RECT 40.110 2366.600 40.390 2366.880 ;
        RECT 684.570 1387.400 684.850 1387.680 ;
      LAYER met3 ;
        RECT 40.545 2656.570 40.875 2656.585 ;
        RECT 41.925 2656.570 42.255 2656.585 ;
        RECT 40.545 2656.270 42.255 2656.570 ;
        RECT 40.545 2656.255 40.875 2656.270 ;
        RECT 41.925 2656.255 42.255 2656.270 ;
        RECT 40.545 2560.010 40.875 2560.025 ;
        RECT 41.925 2560.010 42.255 2560.025 ;
        RECT 40.545 2559.710 42.255 2560.010 ;
        RECT 40.545 2559.695 40.875 2559.710 ;
        RECT 41.925 2559.695 42.255 2559.710 ;
        RECT 39.165 2366.890 39.495 2366.905 ;
        RECT 40.085 2366.890 40.415 2366.905 ;
        RECT 39.165 2366.590 40.415 2366.890 ;
        RECT 39.165 2366.575 39.495 2366.590 ;
        RECT 40.085 2366.575 40.415 2366.590 ;
        RECT 684.545 1387.690 684.875 1387.705 ;
        RECT 715.810 1387.690 719.810 1387.695 ;
        RECT 684.545 1387.390 719.810 1387.690 ;
        RECT 684.545 1387.375 684.875 1387.390 ;
        RECT 715.810 1387.095 719.810 1387.390 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 20.310 3263.900 20.630 3263.960 ;
        RECT 25.830 3263.900 26.150 3263.960 ;
        RECT 20.310 3263.760 26.150 3263.900 ;
        RECT 20.310 3263.700 20.630 3263.760 ;
        RECT 25.830 3263.700 26.150 3263.760 ;
        RECT 25.830 1793.740 26.150 1793.800 ;
        RECT 705.710 1793.740 706.030 1793.800 ;
        RECT 25.830 1793.600 706.030 1793.740 ;
        RECT 25.830 1793.540 26.150 1793.600 ;
        RECT 705.710 1793.540 706.030 1793.600 ;
      LAYER via ;
        RECT 20.340 3263.700 20.600 3263.960 ;
        RECT 25.860 3263.700 26.120 3263.960 ;
        RECT 25.860 1793.540 26.120 1793.800 ;
        RECT 705.740 1793.540 706.000 1793.800 ;
      LAYER met2 ;
        RECT 20.330 3267.555 20.610 3267.925 ;
        RECT 20.400 3263.990 20.540 3267.555 ;
        RECT 20.340 3263.670 20.600 3263.990 ;
        RECT 25.860 3263.670 26.120 3263.990 ;
        RECT 25.920 1793.830 26.060 3263.670 ;
        RECT 25.860 1793.510 26.120 1793.830 ;
        RECT 705.740 1793.510 706.000 1793.830 ;
        RECT 705.800 1788.925 705.940 1793.510 ;
        RECT 705.730 1788.555 706.010 1788.925 ;
      LAYER via2 ;
        RECT 20.330 3267.600 20.610 3267.880 ;
        RECT 705.730 1788.600 706.010 1788.880 ;
      LAYER met3 ;
        RECT -4.800 3267.890 2.400 3268.340 ;
        RECT 20.305 3267.890 20.635 3267.905 ;
        RECT -4.800 3267.590 20.635 3267.890 ;
        RECT -4.800 3267.140 2.400 3267.590 ;
        RECT 20.305 3267.575 20.635 3267.590 ;
        RECT 705.705 1788.890 706.035 1788.905 ;
        RECT 715.810 1788.890 719.810 1788.895 ;
        RECT 705.705 1788.590 719.810 1788.890 ;
        RECT 705.705 1788.575 706.035 1788.590 ;
        RECT 715.810 1788.295 719.810 1788.590 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.170 2974.220 16.490 2974.280 ;
        RECT 700.190 2974.220 700.510 2974.280 ;
        RECT 16.170 2974.080 700.510 2974.220 ;
        RECT 16.170 2974.020 16.490 2974.080 ;
        RECT 700.190 2974.020 700.510 2974.080 ;
        RECT 700.190 1322.160 700.510 1322.220 ;
        RECT 1493.230 1322.160 1493.550 1322.220 ;
        RECT 700.190 1322.020 1493.550 1322.160 ;
        RECT 700.190 1321.960 700.510 1322.020 ;
        RECT 1493.230 1321.960 1493.550 1322.020 ;
      LAYER via ;
        RECT 16.200 2974.020 16.460 2974.280 ;
        RECT 700.220 2974.020 700.480 2974.280 ;
        RECT 700.220 1321.960 700.480 1322.220 ;
        RECT 1493.260 1321.960 1493.520 1322.220 ;
      LAYER met2 ;
        RECT 16.190 2979.915 16.470 2980.285 ;
        RECT 16.260 2974.310 16.400 2979.915 ;
        RECT 16.200 2973.990 16.460 2974.310 ;
        RECT 700.220 2973.990 700.480 2974.310 ;
        RECT 700.280 1393.845 700.420 2973.990 ;
        RECT 700.210 1393.475 700.490 1393.845 ;
        RECT 700.210 1392.115 700.490 1392.485 ;
        RECT 700.280 1322.250 700.420 1392.115 ;
        RECT 1493.300 1323.135 1493.580 1327.135 ;
        RECT 1493.320 1322.250 1493.460 1323.135 ;
        RECT 700.220 1321.930 700.480 1322.250 ;
        RECT 1493.260 1321.930 1493.520 1322.250 ;
      LAYER via2 ;
        RECT 16.190 2979.960 16.470 2980.240 ;
        RECT 700.210 1393.520 700.490 1393.800 ;
        RECT 700.210 1392.160 700.490 1392.440 ;
      LAYER met3 ;
        RECT -4.800 2980.250 2.400 2980.700 ;
        RECT 16.165 2980.250 16.495 2980.265 ;
        RECT -4.800 2979.950 16.495 2980.250 ;
        RECT -4.800 2979.500 2.400 2979.950 ;
        RECT 16.165 2979.935 16.495 2979.950 ;
        RECT 700.185 1393.810 700.515 1393.825 ;
        RECT 700.185 1393.495 700.730 1393.810 ;
        RECT 700.430 1392.465 700.730 1393.495 ;
        RECT 700.185 1392.150 700.730 1392.465 ;
        RECT 700.185 1392.135 700.515 1392.150 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 2691.340 16.030 2691.400 ;
        RECT 30.890 2691.340 31.210 2691.400 ;
        RECT 15.710 2691.200 31.210 2691.340 ;
        RECT 15.710 2691.140 16.030 2691.200 ;
        RECT 30.890 2691.140 31.210 2691.200 ;
        RECT 30.890 1320.800 31.210 1320.860 ;
        RECT 1336.830 1320.800 1337.150 1320.860 ;
        RECT 30.890 1320.660 1337.150 1320.800 ;
        RECT 30.890 1320.600 31.210 1320.660 ;
        RECT 1336.830 1320.600 1337.150 1320.660 ;
      LAYER via ;
        RECT 15.740 2691.140 16.000 2691.400 ;
        RECT 30.920 2691.140 31.180 2691.400 ;
        RECT 30.920 1320.600 31.180 1320.860 ;
        RECT 1336.860 1320.600 1337.120 1320.860 ;
      LAYER met2 ;
        RECT 15.730 2692.955 16.010 2693.325 ;
        RECT 15.800 2691.430 15.940 2692.955 ;
        RECT 15.740 2691.110 16.000 2691.430 ;
        RECT 30.920 2691.110 31.180 2691.430 ;
        RECT 30.980 1320.890 31.120 2691.110 ;
        RECT 1336.900 1323.135 1337.180 1327.135 ;
        RECT 1336.920 1320.890 1337.060 1323.135 ;
        RECT 30.920 1320.570 31.180 1320.890 ;
        RECT 1336.860 1320.570 1337.120 1320.890 ;
      LAYER via2 ;
        RECT 15.730 2693.000 16.010 2693.280 ;
      LAYER met3 ;
        RECT -4.800 2693.290 2.400 2693.740 ;
        RECT 15.705 2693.290 16.035 2693.305 ;
        RECT -4.800 2692.990 16.035 2693.290 ;
        RECT -4.800 2692.540 2.400 2692.990 ;
        RECT 15.705 2692.975 16.035 2692.990 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 20.310 2401.320 20.630 2401.380 ;
        RECT 1745.310 2401.320 1745.630 2401.380 ;
        RECT 20.310 2401.180 1745.630 2401.320 ;
        RECT 20.310 2401.120 20.630 2401.180 ;
        RECT 1745.310 2401.120 1745.630 2401.180 ;
      LAYER via ;
        RECT 20.340 2401.120 20.600 2401.380 ;
        RECT 1745.340 2401.120 1745.600 2401.380 ;
      LAYER met2 ;
        RECT 20.330 2405.315 20.610 2405.685 ;
        RECT 20.400 2401.410 20.540 2405.315 ;
        RECT 20.340 2401.090 20.600 2401.410 ;
        RECT 1745.340 2401.090 1745.600 2401.410 ;
        RECT 1745.400 2377.880 1745.540 2401.090 ;
        RECT 1745.380 2373.880 1745.660 2377.880 ;
      LAYER via2 ;
        RECT 20.330 2405.360 20.610 2405.640 ;
      LAYER met3 ;
        RECT -4.800 2405.650 2.400 2406.100 ;
        RECT 20.305 2405.650 20.635 2405.665 ;
        RECT -4.800 2405.350 20.635 2405.650 ;
        RECT -4.800 2404.900 2.400 2405.350 ;
        RECT 20.305 2405.335 20.635 2405.350 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 673.050 2383.640 673.370 2383.700 ;
        RECT 1641.350 2383.640 1641.670 2383.700 ;
        RECT 673.050 2383.500 1641.670 2383.640 ;
        RECT 673.050 2383.440 673.370 2383.500 ;
        RECT 1641.350 2383.440 1641.670 2383.500 ;
        RECT 19.850 2124.900 20.170 2124.960 ;
        RECT 673.050 2124.900 673.370 2124.960 ;
        RECT 19.850 2124.760 673.370 2124.900 ;
        RECT 19.850 2124.700 20.170 2124.760 ;
        RECT 673.050 2124.700 673.370 2124.760 ;
      LAYER via ;
        RECT 673.080 2383.440 673.340 2383.700 ;
        RECT 1641.380 2383.440 1641.640 2383.700 ;
        RECT 19.880 2124.700 20.140 2124.960 ;
        RECT 673.080 2124.700 673.340 2124.960 ;
      LAYER met2 ;
        RECT 673.080 2383.410 673.340 2383.730 ;
        RECT 1641.380 2383.410 1641.640 2383.730 ;
        RECT 673.140 2124.990 673.280 2383.410 ;
        RECT 1641.440 2377.880 1641.580 2383.410 ;
        RECT 1641.420 2373.880 1641.700 2377.880 ;
        RECT 19.880 2124.670 20.140 2124.990 ;
        RECT 673.080 2124.670 673.340 2124.990 ;
        RECT 19.940 2118.725 20.080 2124.670 ;
        RECT 19.870 2118.355 20.150 2118.725 ;
      LAYER via2 ;
        RECT 19.870 2118.400 20.150 2118.680 ;
      LAYER met3 ;
        RECT -4.800 2118.690 2.400 2119.140 ;
        RECT 19.845 2118.690 20.175 2118.705 ;
        RECT -4.800 2118.390 20.175 2118.690 ;
        RECT -4.800 2117.940 2.400 2118.390 ;
        RECT 19.845 2118.375 20.175 2118.390 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.170 1319.440 16.490 1319.500 ;
        RECT 1649.630 1319.440 1649.950 1319.500 ;
        RECT 16.170 1319.300 1649.950 1319.440 ;
        RECT 16.170 1319.240 16.490 1319.300 ;
        RECT 1649.630 1319.240 1649.950 1319.300 ;
      LAYER via ;
        RECT 16.200 1319.240 16.460 1319.500 ;
        RECT 1649.660 1319.240 1649.920 1319.500 ;
      LAYER met2 ;
        RECT 16.650 1830.715 16.930 1831.085 ;
        RECT 16.720 1329.130 16.860 1830.715 ;
        RECT 16.260 1328.990 16.860 1329.130 ;
        RECT 16.260 1319.530 16.400 1328.990 ;
        RECT 1649.700 1323.135 1649.980 1327.135 ;
        RECT 1649.720 1319.530 1649.860 1323.135 ;
        RECT 16.200 1319.210 16.460 1319.530 ;
        RECT 1649.660 1319.210 1649.920 1319.530 ;
      LAYER via2 ;
        RECT 16.650 1830.760 16.930 1831.040 ;
      LAYER met3 ;
        RECT -4.800 1831.050 2.400 1831.500 ;
        RECT 16.625 1831.050 16.955 1831.065 ;
        RECT -4.800 1830.750 16.955 1831.050 ;
        RECT -4.800 1830.300 2.400 1830.750 ;
        RECT 16.625 1830.735 16.955 1830.750 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1288.070 2386.360 1288.390 2386.420 ;
        RECT 1790.850 2386.360 1791.170 2386.420 ;
        RECT 1288.070 2386.220 1791.170 2386.360 ;
        RECT 1288.070 2386.160 1288.390 2386.220 ;
        RECT 1790.850 2386.160 1791.170 2386.220 ;
        RECT 1790.850 676.160 1791.170 676.220 ;
        RECT 2900.830 676.160 2901.150 676.220 ;
        RECT 1790.850 676.020 2901.150 676.160 ;
        RECT 1790.850 675.960 1791.170 676.020 ;
        RECT 2900.830 675.960 2901.150 676.020 ;
      LAYER via ;
        RECT 1288.100 2386.160 1288.360 2386.420 ;
        RECT 1790.880 2386.160 1791.140 2386.420 ;
        RECT 1790.880 675.960 1791.140 676.220 ;
        RECT 2900.860 675.960 2901.120 676.220 ;
      LAYER met2 ;
        RECT 1288.100 2386.130 1288.360 2386.450 ;
        RECT 1790.880 2386.130 1791.140 2386.450 ;
        RECT 1288.160 2377.880 1288.300 2386.130 ;
        RECT 1288.140 2373.880 1288.420 2377.880 ;
        RECT 1790.940 676.250 1791.080 2386.130 ;
        RECT 1790.880 675.930 1791.140 676.250 ;
        RECT 2900.860 675.930 2901.120 676.250 ;
        RECT 2900.920 674.405 2901.060 675.930 ;
        RECT 2900.850 674.035 2901.130 674.405 ;
      LAYER via2 ;
        RECT 2900.850 674.080 2901.130 674.360 ;
      LAYER met3 ;
        RECT 2900.825 674.370 2901.155 674.385 ;
        RECT 2917.600 674.370 2924.800 674.820 ;
        RECT 2900.825 674.070 2924.800 674.370 ;
        RECT 2900.825 674.055 2901.155 674.070 ;
        RECT 2917.600 673.620 2924.800 674.070 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 19.850 1759.740 20.170 1759.800 ;
        RECT 685.930 1759.740 686.250 1759.800 ;
        RECT 19.850 1759.600 686.250 1759.740 ;
        RECT 19.850 1759.540 20.170 1759.600 ;
        RECT 685.930 1759.540 686.250 1759.600 ;
      LAYER via ;
        RECT 19.880 1759.540 20.140 1759.800 ;
        RECT 685.960 1759.540 686.220 1759.800 ;
      LAYER met2 ;
        RECT 685.950 1762.715 686.230 1763.085 ;
        RECT 686.020 1759.830 686.160 1762.715 ;
        RECT 19.880 1759.510 20.140 1759.830 ;
        RECT 685.960 1759.510 686.220 1759.830 ;
        RECT 19.940 1544.125 20.080 1759.510 ;
        RECT 19.870 1543.755 20.150 1544.125 ;
      LAYER via2 ;
        RECT 685.950 1762.760 686.230 1763.040 ;
        RECT 19.870 1543.800 20.150 1544.080 ;
      LAYER met3 ;
        RECT 685.925 1763.050 686.255 1763.065 ;
        RECT 715.810 1763.050 719.810 1763.055 ;
        RECT 685.925 1762.750 719.810 1763.050 ;
        RECT 685.925 1762.735 686.255 1762.750 ;
        RECT 715.810 1762.455 719.810 1762.750 ;
        RECT -4.800 1544.090 2.400 1544.540 ;
        RECT 19.845 1544.090 20.175 1544.105 ;
        RECT -4.800 1543.790 20.175 1544.090 ;
        RECT -4.800 1543.340 2.400 1543.790 ;
        RECT 19.845 1543.775 20.175 1543.790 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 1324.880 16.950 1324.940 ;
        RECT 694.210 1324.880 694.530 1324.940 ;
        RECT 16.630 1324.740 694.530 1324.880 ;
        RECT 16.630 1324.680 16.950 1324.740 ;
        RECT 694.210 1324.680 694.530 1324.740 ;
        RECT 694.210 1319.780 694.530 1319.840 ;
        RECT 1278.870 1319.780 1279.190 1319.840 ;
        RECT 694.210 1319.640 1279.190 1319.780 ;
        RECT 694.210 1319.580 694.530 1319.640 ;
        RECT 1278.870 1319.580 1279.190 1319.640 ;
      LAYER via ;
        RECT 16.660 1324.680 16.920 1324.940 ;
        RECT 694.240 1324.680 694.500 1324.940 ;
        RECT 694.240 1319.580 694.500 1319.840 ;
        RECT 1278.900 1319.580 1279.160 1319.840 ;
      LAYER met2 ;
        RECT 16.650 1328.195 16.930 1328.565 ;
        RECT 16.720 1324.970 16.860 1328.195 ;
        RECT 16.660 1324.650 16.920 1324.970 ;
        RECT 694.240 1324.650 694.500 1324.970 ;
        RECT 694.300 1319.870 694.440 1324.650 ;
        RECT 1278.940 1323.135 1279.220 1327.135 ;
        RECT 1278.960 1319.870 1279.100 1323.135 ;
        RECT 694.240 1319.550 694.500 1319.870 ;
        RECT 1278.900 1319.550 1279.160 1319.870 ;
      LAYER via2 ;
        RECT 16.650 1328.240 16.930 1328.520 ;
      LAYER met3 ;
        RECT -4.800 1328.530 2.400 1328.980 ;
        RECT 16.625 1328.530 16.955 1328.545 ;
        RECT -4.800 1328.230 16.955 1328.530 ;
        RECT -4.800 1327.780 2.400 1328.230 ;
        RECT 16.625 1328.215 16.955 1328.230 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 691.910 2383.980 692.230 2384.040 ;
        RECT 830.830 2383.980 831.150 2384.040 ;
        RECT 691.910 2383.840 831.150 2383.980 ;
        RECT 691.910 2383.780 692.230 2383.840 ;
        RECT 830.830 2383.780 831.150 2383.840 ;
        RECT 14.790 1117.820 15.110 1117.880 ;
        RECT 691.910 1117.820 692.230 1117.880 ;
        RECT 14.790 1117.680 692.230 1117.820 ;
        RECT 14.790 1117.620 15.110 1117.680 ;
        RECT 691.910 1117.620 692.230 1117.680 ;
      LAYER via ;
        RECT 691.940 2383.780 692.200 2384.040 ;
        RECT 830.860 2383.780 831.120 2384.040 ;
        RECT 14.820 1117.620 15.080 1117.880 ;
        RECT 691.940 1117.620 692.200 1117.880 ;
      LAYER met2 ;
        RECT 691.940 2383.750 692.200 2384.070 ;
        RECT 830.860 2383.750 831.120 2384.070 ;
        RECT 692.000 1393.845 692.140 2383.750 ;
        RECT 830.920 2377.880 831.060 2383.750 ;
        RECT 830.900 2373.880 831.180 2377.880 ;
        RECT 691.930 1393.475 692.210 1393.845 ;
        RECT 691.930 1390.755 692.210 1391.125 ;
        RECT 692.000 1117.910 692.140 1390.755 ;
        RECT 14.820 1117.590 15.080 1117.910 ;
        RECT 691.940 1117.590 692.200 1117.910 ;
        RECT 14.880 1113.005 15.020 1117.590 ;
        RECT 14.810 1112.635 15.090 1113.005 ;
      LAYER via2 ;
        RECT 691.930 1393.520 692.210 1393.800 ;
        RECT 691.930 1390.800 692.210 1391.080 ;
        RECT 14.810 1112.680 15.090 1112.960 ;
      LAYER met3 ;
        RECT 691.905 1393.810 692.235 1393.825 ;
        RECT 691.905 1393.495 692.450 1393.810 ;
        RECT 692.150 1391.105 692.450 1393.495 ;
        RECT 691.905 1390.790 692.450 1391.105 ;
        RECT 691.905 1390.775 692.235 1390.790 ;
        RECT -4.800 1112.970 2.400 1113.420 ;
        RECT 14.785 1112.970 15.115 1112.985 ;
        RECT -4.800 1112.670 15.115 1112.970 ;
        RECT -4.800 1112.220 2.400 1112.670 ;
        RECT 14.785 1112.655 15.115 1112.670 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 707.625 2378.045 707.795 2380.255 ;
      LAYER mcon ;
        RECT 707.625 2380.085 707.795 2380.255 ;
      LAYER met1 ;
        RECT 25.370 2380.240 25.690 2380.300 ;
        RECT 707.565 2380.240 707.855 2380.285 ;
        RECT 25.370 2380.100 707.855 2380.240 ;
        RECT 25.370 2380.040 25.690 2380.100 ;
        RECT 707.565 2380.055 707.855 2380.100 ;
        RECT 707.565 2378.200 707.855 2378.245 ;
        RECT 742.510 2378.200 742.830 2378.260 ;
        RECT 707.565 2378.060 742.830 2378.200 ;
        RECT 707.565 2378.015 707.855 2378.060 ;
        RECT 742.510 2378.000 742.830 2378.060 ;
        RECT 13.870 897.840 14.190 897.900 ;
        RECT 25.370 897.840 25.690 897.900 ;
        RECT 13.870 897.700 25.690 897.840 ;
        RECT 13.870 897.640 14.190 897.700 ;
        RECT 25.370 897.640 25.690 897.700 ;
      LAYER via ;
        RECT 25.400 2380.040 25.660 2380.300 ;
        RECT 742.540 2378.000 742.800 2378.260 ;
        RECT 13.900 897.640 14.160 897.900 ;
        RECT 25.400 897.640 25.660 897.900 ;
      LAYER met2 ;
        RECT 25.400 2380.010 25.660 2380.330 ;
        RECT 25.460 897.930 25.600 2380.010 ;
        RECT 742.540 2377.970 742.800 2378.290 ;
        RECT 742.600 2377.690 742.740 2377.970 ;
        RECT 744.420 2377.690 744.700 2377.880 ;
        RECT 742.600 2377.550 744.700 2377.690 ;
        RECT 744.420 2373.880 744.700 2377.550 ;
        RECT 13.900 897.610 14.160 897.930 ;
        RECT 25.400 897.610 25.660 897.930 ;
        RECT 13.960 897.445 14.100 897.610 ;
        RECT 13.890 897.075 14.170 897.445 ;
      LAYER via2 ;
        RECT 13.890 897.120 14.170 897.400 ;
      LAYER met3 ;
        RECT -4.800 897.410 2.400 897.860 ;
        RECT 13.865 897.410 14.195 897.425 ;
        RECT -4.800 897.110 14.195 897.410 ;
        RECT -4.800 896.660 2.400 897.110 ;
        RECT 13.865 897.095 14.195 897.110 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.550 682.960 17.870 683.020 ;
        RECT 869.930 682.960 870.250 683.020 ;
        RECT 17.550 682.820 870.250 682.960 ;
        RECT 17.550 682.760 17.870 682.820 ;
        RECT 869.930 682.760 870.250 682.820 ;
      LAYER via ;
        RECT 17.580 682.760 17.840 683.020 ;
        RECT 869.960 682.760 870.220 683.020 ;
      LAYER met2 ;
        RECT 874.140 1323.690 874.420 1327.135 ;
        RECT 870.020 1323.550 874.420 1323.690 ;
        RECT 870.020 683.050 870.160 1323.550 ;
        RECT 874.140 1323.135 874.420 1323.550 ;
        RECT 17.580 682.730 17.840 683.050 ;
        RECT 869.960 682.730 870.220 683.050 ;
        RECT 17.640 681.885 17.780 682.730 ;
        RECT 17.570 681.515 17.850 681.885 ;
      LAYER via2 ;
        RECT 17.570 681.560 17.850 681.840 ;
      LAYER met3 ;
        RECT -4.800 681.850 2.400 682.300 ;
        RECT 17.545 681.850 17.875 681.865 ;
        RECT -4.800 681.550 17.875 681.850 ;
        RECT -4.800 681.100 2.400 681.550 ;
        RECT 17.545 681.535 17.875 681.550 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 31.350 1828.760 31.670 1828.820 ;
        RECT 706.170 1828.760 706.490 1828.820 ;
        RECT 31.350 1828.620 706.490 1828.760 ;
        RECT 31.350 1828.560 31.670 1828.620 ;
        RECT 706.170 1828.560 706.490 1828.620 ;
        RECT 15.250 468.080 15.570 468.140 ;
        RECT 31.350 468.080 31.670 468.140 ;
        RECT 15.250 467.940 31.670 468.080 ;
        RECT 15.250 467.880 15.570 467.940 ;
        RECT 31.350 467.880 31.670 467.940 ;
      LAYER via ;
        RECT 31.380 1828.560 31.640 1828.820 ;
        RECT 706.200 1828.560 706.460 1828.820 ;
        RECT 15.280 467.880 15.540 468.140 ;
        RECT 31.380 467.880 31.640 468.140 ;
      LAYER met2 ;
        RECT 706.190 1830.715 706.470 1831.085 ;
        RECT 706.260 1828.850 706.400 1830.715 ;
        RECT 31.380 1828.530 31.640 1828.850 ;
        RECT 706.200 1828.530 706.460 1828.850 ;
        RECT 31.440 468.170 31.580 1828.530 ;
        RECT 15.280 467.850 15.540 468.170 ;
        RECT 31.380 467.850 31.640 468.170 ;
        RECT 15.340 466.325 15.480 467.850 ;
        RECT 15.270 465.955 15.550 466.325 ;
      LAYER via2 ;
        RECT 706.190 1830.760 706.470 1831.040 ;
        RECT 15.270 466.000 15.550 466.280 ;
      LAYER met3 ;
        RECT 706.165 1831.050 706.495 1831.065 ;
        RECT 715.810 1831.050 719.810 1831.055 ;
        RECT 706.165 1830.750 719.810 1831.050 ;
        RECT 706.165 1830.735 706.495 1830.750 ;
        RECT 715.810 1830.455 719.810 1830.750 ;
        RECT -4.800 466.290 2.400 466.740 ;
        RECT 15.245 466.290 15.575 466.305 ;
        RECT -4.800 465.990 15.575 466.290 ;
        RECT -4.800 465.540 2.400 465.990 ;
        RECT 15.245 465.975 15.575 465.990 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 2378.880 17.410 2378.940 ;
        RECT 784.830 2378.880 785.150 2378.940 ;
        RECT 17.090 2378.740 785.150 2378.880 ;
        RECT 17.090 2378.680 17.410 2378.740 ;
        RECT 784.830 2378.680 785.150 2378.740 ;
      LAYER via ;
        RECT 17.120 2378.680 17.380 2378.940 ;
        RECT 784.860 2378.680 785.120 2378.940 ;
      LAYER met2 ;
        RECT 17.120 2378.650 17.380 2378.970 ;
        RECT 784.860 2378.650 785.120 2378.970 ;
        RECT 17.180 250.765 17.320 2378.650 ;
        RECT 784.920 2377.880 785.060 2378.650 ;
        RECT 784.900 2373.880 785.180 2377.880 ;
        RECT 17.110 250.395 17.390 250.765 ;
      LAYER via2 ;
        RECT 17.110 250.440 17.390 250.720 ;
      LAYER met3 ;
        RECT -4.800 250.730 2.400 251.180 ;
        RECT 17.085 250.730 17.415 250.745 ;
        RECT -4.800 250.430 17.415 250.730 ;
        RECT -4.800 249.980 2.400 250.430 ;
        RECT 17.085 250.415 17.415 250.430 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1759.185 1523.625 1759.355 1554.055 ;
      LAYER mcon ;
        RECT 1759.185 1553.885 1759.355 1554.055 ;
      LAYER met1 ;
        RECT 1757.270 1841.680 1757.590 1841.740 ;
        RECT 1758.190 1841.680 1758.510 1841.740 ;
        RECT 1757.270 1841.540 1758.510 1841.680 ;
        RECT 1757.270 1841.480 1757.590 1841.540 ;
        RECT 1758.190 1841.480 1758.510 1841.540 ;
        RECT 1759.110 1554.040 1759.430 1554.100 ;
        RECT 1758.915 1553.900 1759.430 1554.040 ;
        RECT 1759.110 1553.840 1759.430 1553.900 ;
        RECT 1759.110 1523.780 1759.430 1523.840 ;
        RECT 1758.915 1523.640 1759.430 1523.780 ;
        RECT 1759.110 1523.580 1759.430 1523.640 ;
      LAYER via ;
        RECT 1757.300 1841.480 1757.560 1841.740 ;
        RECT 1758.220 1841.480 1758.480 1841.740 ;
        RECT 1759.140 1553.840 1759.400 1554.100 ;
        RECT 1759.140 1523.580 1759.400 1523.840 ;
      LAYER met2 ;
        RECT 1757.750 1878.995 1758.030 1879.365 ;
        RECT 1757.820 1858.850 1757.960 1878.995 ;
        RECT 1757.820 1858.710 1758.420 1858.850 ;
        RECT 1758.280 1841.770 1758.420 1858.710 ;
        RECT 1757.300 1841.450 1757.560 1841.770 ;
        RECT 1758.220 1841.450 1758.480 1841.770 ;
        RECT 1757.360 1837.205 1757.500 1841.450 ;
        RECT 1757.290 1836.835 1757.570 1837.205 ;
        RECT 1758.210 1773.595 1758.490 1773.965 ;
        RECT 1758.280 1705.285 1758.420 1773.595 ;
        RECT 1758.210 1704.915 1758.490 1705.285 ;
        RECT 1758.210 1673.635 1758.490 1674.005 ;
        RECT 1758.280 1642.725 1758.420 1673.635 ;
        RECT 1758.210 1642.355 1758.490 1642.725 ;
        RECT 1759.130 1553.955 1759.410 1554.325 ;
        RECT 1759.140 1553.810 1759.400 1553.955 ;
        RECT 1759.140 1523.550 1759.400 1523.870 ;
        RECT 1759.200 1521.005 1759.340 1523.550 ;
        RECT 1759.130 1520.635 1759.410 1521.005 ;
        RECT 1755.910 1294.875 1756.190 1295.245 ;
        RECT 1755.980 1242.205 1756.120 1294.875 ;
        RECT 1755.910 1241.835 1756.190 1242.205 ;
        RECT 18.030 886.875 18.310 887.245 ;
        RECT 18.100 35.885 18.240 886.875 ;
        RECT 18.030 35.515 18.310 35.885 ;
      LAYER via2 ;
        RECT 1757.750 1879.040 1758.030 1879.320 ;
        RECT 1757.290 1836.880 1757.570 1837.160 ;
        RECT 1758.210 1773.640 1758.490 1773.920 ;
        RECT 1758.210 1704.960 1758.490 1705.240 ;
        RECT 1758.210 1673.680 1758.490 1673.960 ;
        RECT 1758.210 1642.400 1758.490 1642.680 ;
        RECT 1759.130 1554.000 1759.410 1554.280 ;
        RECT 1759.130 1520.680 1759.410 1520.960 ;
        RECT 1755.910 1294.920 1756.190 1295.200 ;
        RECT 1755.910 1241.880 1756.190 1242.160 ;
        RECT 18.030 886.920 18.310 887.200 ;
        RECT 18.030 35.560 18.310 35.840 ;
      LAYER met3 ;
        RECT 1755.835 1946.055 1759.835 1946.655 ;
        RECT 1757.470 1945.290 1757.850 1945.300 ;
        RECT 1758.430 1945.290 1758.730 1946.055 ;
        RECT 1757.470 1944.990 1758.730 1945.290 ;
        RECT 1757.470 1944.980 1757.850 1944.990 ;
        RECT 1757.725 1879.340 1758.055 1879.345 ;
        RECT 1757.470 1879.330 1758.055 1879.340 ;
        RECT 1757.470 1879.030 1758.280 1879.330 ;
        RECT 1757.470 1879.020 1758.055 1879.030 ;
        RECT 1757.725 1879.015 1758.055 1879.020 ;
        RECT 1756.550 1837.170 1756.930 1837.180 ;
        RECT 1757.265 1837.170 1757.595 1837.185 ;
        RECT 1756.550 1836.870 1757.595 1837.170 ;
        RECT 1756.550 1836.860 1756.930 1836.870 ;
        RECT 1757.265 1836.855 1757.595 1836.870 ;
        RECT 1756.550 1817.450 1756.930 1817.460 ;
        RECT 1758.390 1817.450 1758.770 1817.460 ;
        RECT 1756.550 1817.150 1758.770 1817.450 ;
        RECT 1756.550 1817.140 1756.930 1817.150 ;
        RECT 1758.390 1817.140 1758.770 1817.150 ;
        RECT 1758.185 1773.940 1758.515 1773.945 ;
        RECT 1758.185 1773.930 1758.770 1773.940 ;
        RECT 1757.960 1773.630 1758.770 1773.930 ;
        RECT 1758.185 1773.620 1758.770 1773.630 ;
        RECT 1758.185 1773.615 1758.515 1773.620 ;
        RECT 1757.470 1705.250 1757.850 1705.260 ;
        RECT 1758.185 1705.250 1758.515 1705.265 ;
        RECT 1757.470 1704.950 1758.515 1705.250 ;
        RECT 1757.470 1704.940 1757.850 1704.950 ;
        RECT 1758.185 1704.935 1758.515 1704.950 ;
        RECT 1757.470 1673.970 1757.850 1673.980 ;
        RECT 1758.185 1673.970 1758.515 1673.985 ;
        RECT 1757.470 1673.670 1758.515 1673.970 ;
        RECT 1757.470 1673.660 1757.850 1673.670 ;
        RECT 1758.185 1673.655 1758.515 1673.670 ;
        RECT 1758.185 1642.700 1758.515 1642.705 ;
        RECT 1758.185 1642.690 1758.770 1642.700 ;
        RECT 1757.960 1642.390 1758.770 1642.690 ;
        RECT 1758.185 1642.380 1758.770 1642.390 ;
        RECT 1758.185 1642.375 1758.515 1642.380 ;
        RECT 1756.550 1603.930 1756.930 1603.940 ;
        RECT 1758.390 1603.930 1758.770 1603.940 ;
        RECT 1756.550 1603.630 1758.770 1603.930 ;
        RECT 1756.550 1603.620 1756.930 1603.630 ;
        RECT 1758.390 1603.620 1758.770 1603.630 ;
        RECT 1756.550 1554.290 1756.930 1554.300 ;
        RECT 1759.105 1554.290 1759.435 1554.305 ;
        RECT 1756.550 1553.990 1759.435 1554.290 ;
        RECT 1756.550 1553.980 1756.930 1553.990 ;
        RECT 1759.105 1553.975 1759.435 1553.990 ;
        RECT 1756.550 1520.970 1756.930 1520.980 ;
        RECT 1759.105 1520.970 1759.435 1520.985 ;
        RECT 1756.550 1520.670 1759.435 1520.970 ;
        RECT 1756.550 1520.660 1756.930 1520.670 ;
        RECT 1759.105 1520.655 1759.435 1520.670 ;
        RECT 1756.550 1410.130 1756.930 1410.140 ;
        RECT 1765.750 1410.130 1766.130 1410.140 ;
        RECT 1756.550 1409.830 1766.130 1410.130 ;
        RECT 1756.550 1409.820 1756.930 1409.830 ;
        RECT 1765.750 1409.820 1766.130 1409.830 ;
        RECT 1765.750 1364.570 1766.130 1364.580 ;
        RECT 1756.360 1364.270 1766.130 1364.570 ;
        RECT 1756.360 1363.220 1756.660 1364.270 ;
        RECT 1765.750 1364.260 1766.130 1364.270 ;
        RECT 1756.360 1362.910 1756.930 1363.220 ;
        RECT 1756.550 1362.900 1756.930 1362.910 ;
        RECT 1755.885 1295.220 1756.215 1295.225 ;
        RECT 1755.630 1295.210 1756.215 1295.220 ;
        RECT 1755.430 1294.910 1756.215 1295.210 ;
        RECT 1755.630 1294.900 1756.215 1294.910 ;
        RECT 1755.885 1294.895 1756.215 1294.900 ;
        RECT 1755.885 1242.170 1756.215 1242.185 ;
        RECT 1758.390 1242.170 1758.770 1242.180 ;
        RECT 1755.885 1241.870 1758.770 1242.170 ;
        RECT 1755.885 1241.855 1756.215 1241.870 ;
        RECT 1758.390 1241.860 1758.770 1241.870 ;
        RECT 1756.550 1174.850 1756.930 1174.860 ;
        RECT 1758.390 1174.850 1758.770 1174.860 ;
        RECT 1756.550 1174.550 1758.770 1174.850 ;
        RECT 1756.550 1174.540 1756.930 1174.550 ;
        RECT 1758.390 1174.540 1758.770 1174.550 ;
        RECT 1756.550 1125.890 1756.930 1125.900 ;
        RECT 1755.670 1125.590 1756.930 1125.890 ;
        RECT 1755.670 1124.540 1755.970 1125.590 ;
        RECT 1756.550 1125.580 1756.930 1125.590 ;
        RECT 1755.630 1124.220 1756.010 1124.540 ;
        RECT 1755.630 959.660 1756.010 959.980 ;
        RECT 1755.670 959.290 1755.970 959.660 ;
        RECT 1756.550 959.290 1756.930 959.300 ;
        RECT 1755.670 958.990 1756.930 959.290 ;
        RECT 1756.550 958.980 1756.930 958.990 ;
        RECT 1755.630 912.370 1756.010 912.380 ;
        RECT 1756.550 912.370 1756.930 912.380 ;
        RECT 1755.630 912.070 1756.930 912.370 ;
        RECT 1755.630 912.060 1756.010 912.070 ;
        RECT 1756.550 912.060 1756.930 912.070 ;
        RECT 18.005 887.210 18.335 887.225 ;
        RECT 1755.630 887.210 1756.010 887.220 ;
        RECT 18.005 886.910 1756.010 887.210 ;
        RECT 18.005 886.895 18.335 886.910 ;
        RECT 1755.630 886.900 1756.010 886.910 ;
        RECT -4.800 35.850 2.400 36.300 ;
        RECT 18.005 35.850 18.335 35.865 ;
        RECT -4.800 35.550 18.335 35.850 ;
        RECT -4.800 35.100 2.400 35.550 ;
        RECT 18.005 35.535 18.335 35.550 ;
      LAYER via3 ;
        RECT 1757.500 1944.980 1757.820 1945.300 ;
        RECT 1757.500 1879.020 1757.820 1879.340 ;
        RECT 1756.580 1836.860 1756.900 1837.180 ;
        RECT 1756.580 1817.140 1756.900 1817.460 ;
        RECT 1758.420 1817.140 1758.740 1817.460 ;
        RECT 1758.420 1773.620 1758.740 1773.940 ;
        RECT 1757.500 1704.940 1757.820 1705.260 ;
        RECT 1757.500 1673.660 1757.820 1673.980 ;
        RECT 1758.420 1642.380 1758.740 1642.700 ;
        RECT 1756.580 1603.620 1756.900 1603.940 ;
        RECT 1758.420 1603.620 1758.740 1603.940 ;
        RECT 1756.580 1553.980 1756.900 1554.300 ;
        RECT 1756.580 1520.660 1756.900 1520.980 ;
        RECT 1756.580 1409.820 1756.900 1410.140 ;
        RECT 1765.780 1409.820 1766.100 1410.140 ;
        RECT 1765.780 1364.260 1766.100 1364.580 ;
        RECT 1756.580 1362.900 1756.900 1363.220 ;
        RECT 1755.660 1294.900 1755.980 1295.220 ;
        RECT 1758.420 1241.860 1758.740 1242.180 ;
        RECT 1756.580 1174.540 1756.900 1174.860 ;
        RECT 1758.420 1174.540 1758.740 1174.860 ;
        RECT 1756.580 1125.580 1756.900 1125.900 ;
        RECT 1755.660 1124.220 1755.980 1124.540 ;
        RECT 1755.660 959.660 1755.980 959.980 ;
        RECT 1756.580 958.980 1756.900 959.300 ;
        RECT 1755.660 912.060 1755.980 912.380 ;
        RECT 1756.580 912.060 1756.900 912.380 ;
        RECT 1755.660 886.900 1755.980 887.220 ;
      LAYER met4 ;
        RECT 1757.495 1944.975 1757.825 1945.305 ;
        RECT 1757.510 1879.345 1757.810 1944.975 ;
        RECT 1757.495 1879.015 1757.825 1879.345 ;
        RECT 1756.575 1836.855 1756.905 1837.185 ;
        RECT 1756.590 1817.465 1756.890 1836.855 ;
        RECT 1756.575 1817.135 1756.905 1817.465 ;
        RECT 1758.415 1817.135 1758.745 1817.465 ;
        RECT 1758.430 1773.945 1758.730 1817.135 ;
        RECT 1758.415 1773.615 1758.745 1773.945 ;
        RECT 1757.495 1704.935 1757.825 1705.265 ;
        RECT 1757.510 1673.985 1757.810 1704.935 ;
        RECT 1757.495 1673.655 1757.825 1673.985 ;
        RECT 1758.415 1642.375 1758.745 1642.705 ;
        RECT 1758.430 1603.945 1758.730 1642.375 ;
        RECT 1756.575 1603.615 1756.905 1603.945 ;
        RECT 1758.415 1603.615 1758.745 1603.945 ;
        RECT 1756.590 1603.250 1756.890 1603.615 ;
        RECT 1755.670 1602.950 1756.890 1603.250 ;
        RECT 1755.670 1556.330 1755.970 1602.950 ;
        RECT 1755.670 1556.030 1756.890 1556.330 ;
        RECT 1756.590 1554.305 1756.890 1556.030 ;
        RECT 1756.575 1553.975 1756.905 1554.305 ;
        RECT 1756.575 1520.970 1756.905 1520.985 ;
        RECT 1755.670 1520.670 1756.905 1520.970 ;
        RECT 1755.670 1412.850 1755.970 1520.670 ;
        RECT 1756.575 1520.655 1756.905 1520.670 ;
        RECT 1755.670 1412.550 1756.660 1412.850 ;
        RECT 1756.360 1410.145 1756.660 1412.550 ;
        RECT 1756.360 1409.830 1756.905 1410.145 ;
        RECT 1756.575 1409.815 1756.905 1409.830 ;
        RECT 1765.775 1409.815 1766.105 1410.145 ;
        RECT 1765.790 1364.585 1766.090 1409.815 ;
        RECT 1765.775 1364.255 1766.105 1364.585 ;
        RECT 1756.575 1362.895 1756.905 1363.225 ;
        RECT 1756.590 1361.850 1756.890 1362.895 ;
        RECT 1755.670 1361.550 1756.890 1361.850 ;
        RECT 1755.670 1295.225 1755.970 1361.550 ;
        RECT 1755.655 1294.895 1755.985 1295.225 ;
        RECT 1758.415 1241.855 1758.745 1242.185 ;
        RECT 1758.430 1174.865 1758.730 1241.855 ;
        RECT 1756.575 1174.535 1756.905 1174.865 ;
        RECT 1758.415 1174.535 1758.745 1174.865 ;
        RECT 1756.590 1125.905 1756.890 1174.535 ;
        RECT 1756.575 1125.575 1756.905 1125.905 ;
        RECT 1755.655 1124.215 1755.985 1124.545 ;
        RECT 1755.670 959.985 1755.970 1124.215 ;
        RECT 1755.655 959.655 1755.985 959.985 ;
        RECT 1756.575 958.975 1756.905 959.305 ;
        RECT 1756.590 912.385 1756.890 958.975 ;
        RECT 1755.655 912.055 1755.985 912.385 ;
        RECT 1756.575 912.055 1756.905 912.385 ;
        RECT 1755.670 887.225 1755.970 912.055 ;
        RECT 1755.655 886.895 1755.985 887.225 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 690.605 1368.925 690.775 1393.575 ;
      LAYER mcon ;
        RECT 690.605 1393.405 690.775 1393.575 ;
      LAYER met1 ;
        RECT 690.530 1545.880 690.850 1545.940 ;
        RECT 710.310 1545.880 710.630 1545.940 ;
        RECT 690.530 1545.740 710.630 1545.880 ;
        RECT 690.530 1545.680 690.850 1545.740 ;
        RECT 710.310 1545.680 710.630 1545.740 ;
        RECT 690.530 1393.560 690.850 1393.620 ;
        RECT 690.530 1393.420 691.045 1393.560 ;
        RECT 690.530 1393.360 690.850 1393.420 ;
        RECT 690.530 1369.080 690.850 1369.140 ;
        RECT 690.335 1368.940 690.850 1369.080 ;
        RECT 690.530 1368.880 690.850 1368.940 ;
        RECT 690.530 910.760 690.850 910.820 ;
        RECT 2900.830 910.760 2901.150 910.820 ;
        RECT 690.530 910.620 2901.150 910.760 ;
        RECT 690.530 910.560 690.850 910.620 ;
        RECT 2900.830 910.560 2901.150 910.620 ;
      LAYER via ;
        RECT 690.560 1545.680 690.820 1545.940 ;
        RECT 710.340 1545.680 710.600 1545.940 ;
        RECT 690.560 1393.360 690.820 1393.620 ;
        RECT 690.560 1368.880 690.820 1369.140 ;
        RECT 690.560 910.560 690.820 910.820 ;
        RECT 2900.860 910.560 2901.120 910.820 ;
      LAYER met2 ;
        RECT 710.330 1549.195 710.610 1549.565 ;
        RECT 710.400 1545.970 710.540 1549.195 ;
        RECT 690.560 1545.650 690.820 1545.970 ;
        RECT 710.340 1545.650 710.600 1545.970 ;
        RECT 690.620 1393.650 690.760 1545.650 ;
        RECT 690.560 1393.330 690.820 1393.650 ;
        RECT 690.560 1368.850 690.820 1369.170 ;
        RECT 690.620 910.850 690.760 1368.850 ;
        RECT 690.560 910.530 690.820 910.850 ;
        RECT 2900.860 910.530 2901.120 910.850 ;
        RECT 2900.920 909.685 2901.060 910.530 ;
        RECT 2900.850 909.315 2901.130 909.685 ;
      LAYER via2 ;
        RECT 710.330 1549.240 710.610 1549.520 ;
        RECT 2900.850 909.360 2901.130 909.640 ;
      LAYER met3 ;
        RECT 710.305 1549.530 710.635 1549.545 ;
        RECT 715.810 1549.530 719.810 1549.535 ;
        RECT 710.305 1549.230 719.810 1549.530 ;
        RECT 710.305 1549.215 710.635 1549.230 ;
        RECT 715.810 1548.935 719.810 1549.230 ;
        RECT 2900.825 909.650 2901.155 909.665 ;
        RECT 2917.600 909.650 2924.800 910.100 ;
        RECT 2900.825 909.350 2924.800 909.650 ;
        RECT 2900.825 909.335 2901.155 909.350 ;
        RECT 2917.600 908.900 2924.800 909.350 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1687.350 2382.280 1687.670 2382.340 ;
        RECT 1784.410 2382.280 1784.730 2382.340 ;
        RECT 1687.350 2382.140 1784.730 2382.280 ;
        RECT 1687.350 2382.080 1687.670 2382.140 ;
        RECT 1784.410 2382.080 1784.730 2382.140 ;
        RECT 1784.410 1145.360 1784.730 1145.420 ;
        RECT 2900.830 1145.360 2901.150 1145.420 ;
        RECT 1784.410 1145.220 2901.150 1145.360 ;
        RECT 1784.410 1145.160 1784.730 1145.220 ;
        RECT 2900.830 1145.160 2901.150 1145.220 ;
      LAYER via ;
        RECT 1687.380 2382.080 1687.640 2382.340 ;
        RECT 1784.440 2382.080 1784.700 2382.340 ;
        RECT 1784.440 1145.160 1784.700 1145.420 ;
        RECT 2900.860 1145.160 2901.120 1145.420 ;
      LAYER met2 ;
        RECT 1687.380 2382.050 1687.640 2382.370 ;
        RECT 1784.440 2382.050 1784.700 2382.370 ;
        RECT 1687.440 2377.880 1687.580 2382.050 ;
        RECT 1687.420 2373.880 1687.700 2377.880 ;
        RECT 1784.500 1145.450 1784.640 2382.050 ;
        RECT 1784.440 1145.130 1784.700 1145.450 ;
        RECT 2900.860 1145.130 2901.120 1145.450 ;
        RECT 2900.920 1144.285 2901.060 1145.130 ;
        RECT 2900.850 1143.915 2901.130 1144.285 ;
      LAYER via2 ;
        RECT 2900.850 1143.960 2901.130 1144.240 ;
      LAYER met3 ;
        RECT 2900.825 1144.250 2901.155 1144.265 ;
        RECT 2917.600 1144.250 2924.800 1144.700 ;
        RECT 2900.825 1143.950 2924.800 1144.250 ;
        RECT 2900.825 1143.935 2901.155 1143.950 ;
        RECT 2917.600 1143.500 2924.800 1143.950 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1050.710 2385.000 1051.030 2385.060 ;
        RECT 1785.330 2385.000 1785.650 2385.060 ;
        RECT 1050.710 2384.860 1785.650 2385.000 ;
        RECT 1050.710 2384.800 1051.030 2384.860 ;
        RECT 1785.330 2384.800 1785.650 2384.860 ;
        RECT 1785.330 1379.960 1785.650 1380.020 ;
        RECT 2898.990 1379.960 2899.310 1380.020 ;
        RECT 1785.330 1379.820 2899.310 1379.960 ;
        RECT 1785.330 1379.760 1785.650 1379.820 ;
        RECT 2898.990 1379.760 2899.310 1379.820 ;
      LAYER via ;
        RECT 1050.740 2384.800 1051.000 2385.060 ;
        RECT 1785.360 2384.800 1785.620 2385.060 ;
        RECT 1785.360 1379.760 1785.620 1380.020 ;
        RECT 2899.020 1379.760 2899.280 1380.020 ;
      LAYER met2 ;
        RECT 1050.740 2384.770 1051.000 2385.090 ;
        RECT 1785.360 2384.770 1785.620 2385.090 ;
        RECT 1050.800 2377.880 1050.940 2384.770 ;
        RECT 1050.780 2373.880 1051.060 2377.880 ;
        RECT 1785.420 1380.050 1785.560 2384.770 ;
        RECT 1785.360 1379.730 1785.620 1380.050 ;
        RECT 2899.020 1379.730 2899.280 1380.050 ;
        RECT 2899.080 1378.885 2899.220 1379.730 ;
        RECT 2899.010 1378.515 2899.290 1378.885 ;
      LAYER via2 ;
        RECT 2899.010 1378.560 2899.290 1378.840 ;
      LAYER met3 ;
        RECT 2898.985 1378.850 2899.315 1378.865 ;
        RECT 2917.600 1378.850 2924.800 1379.300 ;
        RECT 2898.985 1378.550 2924.800 1378.850 ;
        RECT 2898.985 1378.535 2899.315 1378.550 ;
        RECT 2917.600 1378.100 2924.800 1378.550 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1733.350 2380.580 1733.670 2380.640 ;
        RECT 1786.250 2380.580 1786.570 2380.640 ;
        RECT 1733.350 2380.440 1786.570 2380.580 ;
        RECT 1733.350 2380.380 1733.670 2380.440 ;
        RECT 1786.250 2380.380 1786.570 2380.440 ;
        RECT 1786.250 1614.560 1786.570 1614.620 ;
        RECT 2898.990 1614.560 2899.310 1614.620 ;
        RECT 1786.250 1614.420 2899.310 1614.560 ;
        RECT 1786.250 1614.360 1786.570 1614.420 ;
        RECT 2898.990 1614.360 2899.310 1614.420 ;
      LAYER via ;
        RECT 1733.380 2380.380 1733.640 2380.640 ;
        RECT 1786.280 2380.380 1786.540 2380.640 ;
        RECT 1786.280 1614.360 1786.540 1614.620 ;
        RECT 2899.020 1614.360 2899.280 1614.620 ;
      LAYER met2 ;
        RECT 1733.380 2380.350 1733.640 2380.670 ;
        RECT 1786.280 2380.350 1786.540 2380.670 ;
        RECT 1733.440 2377.880 1733.580 2380.350 ;
        RECT 1733.420 2373.880 1733.700 2377.880 ;
        RECT 1786.340 1614.650 1786.480 2380.350 ;
        RECT 1786.280 1614.330 1786.540 1614.650 ;
        RECT 2899.020 1614.330 2899.280 1614.650 ;
        RECT 2899.080 1613.485 2899.220 1614.330 ;
        RECT 2899.010 1613.115 2899.290 1613.485 ;
      LAYER via2 ;
        RECT 2899.010 1613.160 2899.290 1613.440 ;
      LAYER met3 ;
        RECT 2898.985 1613.450 2899.315 1613.465 ;
        RECT 2917.600 1613.450 2924.800 1613.900 ;
        RECT 2898.985 1613.150 2924.800 1613.450 ;
        RECT 2898.985 1613.135 2899.315 1613.150 ;
        RECT 2917.600 1612.700 2924.800 1613.150 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1209.870 1319.100 1210.190 1319.160 ;
        RECT 2903.590 1319.100 2903.910 1319.160 ;
        RECT 1209.870 1318.960 2903.910 1319.100 ;
        RECT 1209.870 1318.900 1210.190 1318.960 ;
        RECT 2903.590 1318.900 2903.910 1318.960 ;
      LAYER via ;
        RECT 1209.900 1318.900 1210.160 1319.160 ;
        RECT 2903.620 1318.900 2903.880 1319.160 ;
      LAYER met2 ;
        RECT 2903.610 1847.715 2903.890 1848.085 ;
        RECT 1209.940 1323.135 1210.220 1327.135 ;
        RECT 1209.960 1319.190 1210.100 1323.135 ;
        RECT 2903.680 1319.190 2903.820 1847.715 ;
        RECT 1209.900 1318.870 1210.160 1319.190 ;
        RECT 2903.620 1318.870 2903.880 1319.190 ;
      LAYER via2 ;
        RECT 2903.610 1847.760 2903.890 1848.040 ;
      LAYER met3 ;
        RECT 2903.585 1848.050 2903.915 1848.065 ;
        RECT 2917.600 1848.050 2924.800 1848.500 ;
        RECT 2903.585 1847.750 2924.800 1848.050 ;
        RECT 2903.585 1847.735 2903.915 1847.750 ;
        RECT 2917.600 1847.300 2924.800 1847.750 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1548.430 2387.040 1548.750 2387.100 ;
        RECT 1764.170 2387.040 1764.490 2387.100 ;
        RECT 1548.430 2386.900 1764.490 2387.040 ;
        RECT 1548.430 2386.840 1548.750 2386.900 ;
        RECT 1764.170 2386.840 1764.490 2386.900 ;
        RECT 1764.170 2083.760 1764.490 2083.820 ;
        RECT 2900.830 2083.760 2901.150 2083.820 ;
        RECT 1764.170 2083.620 2901.150 2083.760 ;
        RECT 1764.170 2083.560 1764.490 2083.620 ;
        RECT 2900.830 2083.560 2901.150 2083.620 ;
      LAYER via ;
        RECT 1548.460 2386.840 1548.720 2387.100 ;
        RECT 1764.200 2386.840 1764.460 2387.100 ;
        RECT 1764.200 2083.560 1764.460 2083.820 ;
        RECT 2900.860 2083.560 2901.120 2083.820 ;
      LAYER met2 ;
        RECT 1548.460 2386.810 1548.720 2387.130 ;
        RECT 1764.200 2386.810 1764.460 2387.130 ;
        RECT 1548.520 2377.880 1548.660 2386.810 ;
        RECT 1548.500 2373.880 1548.780 2377.880 ;
        RECT 1764.260 2083.850 1764.400 2386.810 ;
        RECT 1764.200 2083.530 1764.460 2083.850 ;
        RECT 2900.860 2083.530 2901.120 2083.850 ;
        RECT 2900.920 2082.685 2901.060 2083.530 ;
        RECT 2900.850 2082.315 2901.130 2082.685 ;
      LAYER via2 ;
        RECT 2900.850 2082.360 2901.130 2082.640 ;
      LAYER met3 ;
        RECT 2900.825 2082.650 2901.155 2082.665 ;
        RECT 2917.600 2082.650 2924.800 2083.100 ;
        RECT 2900.825 2082.350 2924.800 2082.650 ;
        RECT 2900.825 2082.335 2901.155 2082.350 ;
        RECT 2917.600 2081.900 2924.800 2082.350 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 920.990 1318.080 921.310 1318.140 ;
        RECT 2902.670 1318.080 2902.990 1318.140 ;
        RECT 920.990 1317.940 2902.990 1318.080 ;
        RECT 920.990 1317.880 921.310 1317.940 ;
        RECT 2902.670 1317.880 2902.990 1317.940 ;
      LAYER via ;
        RECT 921.020 1317.880 921.280 1318.140 ;
        RECT 2902.700 1317.880 2902.960 1318.140 ;
      LAYER met2 ;
        RECT 2902.690 2316.915 2902.970 2317.285 ;
        RECT 921.060 1323.135 921.340 1327.135 ;
        RECT 921.080 1318.170 921.220 1323.135 ;
        RECT 2902.760 1318.170 2902.900 2316.915 ;
        RECT 921.020 1317.850 921.280 1318.170 ;
        RECT 2902.700 1317.850 2902.960 1318.170 ;
      LAYER via2 ;
        RECT 2902.690 2316.960 2902.970 2317.240 ;
      LAYER met3 ;
        RECT 2902.665 2317.250 2902.995 2317.265 ;
        RECT 2917.600 2317.250 2924.800 2317.700 ;
        RECT 2902.665 2316.950 2924.800 2317.250 ;
        RECT 2902.665 2316.935 2902.995 2316.950 ;
        RECT 2917.600 2316.500 2924.800 2316.950 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2089.390 146.100 2089.710 146.160 ;
        RECT 2124.810 146.100 2125.130 146.160 ;
        RECT 2089.390 145.960 2125.130 146.100 ;
        RECT 2089.390 145.900 2089.710 145.960 ;
        RECT 2124.810 145.900 2125.130 145.960 ;
        RECT 2208.070 146.100 2208.390 146.160 ;
        RECT 2255.910 146.100 2256.230 146.160 ;
        RECT 2208.070 145.960 2256.230 146.100 ;
        RECT 2208.070 145.900 2208.390 145.960 ;
        RECT 2255.910 145.900 2256.230 145.960 ;
      LAYER via ;
        RECT 2089.420 145.900 2089.680 146.160 ;
        RECT 2124.840 145.900 2125.100 146.160 ;
        RECT 2208.100 145.900 2208.360 146.160 ;
        RECT 2255.940 145.900 2256.200 146.160 ;
      LAYER met2 ;
        RECT 992.770 2382.195 993.050 2382.565 ;
        RECT 992.840 2377.880 992.980 2382.195 ;
        RECT 992.820 2373.880 993.100 2377.880 ;
        RECT 2285.370 147.715 2285.650 148.085 ;
        RECT 2285.440 146.725 2285.580 147.715 ;
        RECT 1945.890 146.610 1946.170 146.725 ;
        RECT 1945.890 146.470 1946.560 146.610 ;
        RECT 1945.890 146.355 1946.170 146.470 ;
        RECT 1946.420 145.365 1946.560 146.470 ;
        RECT 2124.830 146.355 2125.110 146.725 ;
        RECT 2255.930 146.355 2256.210 146.725 ;
        RECT 2285.370 146.355 2285.650 146.725 ;
        RECT 2632.210 146.355 2632.490 146.725 ;
        RECT 2124.900 146.190 2125.040 146.355 ;
        RECT 2256.000 146.190 2256.140 146.355 ;
        RECT 2089.420 146.045 2089.680 146.190 ;
        RECT 2089.410 145.675 2089.690 146.045 ;
        RECT 2124.840 145.870 2125.100 146.190 ;
        RECT 2208.100 146.045 2208.360 146.190 ;
        RECT 2166.690 145.675 2166.970 146.045 ;
        RECT 2208.090 145.675 2208.370 146.045 ;
        RECT 2255.940 145.870 2256.200 146.190 ;
        RECT 2166.760 145.365 2166.900 145.675 ;
        RECT 2632.280 145.365 2632.420 146.355 ;
        RECT 1946.350 144.995 1946.630 145.365 ;
        RECT 2166.690 144.995 2166.970 145.365 ;
        RECT 2632.210 144.995 2632.490 145.365 ;
      LAYER via2 ;
        RECT 992.770 2382.240 993.050 2382.520 ;
        RECT 2285.370 147.760 2285.650 148.040 ;
        RECT 1945.890 146.400 1946.170 146.680 ;
        RECT 2124.830 146.400 2125.110 146.680 ;
        RECT 2255.930 146.400 2256.210 146.680 ;
        RECT 2285.370 146.400 2285.650 146.680 ;
        RECT 2632.210 146.400 2632.490 146.680 ;
        RECT 2089.410 145.720 2089.690 146.000 ;
        RECT 2166.690 145.720 2166.970 146.000 ;
        RECT 2208.090 145.720 2208.370 146.000 ;
        RECT 1946.350 145.040 1946.630 145.320 ;
        RECT 2166.690 145.040 2166.970 145.320 ;
        RECT 2632.210 145.040 2632.490 145.320 ;
      LAYER met3 ;
        RECT 992.745 2382.530 993.075 2382.545 ;
        RECT 1784.150 2382.530 1784.530 2382.540 ;
        RECT 992.745 2382.230 1784.530 2382.530 ;
        RECT 992.745 2382.215 993.075 2382.230 ;
        RECT 1784.150 2382.220 1784.530 2382.230 ;
        RECT 2285.345 148.050 2285.675 148.065 ;
        RECT 2263.510 147.750 2285.675 148.050 ;
        RECT 1945.865 146.690 1946.195 146.705 ;
        RECT 1800.750 146.390 1946.195 146.690 ;
        RECT 1784.150 145.330 1784.530 145.340 ;
        RECT 1800.750 145.330 1801.050 146.390 ;
        RECT 1945.865 146.375 1946.195 146.390 ;
        RECT 1980.110 146.690 1980.490 146.700 ;
        RECT 2124.805 146.690 2125.135 146.705 ;
        RECT 2255.905 146.690 2256.235 146.705 ;
        RECT 2263.510 146.690 2263.810 147.750 ;
        RECT 2285.345 147.735 2285.675 147.750 ;
        RECT 1980.110 146.390 2043.010 146.690 ;
        RECT 1980.110 146.380 1980.490 146.390 ;
        RECT 2042.710 146.010 2043.010 146.390 ;
        RECT 2124.805 146.390 2139.610 146.690 ;
        RECT 2124.805 146.375 2125.135 146.390 ;
        RECT 2089.385 146.010 2089.715 146.025 ;
        RECT 2042.710 145.710 2089.715 146.010 ;
        RECT 2089.385 145.695 2089.715 145.710 ;
        RECT 1784.150 145.030 1801.050 145.330 ;
        RECT 1946.325 145.330 1946.655 145.345 ;
        RECT 1980.110 145.330 1980.490 145.340 ;
        RECT 1946.325 145.030 1980.490 145.330 ;
        RECT 2139.310 145.330 2139.610 146.390 ;
        RECT 2255.905 146.390 2263.810 146.690 ;
        RECT 2285.345 146.690 2285.675 146.705 ;
        RECT 2632.185 146.690 2632.515 146.705 ;
        RECT 2285.345 146.390 2380.650 146.690 ;
        RECT 2255.905 146.375 2256.235 146.390 ;
        RECT 2285.345 146.375 2285.675 146.390 ;
        RECT 2166.665 146.010 2166.995 146.025 ;
        RECT 2208.065 146.010 2208.395 146.025 ;
        RECT 2166.665 145.710 2208.395 146.010 ;
        RECT 2380.350 146.010 2380.650 146.390 ;
        RECT 2524.790 146.390 2546.250 146.690 ;
        RECT 2524.790 146.010 2525.090 146.390 ;
        RECT 2380.350 145.710 2428.490 146.010 ;
        RECT 2166.665 145.695 2166.995 145.710 ;
        RECT 2208.065 145.695 2208.395 145.710 ;
        RECT 2166.665 145.330 2166.995 145.345 ;
        RECT 2139.310 145.030 2166.995 145.330 ;
        RECT 2428.190 145.330 2428.490 145.710 ;
        RECT 2476.950 145.710 2525.090 146.010 ;
        RECT 2545.950 146.010 2546.250 146.390 ;
        RECT 2594.710 146.390 2632.515 146.690 ;
        RECT 2545.950 145.710 2594.090 146.010 ;
        RECT 2476.950 145.330 2477.250 145.710 ;
        RECT 2428.190 145.030 2477.250 145.330 ;
        RECT 2593.790 145.330 2594.090 145.710 ;
        RECT 2594.710 145.330 2595.010 146.390 ;
        RECT 2632.185 146.375 2632.515 146.390 ;
        RECT 2656.310 146.690 2656.690 146.700 ;
        RECT 2917.600 146.690 2924.800 147.140 ;
        RECT 2656.310 146.390 2739.450 146.690 ;
        RECT 2656.310 146.380 2656.690 146.390 ;
        RECT 2739.150 146.010 2739.450 146.390 ;
        RECT 2787.910 146.390 2836.050 146.690 ;
        RECT 2739.150 145.710 2787.290 146.010 ;
        RECT 2593.790 145.030 2595.010 145.330 ;
        RECT 2632.185 145.330 2632.515 145.345 ;
        RECT 2656.310 145.330 2656.690 145.340 ;
        RECT 2632.185 145.030 2656.690 145.330 ;
        RECT 2786.990 145.330 2787.290 145.710 ;
        RECT 2787.910 145.330 2788.210 146.390 ;
        RECT 2835.750 146.010 2836.050 146.390 ;
        RECT 2916.710 146.390 2924.800 146.690 ;
        RECT 2916.710 146.010 2917.010 146.390 ;
        RECT 2835.750 145.710 2883.890 146.010 ;
        RECT 2786.990 145.030 2788.210 145.330 ;
        RECT 2883.590 145.330 2883.890 145.710 ;
        RECT 2884.510 145.710 2917.010 146.010 ;
        RECT 2917.600 145.940 2924.800 146.390 ;
        RECT 2884.510 145.330 2884.810 145.710 ;
        RECT 2883.590 145.030 2884.810 145.330 ;
        RECT 1784.150 145.020 1784.530 145.030 ;
        RECT 1946.325 145.015 1946.655 145.030 ;
        RECT 1980.110 145.020 1980.490 145.030 ;
        RECT 2166.665 145.015 2166.995 145.030 ;
        RECT 2632.185 145.015 2632.515 145.030 ;
        RECT 2656.310 145.020 2656.690 145.030 ;
      LAYER via3 ;
        RECT 1784.180 2382.220 1784.500 2382.540 ;
        RECT 1784.180 145.020 1784.500 145.340 ;
        RECT 1980.140 146.380 1980.460 146.700 ;
        RECT 1980.140 145.020 1980.460 145.340 ;
        RECT 2656.340 146.380 2656.660 146.700 ;
        RECT 2656.340 145.020 2656.660 145.340 ;
      LAYER met4 ;
        RECT 1784.175 2382.215 1784.505 2382.545 ;
        RECT 1784.190 145.345 1784.490 2382.215 ;
        RECT 1980.135 146.375 1980.465 146.705 ;
        RECT 2656.335 146.375 2656.665 146.705 ;
        RECT 1980.150 145.345 1980.450 146.375 ;
        RECT 2656.350 145.345 2656.650 146.375 ;
        RECT 1784.175 145.015 1784.505 145.345 ;
        RECT 1980.135 145.015 1980.465 145.345 ;
        RECT 2656.335 145.015 2656.665 145.345 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 951.810 2491.080 952.130 2491.140 ;
        RECT 2900.830 2491.080 2901.150 2491.140 ;
        RECT 951.810 2490.940 2901.150 2491.080 ;
        RECT 951.810 2490.880 952.130 2490.940 ;
        RECT 2900.830 2490.880 2901.150 2490.940 ;
        RECT 946.750 2388.060 947.070 2388.120 ;
        RECT 951.810 2388.060 952.130 2388.120 ;
        RECT 946.750 2387.920 952.130 2388.060 ;
        RECT 946.750 2387.860 947.070 2387.920 ;
        RECT 951.810 2387.860 952.130 2387.920 ;
      LAYER via ;
        RECT 951.840 2490.880 952.100 2491.140 ;
        RECT 2900.860 2490.880 2901.120 2491.140 ;
        RECT 946.780 2387.860 947.040 2388.120 ;
        RECT 951.840 2387.860 952.100 2388.120 ;
      LAYER met2 ;
        RECT 2900.850 2493.035 2901.130 2493.405 ;
        RECT 2900.920 2491.170 2901.060 2493.035 ;
        RECT 951.840 2490.850 952.100 2491.170 ;
        RECT 2900.860 2490.850 2901.120 2491.170 ;
        RECT 951.900 2388.150 952.040 2490.850 ;
        RECT 946.780 2387.830 947.040 2388.150 ;
        RECT 951.840 2387.830 952.100 2388.150 ;
        RECT 946.840 2377.880 946.980 2387.830 ;
        RECT 946.820 2373.880 947.100 2377.880 ;
      LAYER via2 ;
        RECT 2900.850 2493.080 2901.130 2493.360 ;
      LAYER met3 ;
        RECT 2900.825 2493.370 2901.155 2493.385 ;
        RECT 2917.600 2493.370 2924.800 2493.820 ;
        RECT 2900.825 2493.070 2924.800 2493.370 ;
        RECT 2900.825 2493.055 2901.155 2493.070 ;
        RECT 2917.600 2492.620 2924.800 2493.070 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 972.510 1318.420 972.830 1318.480 ;
        RECT 2902.210 1318.420 2902.530 1318.480 ;
        RECT 972.510 1318.280 2902.530 1318.420 ;
        RECT 972.510 1318.220 972.830 1318.280 ;
        RECT 2902.210 1318.220 2902.530 1318.280 ;
      LAYER via ;
        RECT 972.540 1318.220 972.800 1318.480 ;
        RECT 2902.240 1318.220 2902.500 1318.480 ;
      LAYER met2 ;
        RECT 2902.230 2727.635 2902.510 2728.005 ;
        RECT 972.580 1323.135 972.860 1327.135 ;
        RECT 972.600 1318.510 972.740 1323.135 ;
        RECT 2902.300 1318.510 2902.440 2727.635 ;
        RECT 972.540 1318.190 972.800 1318.510 ;
        RECT 2902.240 1318.190 2902.500 1318.510 ;
      LAYER via2 ;
        RECT 2902.230 2727.680 2902.510 2727.960 ;
      LAYER met3 ;
        RECT 2902.205 2727.970 2902.535 2727.985 ;
        RECT 2917.600 2727.970 2924.800 2728.420 ;
        RECT 2902.205 2727.670 2924.800 2727.970 ;
        RECT 2902.205 2727.655 2902.535 2727.670 ;
        RECT 2917.600 2727.220 2924.800 2727.670 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1435.270 1320.800 1435.590 1320.860 ;
        RECT 2901.750 1320.800 2902.070 1320.860 ;
        RECT 1435.270 1320.660 2902.070 1320.800 ;
        RECT 1435.270 1320.600 1435.590 1320.660 ;
        RECT 2901.750 1320.600 2902.070 1320.660 ;
      LAYER via ;
        RECT 1435.300 1320.600 1435.560 1320.860 ;
        RECT 2901.780 1320.600 2902.040 1320.860 ;
      LAYER met2 ;
        RECT 2901.770 2962.235 2902.050 2962.605 ;
        RECT 1435.340 1323.135 1435.620 1327.135 ;
        RECT 1435.360 1320.890 1435.500 1323.135 ;
        RECT 2901.840 1320.890 2901.980 2962.235 ;
        RECT 1435.300 1320.570 1435.560 1320.890 ;
        RECT 2901.780 1320.570 2902.040 1320.890 ;
      LAYER via2 ;
        RECT 2901.770 2962.280 2902.050 2962.560 ;
      LAYER met3 ;
        RECT 2901.745 2962.570 2902.075 2962.585 ;
        RECT 2917.600 2962.570 2924.800 2963.020 ;
        RECT 2901.745 2962.270 2924.800 2962.570 ;
        RECT 2901.745 2962.255 2902.075 2962.270 ;
        RECT 2917.600 2961.820 2924.800 2962.270 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1470.230 1321.140 1470.550 1321.200 ;
        RECT 2901.290 1321.140 2901.610 1321.200 ;
        RECT 1470.230 1321.000 2901.610 1321.140 ;
        RECT 1470.230 1320.940 1470.550 1321.000 ;
        RECT 2901.290 1320.940 2901.610 1321.000 ;
      LAYER via ;
        RECT 1470.260 1320.940 1470.520 1321.200 ;
        RECT 2901.320 1320.940 2901.580 1321.200 ;
      LAYER met2 ;
        RECT 2901.310 3196.835 2901.590 3197.205 ;
        RECT 1470.300 1323.135 1470.580 1327.135 ;
        RECT 1470.320 1321.230 1470.460 1323.135 ;
        RECT 2901.380 1321.230 2901.520 3196.835 ;
        RECT 1470.260 1320.910 1470.520 1321.230 ;
        RECT 2901.320 1320.910 2901.580 1321.230 ;
      LAYER via2 ;
        RECT 2901.310 3196.880 2901.590 3197.160 ;
      LAYER met3 ;
        RECT 2901.285 3197.170 2901.615 3197.185 ;
        RECT 2917.600 3197.170 2924.800 3197.620 ;
        RECT 2901.285 3196.870 2924.800 3197.170 ;
        RECT 2901.285 3196.855 2901.615 3196.870 ;
        RECT 2917.600 3196.420 2924.800 3196.870 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1783.490 3429.480 1783.810 3429.540 ;
        RECT 2900.830 3429.480 2901.150 3429.540 ;
        RECT 1783.490 3429.340 2901.150 3429.480 ;
        RECT 1783.490 3429.280 1783.810 3429.340 ;
        RECT 2900.830 3429.280 2901.150 3429.340 ;
        RECT 1768.770 1882.820 1769.090 1882.880 ;
        RECT 1783.490 1882.820 1783.810 1882.880 ;
        RECT 1768.770 1882.680 1783.810 1882.820 ;
        RECT 1768.770 1882.620 1769.090 1882.680 ;
        RECT 1783.490 1882.620 1783.810 1882.680 ;
      LAYER via ;
        RECT 1783.520 3429.280 1783.780 3429.540 ;
        RECT 2900.860 3429.280 2901.120 3429.540 ;
        RECT 1768.800 1882.620 1769.060 1882.880 ;
        RECT 1783.520 1882.620 1783.780 1882.880 ;
      LAYER met2 ;
        RECT 2900.850 3431.435 2901.130 3431.805 ;
        RECT 2900.920 3429.570 2901.060 3431.435 ;
        RECT 1783.520 3429.250 1783.780 3429.570 ;
        RECT 2900.860 3429.250 2901.120 3429.570 ;
        RECT 1783.580 1882.910 1783.720 3429.250 ;
        RECT 1768.800 1882.590 1769.060 1882.910 ;
        RECT 1783.520 1882.590 1783.780 1882.910 ;
        RECT 1768.860 1878.685 1769.000 1882.590 ;
        RECT 1768.790 1878.315 1769.070 1878.685 ;
      LAYER via2 ;
        RECT 2900.850 3431.480 2901.130 3431.760 ;
        RECT 1768.790 1878.360 1769.070 1878.640 ;
      LAYER met3 ;
        RECT 2900.825 3431.770 2901.155 3431.785 ;
        RECT 2917.600 3431.770 2924.800 3432.220 ;
        RECT 2900.825 3431.470 2924.800 3431.770 ;
        RECT 2900.825 3431.455 2901.155 3431.470 ;
        RECT 2917.600 3431.020 2924.800 3431.470 ;
        RECT 1755.835 1878.650 1759.835 1878.655 ;
        RECT 1768.765 1878.650 1769.095 1878.665 ;
        RECT 1755.835 1878.350 1769.095 1878.650 ;
        RECT 1755.835 1878.055 1759.835 1878.350 ;
        RECT 1768.765 1878.335 1769.095 1878.350 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1769.690 3502.580 1770.010 3502.640 ;
        RECT 2717.290 3502.580 2717.610 3502.640 ;
        RECT 1769.690 3502.440 2717.610 3502.580 ;
        RECT 1769.690 3502.380 1770.010 3502.440 ;
        RECT 2717.290 3502.380 2717.610 3502.440 ;
      LAYER via ;
        RECT 1769.720 3502.380 1769.980 3502.640 ;
        RECT 2717.320 3502.380 2717.580 3502.640 ;
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
        RECT 2717.380 3502.670 2717.520 3517.600 ;
        RECT 1769.720 3502.350 1769.980 3502.670 ;
        RECT 2717.320 3502.350 2717.580 3502.670 ;
        RECT 1769.780 2297.565 1769.920 3502.350 ;
        RECT 1769.710 2297.195 1769.990 2297.565 ;
      LAYER via2 ;
        RECT 1769.710 2297.240 1769.990 2297.520 ;
      LAYER met3 ;
        RECT 1755.835 2297.530 1759.835 2297.535 ;
        RECT 1769.685 2297.530 1770.015 2297.545 ;
        RECT 1755.835 2297.230 1770.015 2297.530 ;
        RECT 1755.835 2296.935 1759.835 2297.230 ;
        RECT 1769.685 2297.215 1770.015 2297.230 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 709.850 3501.900 710.170 3501.960 ;
        RECT 2392.530 3501.900 2392.850 3501.960 ;
        RECT 709.850 3501.760 2392.850 3501.900 ;
        RECT 709.850 3501.700 710.170 3501.760 ;
        RECT 2392.530 3501.700 2392.850 3501.760 ;
      LAYER via ;
        RECT 709.880 3501.700 710.140 3501.960 ;
        RECT 2392.560 3501.700 2392.820 3501.960 ;
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
        RECT 2392.620 3501.990 2392.760 3517.600 ;
        RECT 709.880 3501.670 710.140 3501.990 ;
        RECT 2392.560 3501.670 2392.820 3501.990 ;
        RECT 709.940 2259.485 710.080 3501.670 ;
        RECT 709.870 2259.115 710.150 2259.485 ;
      LAYER via2 ;
        RECT 709.870 2259.160 710.150 2259.440 ;
      LAYER met3 ;
        RECT 709.845 2259.450 710.175 2259.465 ;
        RECT 715.810 2259.450 719.810 2259.455 ;
        RECT 709.845 2259.150 719.810 2259.450 ;
        RECT 709.845 2259.135 710.175 2259.150 ;
        RECT 715.810 2258.855 719.810 2259.150 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
        RECT 2068.320 3501.845 2068.460 3517.600 ;
        RECT 2068.250 3501.475 2068.530 3501.845 ;
        RECT 729.700 1323.135 729.980 1327.135 ;
        RECT 729.720 1318.365 729.860 1323.135 ;
        RECT 729.650 1317.995 729.930 1318.365 ;
      LAYER via2 ;
        RECT 2068.250 3501.520 2068.530 3501.800 ;
        RECT 729.650 1318.040 729.930 1318.320 ;
      LAYER met3 ;
        RECT 1785.070 3501.810 1785.450 3501.820 ;
        RECT 2068.225 3501.810 2068.555 3501.825 ;
        RECT 1785.070 3501.510 2068.555 3501.810 ;
        RECT 1785.070 3501.500 1785.450 3501.510 ;
        RECT 2068.225 3501.495 2068.555 3501.510 ;
        RECT 729.625 1318.330 729.955 1318.345 ;
        RECT 1785.070 1318.330 1785.450 1318.340 ;
        RECT 729.625 1318.030 1785.450 1318.330 ;
        RECT 729.625 1318.015 729.955 1318.030 ;
        RECT 1785.070 1318.020 1785.450 1318.030 ;
      LAYER via3 ;
        RECT 1785.100 3501.500 1785.420 3501.820 ;
        RECT 1785.100 1318.020 1785.420 1318.340 ;
      LAYER met4 ;
        RECT 1785.095 3501.495 1785.425 3501.825 ;
        RECT 1785.110 1318.345 1785.410 3501.495 ;
        RECT 1785.095 1318.015 1785.425 1318.345 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
        RECT 1744.020 3504.565 1744.160 3517.600 ;
        RECT 1743.950 3504.195 1744.230 3504.565 ;
        RECT 816.180 1323.135 816.460 1327.135 ;
        RECT 816.200 1319.045 816.340 1323.135 ;
        RECT 816.130 1318.675 816.410 1319.045 ;
      LAYER via2 ;
        RECT 1743.950 3504.240 1744.230 3504.520 ;
        RECT 816.130 1318.720 816.410 1319.000 ;
      LAYER met3 ;
        RECT 1743.925 3504.530 1744.255 3504.545 ;
        RECT 1744.590 3504.530 1744.970 3504.540 ;
        RECT 1743.925 3504.230 1744.970 3504.530 ;
        RECT 1743.925 3504.215 1744.255 3504.230 ;
        RECT 1744.590 3504.220 1744.970 3504.230 ;
        RECT 816.105 1319.010 816.435 1319.025 ;
        RECT 1744.590 1319.010 1744.970 1319.020 ;
        RECT 816.105 1318.710 1744.970 1319.010 ;
        RECT 816.105 1318.695 816.435 1318.710 ;
        RECT 1744.590 1318.700 1744.970 1318.710 ;
      LAYER via3 ;
        RECT 1744.620 3504.220 1744.940 3504.540 ;
        RECT 1744.620 1318.700 1744.940 1319.020 ;
      LAYER met4 ;
        RECT 1744.615 3504.215 1744.945 3504.545 ;
        RECT 1744.630 1319.025 1744.930 3504.215 ;
        RECT 1744.615 1318.695 1744.945 1319.025 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1352.010 3504.280 1352.330 3504.340 ;
        RECT 1419.170 3504.280 1419.490 3504.340 ;
        RECT 1352.010 3504.140 1419.490 3504.280 ;
        RECT 1352.010 3504.080 1352.330 3504.140 ;
        RECT 1419.170 3504.080 1419.490 3504.140 ;
      LAYER via ;
        RECT 1352.040 3504.080 1352.300 3504.340 ;
        RECT 1419.200 3504.080 1419.460 3504.340 ;
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
        RECT 1419.260 3504.370 1419.400 3517.600 ;
        RECT 1352.040 3504.050 1352.300 3504.370 ;
        RECT 1419.200 3504.050 1419.460 3504.370 ;
        RECT 1351.620 2377.690 1351.900 2377.880 ;
        RECT 1352.100 2377.690 1352.240 3504.050 ;
        RECT 1351.620 2377.550 1352.240 2377.690 ;
        RECT 1351.620 2373.880 1351.900 2377.550 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2263.730 381.380 2264.050 381.440 ;
        RECT 2284.430 381.380 2284.750 381.440 ;
        RECT 2263.730 381.240 2284.750 381.380 ;
        RECT 2263.730 381.180 2264.050 381.240 ;
        RECT 2284.430 381.180 2284.750 381.240 ;
        RECT 1027.710 380.700 1028.030 380.760 ;
        RECT 1028.630 380.700 1028.950 380.760 ;
        RECT 1027.710 380.560 1028.950 380.700 ;
        RECT 1027.710 380.500 1028.030 380.560 ;
        RECT 1028.630 380.500 1028.950 380.560 ;
        RECT 1317.510 380.700 1317.830 380.760 ;
        RECT 1352.010 380.700 1352.330 380.760 ;
        RECT 1317.510 380.560 1352.330 380.700 ;
        RECT 1317.510 380.500 1317.830 380.560 ;
        RECT 1352.010 380.500 1352.330 380.560 ;
        RECT 1400.770 380.700 1401.090 380.760 ;
        RECT 1421.930 380.700 1422.250 380.760 ;
        RECT 1400.770 380.560 1422.250 380.700 ;
        RECT 1400.770 380.500 1401.090 380.560 ;
        RECT 1421.930 380.500 1422.250 380.560 ;
        RECT 1993.710 380.700 1994.030 380.760 ;
        RECT 2028.210 380.700 2028.530 380.760 ;
        RECT 1993.710 380.560 2028.530 380.700 ;
        RECT 1993.710 380.500 1994.030 380.560 ;
        RECT 2028.210 380.500 2028.530 380.560 ;
        RECT 2090.310 380.700 2090.630 380.760 ;
        RECT 2124.810 380.700 2125.130 380.760 ;
        RECT 2090.310 380.560 2125.130 380.700 ;
        RECT 2090.310 380.500 2090.630 380.560 ;
        RECT 2124.810 380.500 2125.130 380.560 ;
        RECT 2235.210 380.700 2235.530 380.760 ;
        RECT 2238.890 380.700 2239.210 380.760 ;
        RECT 2235.210 380.560 2239.210 380.700 ;
        RECT 2235.210 380.500 2235.530 380.560 ;
        RECT 2238.890 380.500 2239.210 380.560 ;
        RECT 2380.110 380.700 2380.430 380.760 ;
        RECT 2414.610 380.700 2414.930 380.760 ;
        RECT 2380.110 380.560 2414.930 380.700 ;
        RECT 2380.110 380.500 2380.430 380.560 ;
        RECT 2414.610 380.500 2414.930 380.560 ;
        RECT 1795.910 380.360 1796.230 380.420 ;
        RECT 1835.010 380.360 1835.330 380.420 ;
        RECT 1795.910 380.220 1835.330 380.360 ;
        RECT 1795.910 380.160 1796.230 380.220 ;
        RECT 1835.010 380.160 1835.330 380.220 ;
      LAYER via ;
        RECT 2263.760 381.180 2264.020 381.440 ;
        RECT 2284.460 381.180 2284.720 381.440 ;
        RECT 1027.740 380.500 1028.000 380.760 ;
        RECT 1028.660 380.500 1028.920 380.760 ;
        RECT 1317.540 380.500 1317.800 380.760 ;
        RECT 1352.040 380.500 1352.300 380.760 ;
        RECT 1400.800 380.500 1401.060 380.760 ;
        RECT 1421.960 380.500 1422.220 380.760 ;
        RECT 1993.740 380.500 1994.000 380.760 ;
        RECT 2028.240 380.500 2028.500 380.760 ;
        RECT 2090.340 380.500 2090.600 380.760 ;
        RECT 2124.840 380.500 2125.100 380.760 ;
        RECT 2235.240 380.500 2235.500 380.760 ;
        RECT 2238.920 380.500 2239.180 380.760 ;
        RECT 2380.140 380.500 2380.400 380.760 ;
        RECT 2414.640 380.500 2414.900 380.760 ;
        RECT 1795.940 380.160 1796.200 380.420 ;
        RECT 1835.040 380.160 1835.300 380.420 ;
      LAYER met2 ;
        RECT 1973.030 381.635 1973.310 382.005 ;
        RECT 1352.030 380.955 1352.310 381.325 ;
        RECT 1642.290 380.955 1642.570 381.325 ;
        RECT 1795.930 380.955 1796.210 381.325 ;
        RECT 1897.130 380.955 1897.410 381.325 ;
        RECT 1352.100 380.790 1352.240 380.955 ;
        RECT 1027.740 380.645 1028.000 380.790 ;
        RECT 1028.660 380.645 1028.920 380.790 ;
        RECT 1317.540 380.645 1317.800 380.790 ;
        RECT 1027.730 380.275 1028.010 380.645 ;
        RECT 1028.650 380.275 1028.930 380.645 ;
        RECT 1317.530 380.275 1317.810 380.645 ;
        RECT 1352.040 380.470 1352.300 380.790 ;
        RECT 1400.800 380.645 1401.060 380.790 ;
        RECT 1421.960 380.645 1422.220 380.790 ;
        RECT 1400.790 380.275 1401.070 380.645 ;
        RECT 1421.950 380.275 1422.230 380.645 ;
        RECT 1642.360 379.285 1642.500 380.955 ;
        RECT 1796.000 380.450 1796.140 380.955 ;
        RECT 1897.200 380.530 1897.340 380.955 ;
        RECT 1898.050 380.530 1898.330 380.645 ;
        RECT 1795.940 380.130 1796.200 380.450 ;
        RECT 1835.040 380.130 1835.300 380.450 ;
        RECT 1897.200 380.390 1898.330 380.530 ;
        RECT 1898.050 380.275 1898.330 380.390 ;
        RECT 1835.100 379.965 1835.240 380.130 ;
        RECT 1973.100 379.965 1973.240 381.635 ;
        RECT 2263.760 381.325 2264.020 381.470 ;
        RECT 2284.460 381.325 2284.720 381.470 ;
        RECT 2028.230 380.955 2028.510 381.325 ;
        RECT 2124.830 380.955 2125.110 381.325 ;
        RECT 2263.750 380.955 2264.030 381.325 ;
        RECT 2284.450 380.955 2284.730 381.325 ;
        RECT 2414.630 380.955 2414.910 381.325 ;
        RECT 2632.210 380.955 2632.490 381.325 ;
        RECT 2028.300 380.790 2028.440 380.955 ;
        RECT 2124.900 380.790 2125.040 380.955 ;
        RECT 2414.700 380.790 2414.840 380.955 ;
        RECT 1993.740 380.645 1994.000 380.790 ;
        RECT 1993.730 380.275 1994.010 380.645 ;
        RECT 2028.240 380.470 2028.500 380.790 ;
        RECT 2090.340 380.645 2090.600 380.790 ;
        RECT 2090.330 380.275 2090.610 380.645 ;
        RECT 2124.840 380.470 2125.100 380.790 ;
        RECT 2235.240 380.645 2235.500 380.790 ;
        RECT 2238.920 380.645 2239.180 380.790 ;
        RECT 2380.140 380.645 2380.400 380.790 ;
        RECT 2187.850 380.530 2188.130 380.645 ;
        RECT 2187.000 380.390 2188.130 380.530 ;
        RECT 2187.000 379.965 2187.140 380.390 ;
        RECT 2187.850 380.275 2188.130 380.390 ;
        RECT 2235.230 380.275 2235.510 380.645 ;
        RECT 2238.910 380.275 2239.190 380.645 ;
        RECT 2380.130 380.275 2380.410 380.645 ;
        RECT 2414.640 380.470 2414.900 380.790 ;
        RECT 1835.030 379.595 1835.310 379.965 ;
        RECT 1973.030 379.595 1973.310 379.965 ;
        RECT 2138.630 379.850 2138.910 379.965 ;
        RECT 2139.550 379.850 2139.830 379.965 ;
        RECT 2138.630 379.710 2139.830 379.850 ;
        RECT 2138.630 379.595 2138.910 379.710 ;
        RECT 2139.550 379.595 2139.830 379.710 ;
        RECT 2186.930 379.595 2187.210 379.965 ;
        RECT 1642.290 378.915 1642.570 379.285 ;
        RECT 2632.280 378.605 2632.420 380.955 ;
        RECT 2632.210 378.235 2632.490 378.605 ;
      LAYER via2 ;
        RECT 1973.030 381.680 1973.310 381.960 ;
        RECT 1352.030 381.000 1352.310 381.280 ;
        RECT 1642.290 381.000 1642.570 381.280 ;
        RECT 1795.930 381.000 1796.210 381.280 ;
        RECT 1897.130 381.000 1897.410 381.280 ;
        RECT 1027.730 380.320 1028.010 380.600 ;
        RECT 1028.650 380.320 1028.930 380.600 ;
        RECT 1317.530 380.320 1317.810 380.600 ;
        RECT 1400.790 380.320 1401.070 380.600 ;
        RECT 1421.950 380.320 1422.230 380.600 ;
        RECT 1898.050 380.320 1898.330 380.600 ;
        RECT 2028.230 381.000 2028.510 381.280 ;
        RECT 2124.830 381.000 2125.110 381.280 ;
        RECT 2263.750 381.000 2264.030 381.280 ;
        RECT 2284.450 381.000 2284.730 381.280 ;
        RECT 2414.630 381.000 2414.910 381.280 ;
        RECT 2632.210 381.000 2632.490 381.280 ;
        RECT 1993.730 380.320 1994.010 380.600 ;
        RECT 2090.330 380.320 2090.610 380.600 ;
        RECT 2187.850 380.320 2188.130 380.600 ;
        RECT 2235.230 380.320 2235.510 380.600 ;
        RECT 2238.910 380.320 2239.190 380.600 ;
        RECT 2380.130 380.320 2380.410 380.600 ;
        RECT 1835.030 379.640 1835.310 379.920 ;
        RECT 1973.030 379.640 1973.310 379.920 ;
        RECT 2138.630 379.640 2138.910 379.920 ;
        RECT 2139.550 379.640 2139.830 379.920 ;
        RECT 2186.930 379.640 2187.210 379.920 ;
        RECT 1642.290 378.960 1642.570 379.240 ;
        RECT 2632.210 378.280 2632.490 378.560 ;
      LAYER met3 ;
        RECT 693.030 1515.530 693.410 1515.540 ;
        RECT 715.810 1515.530 719.810 1515.535 ;
        RECT 693.030 1515.230 719.810 1515.530 ;
        RECT 693.030 1515.220 693.410 1515.230 ;
        RECT 715.810 1514.935 719.810 1515.230 ;
        RECT 1731.710 381.970 1732.090 381.980 ;
        RECT 1924.910 381.970 1925.290 381.980 ;
        RECT 1973.005 381.970 1973.335 381.985 ;
        RECT 1731.710 381.670 1732.970 381.970 ;
        RECT 1731.710 381.660 1732.090 381.670 ;
        RECT 693.030 381.290 693.410 381.300 ;
        RECT 1352.005 381.290 1352.335 381.305 ;
        RECT 1544.950 381.290 1545.330 381.300 ;
        RECT 1642.265 381.290 1642.595 381.305 ;
        RECT 693.030 380.990 738.450 381.290 ;
        RECT 693.030 380.980 693.410 380.990 ;
        RECT 738.150 379.930 738.450 380.990 ;
        RECT 834.750 380.990 931.650 381.290 ;
        RECT 834.750 379.930 835.050 380.990 ;
        RECT 738.150 379.630 835.050 379.930 ;
        RECT 931.350 379.930 931.650 380.990 ;
        RECT 1076.710 380.990 1124.850 381.290 ;
        RECT 1027.705 380.610 1028.035 380.625 ;
        RECT 980.110 380.310 1028.035 380.610 ;
        RECT 980.110 379.930 980.410 380.310 ;
        RECT 1027.705 380.295 1028.035 380.310 ;
        RECT 1028.625 380.610 1028.955 380.625 ;
        RECT 1028.625 380.310 1076.090 380.610 ;
        RECT 1028.625 380.295 1028.955 380.310 ;
        RECT 931.350 379.630 980.410 379.930 ;
        RECT 1075.790 379.930 1076.090 380.310 ;
        RECT 1076.710 379.930 1077.010 380.990 ;
        RECT 1075.790 379.630 1077.010 379.930 ;
        RECT 1124.550 379.930 1124.850 380.990 ;
        RECT 1221.150 380.990 1270.210 381.290 ;
        RECT 1221.150 379.930 1221.450 380.990 ;
        RECT 1269.910 380.610 1270.210 380.990 ;
        RECT 1352.005 380.990 1366.810 381.290 ;
        RECT 1352.005 380.975 1352.335 380.990 ;
        RECT 1317.505 380.610 1317.835 380.625 ;
        RECT 1269.910 380.310 1317.835 380.610 ;
        RECT 1366.510 380.610 1366.810 380.990 ;
        RECT 1448.390 380.990 1463.410 381.290 ;
        RECT 1400.765 380.610 1401.095 380.625 ;
        RECT 1366.510 380.310 1401.095 380.610 ;
        RECT 1317.505 380.295 1317.835 380.310 ;
        RECT 1400.765 380.295 1401.095 380.310 ;
        RECT 1421.925 380.610 1422.255 380.625 ;
        RECT 1448.390 380.610 1448.690 380.990 ;
        RECT 1421.925 380.310 1448.690 380.610 ;
        RECT 1463.110 380.610 1463.410 380.990 ;
        RECT 1544.950 380.990 1560.010 381.290 ;
        RECT 1544.950 380.980 1545.330 380.990 ;
        RECT 1559.710 380.610 1560.010 380.990 ;
        RECT 1641.590 380.990 1642.595 381.290 ;
        RECT 1732.670 381.290 1732.970 381.670 ;
        RECT 1924.910 381.670 1973.335 381.970 ;
        RECT 1924.910 381.660 1925.290 381.670 ;
        RECT 1973.005 381.655 1973.335 381.670 ;
        RECT 1795.905 381.290 1796.235 381.305 ;
        RECT 1897.105 381.290 1897.435 381.305 ;
        RECT 1732.670 380.990 1796.235 381.290 ;
        RECT 1641.590 380.610 1641.890 380.990 ;
        RECT 1642.265 380.975 1642.595 380.990 ;
        RECT 1795.905 380.975 1796.235 380.990 ;
        RECT 1849.510 380.990 1897.435 381.290 ;
        RECT 1731.710 380.610 1732.090 380.620 ;
        RECT 1463.110 380.310 1510.330 380.610 ;
        RECT 1559.710 380.310 1641.890 380.610 ;
        RECT 1704.150 380.310 1732.090 380.610 ;
        RECT 1421.925 380.295 1422.255 380.310 ;
        RECT 1124.550 379.630 1221.450 379.930 ;
        RECT 1510.030 379.250 1510.330 380.310 ;
        RECT 1544.950 379.620 1545.330 379.940 ;
        RECT 1704.150 379.930 1704.450 380.310 ;
        RECT 1731.710 380.300 1732.090 380.310 ;
        RECT 1690.350 379.630 1704.450 379.930 ;
        RECT 1835.005 379.930 1835.335 379.945 ;
        RECT 1849.510 379.930 1849.810 380.990 ;
        RECT 1897.105 380.975 1897.435 380.990 ;
        RECT 2028.205 381.290 2028.535 381.305 ;
        RECT 2124.805 381.290 2125.135 381.305 ;
        RECT 2125.470 381.290 2125.850 381.300 ;
        RECT 2263.725 381.290 2264.055 381.305 ;
        RECT 2028.205 380.990 2043.010 381.290 ;
        RECT 2028.205 380.975 2028.535 380.990 ;
        RECT 1898.025 380.610 1898.355 380.625 ;
        RECT 1924.910 380.610 1925.290 380.620 ;
        RECT 1993.705 380.610 1994.035 380.625 ;
        RECT 1898.025 380.310 1925.290 380.610 ;
        RECT 1898.025 380.295 1898.355 380.310 ;
        RECT 1924.910 380.300 1925.290 380.310 ;
        RECT 1980.150 380.310 1994.035 380.610 ;
        RECT 2042.710 380.610 2043.010 380.990 ;
        RECT 2124.805 380.990 2125.850 381.290 ;
        RECT 2124.805 380.975 2125.135 380.990 ;
        RECT 2125.470 380.980 2125.850 380.990 ;
        RECT 2262.590 380.990 2264.055 381.290 ;
        RECT 2090.305 380.610 2090.635 380.625 ;
        RECT 2042.710 380.310 2090.635 380.610 ;
        RECT 1835.005 379.630 1849.810 379.930 ;
        RECT 1973.005 379.930 1973.335 379.945 ;
        RECT 1980.150 379.930 1980.450 380.310 ;
        RECT 1993.705 380.295 1994.035 380.310 ;
        RECT 2090.305 380.295 2090.635 380.310 ;
        RECT 2187.825 380.610 2188.155 380.625 ;
        RECT 2235.205 380.610 2235.535 380.625 ;
        RECT 2187.825 380.310 2235.535 380.610 ;
        RECT 2187.825 380.295 2188.155 380.310 ;
        RECT 2235.205 380.295 2235.535 380.310 ;
        RECT 2238.885 380.610 2239.215 380.625 ;
        RECT 2262.590 380.610 2262.890 380.990 ;
        RECT 2263.725 380.975 2264.055 380.990 ;
        RECT 2284.425 381.290 2284.755 381.305 ;
        RECT 2414.605 381.290 2414.935 381.305 ;
        RECT 2632.185 381.290 2632.515 381.305 ;
        RECT 2284.425 380.990 2332.810 381.290 ;
        RECT 2284.425 380.975 2284.755 380.990 ;
        RECT 2238.885 380.310 2262.890 380.610 ;
        RECT 2332.510 380.610 2332.810 380.990 ;
        RECT 2414.605 380.990 2477.250 381.290 ;
        RECT 2414.605 380.975 2414.935 380.990 ;
        RECT 2380.105 380.610 2380.435 380.625 ;
        RECT 2332.510 380.310 2380.435 380.610 ;
        RECT 2476.950 380.610 2477.250 380.990 ;
        RECT 2545.950 380.990 2594.090 381.290 ;
        RECT 2476.950 380.310 2525.090 380.610 ;
        RECT 2238.885 380.295 2239.215 380.310 ;
        RECT 2380.105 380.295 2380.435 380.310 ;
        RECT 1973.005 379.630 1980.450 379.930 ;
        RECT 2125.470 379.930 2125.850 379.940 ;
        RECT 2138.605 379.930 2138.935 379.945 ;
        RECT 2125.470 379.630 2138.935 379.930 ;
        RECT 1544.990 379.250 1545.290 379.620 ;
        RECT 1510.030 378.950 1545.290 379.250 ;
        RECT 1642.265 379.250 1642.595 379.265 ;
        RECT 1690.350 379.250 1690.650 379.630 ;
        RECT 1835.005 379.615 1835.335 379.630 ;
        RECT 1973.005 379.615 1973.335 379.630 ;
        RECT 2125.470 379.620 2125.850 379.630 ;
        RECT 2138.605 379.615 2138.935 379.630 ;
        RECT 2139.525 379.930 2139.855 379.945 ;
        RECT 2186.905 379.930 2187.235 379.945 ;
        RECT 2139.525 379.630 2187.235 379.930 ;
        RECT 2524.790 379.930 2525.090 380.310 ;
        RECT 2545.950 379.930 2546.250 380.990 ;
        RECT 2524.790 379.630 2546.250 379.930 ;
        RECT 2593.790 379.930 2594.090 380.990 ;
        RECT 2594.710 380.990 2632.515 381.290 ;
        RECT 2594.710 379.930 2595.010 380.990 ;
        RECT 2632.185 380.975 2632.515 380.990 ;
        RECT 2656.310 381.290 2656.690 381.300 ;
        RECT 2917.600 381.290 2924.800 381.740 ;
        RECT 2656.310 380.990 2739.450 381.290 ;
        RECT 2656.310 380.980 2656.690 380.990 ;
        RECT 2739.150 380.610 2739.450 380.990 ;
        RECT 2787.910 380.990 2836.050 381.290 ;
        RECT 2739.150 380.310 2787.290 380.610 ;
        RECT 2593.790 379.630 2595.010 379.930 ;
        RECT 2786.990 379.930 2787.290 380.310 ;
        RECT 2787.910 379.930 2788.210 380.990 ;
        RECT 2835.750 380.610 2836.050 380.990 ;
        RECT 2916.710 380.990 2924.800 381.290 ;
        RECT 2916.710 380.610 2917.010 380.990 ;
        RECT 2835.750 380.310 2883.890 380.610 ;
        RECT 2786.990 379.630 2788.210 379.930 ;
        RECT 2883.590 379.930 2883.890 380.310 ;
        RECT 2884.510 380.310 2917.010 380.610 ;
        RECT 2917.600 380.540 2924.800 380.990 ;
        RECT 2884.510 379.930 2884.810 380.310 ;
        RECT 2883.590 379.630 2884.810 379.930 ;
        RECT 2139.525 379.615 2139.855 379.630 ;
        RECT 2186.905 379.615 2187.235 379.630 ;
        RECT 1642.265 378.950 1690.650 379.250 ;
        RECT 1642.265 378.935 1642.595 378.950 ;
        RECT 2632.185 378.570 2632.515 378.585 ;
        RECT 2656.310 378.570 2656.690 378.580 ;
        RECT 2632.185 378.270 2656.690 378.570 ;
        RECT 2632.185 378.255 2632.515 378.270 ;
        RECT 2656.310 378.260 2656.690 378.270 ;
      LAYER via3 ;
        RECT 693.060 1515.220 693.380 1515.540 ;
        RECT 1731.740 381.660 1732.060 381.980 ;
        RECT 693.060 380.980 693.380 381.300 ;
        RECT 1544.980 380.980 1545.300 381.300 ;
        RECT 1924.940 381.660 1925.260 381.980 ;
        RECT 1544.980 379.620 1545.300 379.940 ;
        RECT 1731.740 380.300 1732.060 380.620 ;
        RECT 1924.940 380.300 1925.260 380.620 ;
        RECT 2125.500 380.980 2125.820 381.300 ;
        RECT 2125.500 379.620 2125.820 379.940 ;
        RECT 2656.340 380.980 2656.660 381.300 ;
        RECT 2656.340 378.260 2656.660 378.580 ;
      LAYER met4 ;
        RECT 693.055 1515.215 693.385 1515.545 ;
        RECT 693.070 381.305 693.370 1515.215 ;
        RECT 1731.735 381.655 1732.065 381.985 ;
        RECT 1924.935 381.655 1925.265 381.985 ;
        RECT 693.055 380.975 693.385 381.305 ;
        RECT 1544.975 380.975 1545.305 381.305 ;
        RECT 1544.990 379.945 1545.290 380.975 ;
        RECT 1731.750 380.625 1732.050 381.655 ;
        RECT 1924.950 380.625 1925.250 381.655 ;
        RECT 2125.495 380.975 2125.825 381.305 ;
        RECT 2656.335 380.975 2656.665 381.305 ;
        RECT 1731.735 380.295 1732.065 380.625 ;
        RECT 1924.935 380.295 1925.265 380.625 ;
        RECT 2125.510 379.945 2125.810 380.975 ;
        RECT 1544.975 379.615 1545.305 379.945 ;
        RECT 2125.495 379.615 2125.825 379.945 ;
        RECT 2656.350 378.585 2656.650 380.975 ;
        RECT 2656.335 378.255 2656.665 378.585 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 717.285 1452.225 717.455 1469.735 ;
      LAYER mcon ;
        RECT 717.285 1469.565 717.455 1469.735 ;
      LAYER met1 ;
        RECT 716.290 2163.320 716.610 2163.380 ;
        RECT 717.210 2163.320 717.530 2163.380 ;
        RECT 716.290 2163.180 717.530 2163.320 ;
        RECT 716.290 2163.120 716.610 2163.180 ;
        RECT 717.210 2163.120 717.530 2163.180 ;
        RECT 717.210 1469.720 717.530 1469.780 ;
        RECT 717.015 1469.580 717.530 1469.720 ;
        RECT 717.210 1469.520 717.530 1469.580 ;
        RECT 716.750 1452.380 717.070 1452.440 ;
        RECT 717.225 1452.380 717.515 1452.425 ;
        RECT 716.750 1452.240 717.515 1452.380 ;
        RECT 716.750 1452.180 717.070 1452.240 ;
        RECT 717.225 1452.195 717.515 1452.240 ;
      LAYER via ;
        RECT 716.320 2163.120 716.580 2163.380 ;
        RECT 717.240 2163.120 717.500 2163.380 ;
        RECT 717.240 1469.520 717.500 1469.780 ;
        RECT 716.780 1452.180 717.040 1452.440 ;
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
        RECT 1094.960 3501.845 1095.100 3517.600 ;
        RECT 1094.890 3501.475 1095.170 3501.845 ;
        RECT 717.230 3470.195 717.510 3470.565 ;
        RECT 717.300 3423.645 717.440 3470.195 ;
        RECT 717.230 3423.275 717.510 3423.645 ;
        RECT 717.230 3373.635 717.510 3374.005 ;
        RECT 717.300 3327.085 717.440 3373.635 ;
        RECT 717.230 3326.715 717.510 3327.085 ;
        RECT 717.230 3277.075 717.510 3277.445 ;
        RECT 717.300 3230.525 717.440 3277.075 ;
        RECT 717.230 3230.155 717.510 3230.525 ;
        RECT 716.770 3180.515 717.050 3180.885 ;
        RECT 716.840 3133.965 716.980 3180.515 ;
        RECT 716.770 3133.595 717.050 3133.965 ;
        RECT 716.770 3083.955 717.050 3084.325 ;
        RECT 716.840 3037.405 716.980 3083.955 ;
        RECT 716.770 3037.035 717.050 3037.405 ;
        RECT 716.770 2987.395 717.050 2987.765 ;
        RECT 716.840 2940.845 716.980 2987.395 ;
        RECT 716.770 2940.475 717.050 2940.845 ;
        RECT 717.230 2890.835 717.510 2891.205 ;
        RECT 717.300 2844.285 717.440 2890.835 ;
        RECT 717.230 2843.915 717.510 2844.285 ;
        RECT 717.230 2794.275 717.510 2794.645 ;
        RECT 717.300 2747.725 717.440 2794.275 ;
        RECT 717.230 2747.355 717.510 2747.725 ;
        RECT 716.770 2697.035 717.050 2697.405 ;
        RECT 716.840 2649.805 716.980 2697.035 ;
        RECT 716.770 2649.435 717.050 2649.805 ;
        RECT 717.230 2600.475 717.510 2600.845 ;
        RECT 717.300 2553.245 717.440 2600.475 ;
        RECT 717.230 2552.875 717.510 2553.245 ;
        RECT 717.230 2503.915 717.510 2504.285 ;
        RECT 717.300 2456.685 717.440 2503.915 ;
        RECT 717.230 2456.315 717.510 2456.685 ;
        RECT 716.770 2407.355 717.050 2407.725 ;
        RECT 716.840 2360.125 716.980 2407.355 ;
        RECT 716.770 2359.755 717.050 2360.125 ;
        RECT 717.230 2359.075 717.510 2359.445 ;
        RECT 717.300 2314.565 717.440 2359.075 ;
        RECT 717.230 2314.195 717.510 2314.565 ;
        RECT 717.230 2214.235 717.510 2214.605 ;
        RECT 717.300 2163.410 717.440 2214.235 ;
        RECT 716.320 2163.090 716.580 2163.410 ;
        RECT 717.240 2163.090 717.500 2163.410 ;
        RECT 716.380 2128.245 716.520 2163.090 ;
        RECT 716.310 2127.875 716.590 2128.245 ;
        RECT 717.230 2100.675 717.510 2101.045 ;
        RECT 717.300 2084.725 717.440 2100.675 ;
        RECT 717.230 2084.355 717.510 2084.725 ;
        RECT 714.010 1945.635 714.290 1946.005 ;
        RECT 714.080 1905.205 714.220 1945.635 ;
        RECT 714.010 1904.835 714.290 1905.205 ;
        RECT 717.230 1552.595 717.510 1552.965 ;
        RECT 717.300 1546.165 717.440 1552.595 ;
        RECT 717.230 1545.795 717.510 1546.165 ;
        RECT 717.230 1475.075 717.510 1475.445 ;
        RECT 717.300 1469.810 717.440 1475.075 ;
        RECT 717.240 1469.490 717.500 1469.810 ;
        RECT 716.780 1452.325 717.040 1452.470 ;
        RECT 716.770 1451.955 717.050 1452.325 ;
        RECT 1294.990 1326.410 1295.270 1326.525 ;
        RECT 1296.420 1326.410 1296.700 1327.135 ;
        RECT 1294.990 1326.270 1296.700 1326.410 ;
        RECT 1294.990 1326.155 1295.270 1326.270 ;
        RECT 1296.420 1323.135 1296.700 1326.270 ;
      LAYER via2 ;
        RECT 1094.890 3501.520 1095.170 3501.800 ;
        RECT 717.230 3470.240 717.510 3470.520 ;
        RECT 717.230 3423.320 717.510 3423.600 ;
        RECT 717.230 3373.680 717.510 3373.960 ;
        RECT 717.230 3326.760 717.510 3327.040 ;
        RECT 717.230 3277.120 717.510 3277.400 ;
        RECT 717.230 3230.200 717.510 3230.480 ;
        RECT 716.770 3180.560 717.050 3180.840 ;
        RECT 716.770 3133.640 717.050 3133.920 ;
        RECT 716.770 3084.000 717.050 3084.280 ;
        RECT 716.770 3037.080 717.050 3037.360 ;
        RECT 716.770 2987.440 717.050 2987.720 ;
        RECT 716.770 2940.520 717.050 2940.800 ;
        RECT 717.230 2890.880 717.510 2891.160 ;
        RECT 717.230 2843.960 717.510 2844.240 ;
        RECT 717.230 2794.320 717.510 2794.600 ;
        RECT 717.230 2747.400 717.510 2747.680 ;
        RECT 716.770 2697.080 717.050 2697.360 ;
        RECT 716.770 2649.480 717.050 2649.760 ;
        RECT 717.230 2600.520 717.510 2600.800 ;
        RECT 717.230 2552.920 717.510 2553.200 ;
        RECT 717.230 2503.960 717.510 2504.240 ;
        RECT 717.230 2456.360 717.510 2456.640 ;
        RECT 716.770 2407.400 717.050 2407.680 ;
        RECT 716.770 2359.800 717.050 2360.080 ;
        RECT 717.230 2359.120 717.510 2359.400 ;
        RECT 717.230 2314.240 717.510 2314.520 ;
        RECT 717.230 2214.280 717.510 2214.560 ;
        RECT 716.310 2127.920 716.590 2128.200 ;
        RECT 717.230 2100.720 717.510 2101.000 ;
        RECT 717.230 2084.400 717.510 2084.680 ;
        RECT 714.010 1945.680 714.290 1945.960 ;
        RECT 714.010 1904.880 714.290 1905.160 ;
        RECT 717.230 1552.640 717.510 1552.920 ;
        RECT 717.230 1545.840 717.510 1546.120 ;
        RECT 717.230 1475.120 717.510 1475.400 ;
        RECT 716.770 1452.000 717.050 1452.280 ;
        RECT 1294.990 1326.200 1295.270 1326.480 ;
      LAYER met3 ;
        RECT 716.950 3501.810 717.330 3501.820 ;
        RECT 1094.865 3501.810 1095.195 3501.825 ;
        RECT 716.950 3501.510 1095.195 3501.810 ;
        RECT 716.950 3501.500 717.330 3501.510 ;
        RECT 1094.865 3501.495 1095.195 3501.510 ;
        RECT 717.205 3470.540 717.535 3470.545 ;
        RECT 716.950 3470.530 717.535 3470.540 ;
        RECT 716.750 3470.230 717.535 3470.530 ;
        RECT 716.950 3470.220 717.535 3470.230 ;
        RECT 717.205 3470.215 717.535 3470.220 ;
        RECT 717.205 3423.610 717.535 3423.625 ;
        RECT 716.990 3423.295 717.535 3423.610 ;
        RECT 716.990 3422.940 717.290 3423.295 ;
        RECT 716.950 3422.620 717.330 3422.940 ;
        RECT 717.205 3373.980 717.535 3373.985 ;
        RECT 716.950 3373.970 717.535 3373.980 ;
        RECT 716.750 3373.670 717.535 3373.970 ;
        RECT 716.950 3373.660 717.535 3373.670 ;
        RECT 717.205 3373.655 717.535 3373.660 ;
        RECT 717.205 3327.050 717.535 3327.065 ;
        RECT 716.990 3326.735 717.535 3327.050 ;
        RECT 716.990 3326.380 717.290 3326.735 ;
        RECT 716.950 3326.060 717.330 3326.380 ;
        RECT 717.205 3277.420 717.535 3277.425 ;
        RECT 716.950 3277.410 717.535 3277.420 ;
        RECT 716.750 3277.110 717.535 3277.410 ;
        RECT 716.950 3277.100 717.535 3277.110 ;
        RECT 717.205 3277.095 717.535 3277.100 ;
        RECT 717.205 3230.490 717.535 3230.505 ;
        RECT 716.990 3230.175 717.535 3230.490 ;
        RECT 716.990 3229.820 717.290 3230.175 ;
        RECT 716.950 3229.500 717.330 3229.820 ;
        RECT 716.745 3180.860 717.075 3180.865 ;
        RECT 716.745 3180.850 717.330 3180.860 ;
        RECT 716.520 3180.550 717.330 3180.850 ;
        RECT 716.745 3180.540 717.330 3180.550 ;
        RECT 716.745 3180.535 717.075 3180.540 ;
        RECT 716.745 3133.930 717.075 3133.945 ;
        RECT 716.745 3133.615 717.290 3133.930 ;
        RECT 716.990 3133.260 717.290 3133.615 ;
        RECT 716.950 3132.940 717.330 3133.260 ;
        RECT 716.745 3084.300 717.075 3084.305 ;
        RECT 716.745 3084.290 717.330 3084.300 ;
        RECT 716.520 3083.990 717.330 3084.290 ;
        RECT 716.745 3083.980 717.330 3083.990 ;
        RECT 716.745 3083.975 717.075 3083.980 ;
        RECT 716.745 3037.370 717.075 3037.385 ;
        RECT 716.745 3037.055 717.290 3037.370 ;
        RECT 716.990 3036.700 717.290 3037.055 ;
        RECT 716.950 3036.380 717.330 3036.700 ;
        RECT 716.745 2987.740 717.075 2987.745 ;
        RECT 716.745 2987.730 717.330 2987.740 ;
        RECT 716.520 2987.430 717.330 2987.730 ;
        RECT 716.745 2987.420 717.330 2987.430 ;
        RECT 716.745 2987.415 717.075 2987.420 ;
        RECT 716.745 2940.810 717.075 2940.825 ;
        RECT 716.745 2940.495 717.290 2940.810 ;
        RECT 716.990 2940.140 717.290 2940.495 ;
        RECT 716.950 2939.820 717.330 2940.140 ;
        RECT 717.205 2891.180 717.535 2891.185 ;
        RECT 716.950 2891.170 717.535 2891.180 ;
        RECT 716.750 2890.870 717.535 2891.170 ;
        RECT 716.950 2890.860 717.535 2890.870 ;
        RECT 717.205 2890.855 717.535 2890.860 ;
        RECT 717.205 2844.250 717.535 2844.265 ;
        RECT 716.990 2843.935 717.535 2844.250 ;
        RECT 716.990 2843.580 717.290 2843.935 ;
        RECT 716.950 2843.260 717.330 2843.580 ;
        RECT 717.205 2794.620 717.535 2794.625 ;
        RECT 716.950 2794.610 717.535 2794.620 ;
        RECT 716.750 2794.310 717.535 2794.610 ;
        RECT 716.950 2794.300 717.535 2794.310 ;
        RECT 717.205 2794.295 717.535 2794.300 ;
        RECT 717.205 2747.690 717.535 2747.705 ;
        RECT 716.990 2747.375 717.535 2747.690 ;
        RECT 716.990 2747.020 717.290 2747.375 ;
        RECT 716.950 2746.700 717.330 2747.020 ;
        RECT 716.745 2697.380 717.075 2697.385 ;
        RECT 716.745 2697.370 717.330 2697.380 ;
        RECT 716.520 2697.070 717.330 2697.370 ;
        RECT 716.745 2697.060 717.330 2697.070 ;
        RECT 716.745 2697.055 717.075 2697.060 ;
        RECT 716.745 2649.780 717.075 2649.785 ;
        RECT 716.745 2649.770 717.330 2649.780 ;
        RECT 716.745 2649.470 717.530 2649.770 ;
        RECT 716.745 2649.460 717.330 2649.470 ;
        RECT 716.745 2649.455 717.075 2649.460 ;
        RECT 717.205 2600.820 717.535 2600.825 ;
        RECT 716.950 2600.810 717.535 2600.820 ;
        RECT 716.750 2600.510 717.535 2600.810 ;
        RECT 716.950 2600.500 717.535 2600.510 ;
        RECT 717.205 2600.495 717.535 2600.500 ;
        RECT 717.205 2553.220 717.535 2553.225 ;
        RECT 716.950 2553.210 717.535 2553.220 ;
        RECT 716.750 2552.910 717.535 2553.210 ;
        RECT 716.950 2552.900 717.535 2552.910 ;
        RECT 717.205 2552.895 717.535 2552.900 ;
        RECT 717.205 2504.260 717.535 2504.265 ;
        RECT 716.950 2504.250 717.535 2504.260 ;
        RECT 716.750 2503.950 717.535 2504.250 ;
        RECT 716.950 2503.940 717.535 2503.950 ;
        RECT 717.205 2503.935 717.535 2503.940 ;
        RECT 717.205 2456.660 717.535 2456.665 ;
        RECT 716.950 2456.650 717.535 2456.660 ;
        RECT 716.750 2456.350 717.535 2456.650 ;
        RECT 716.950 2456.340 717.535 2456.350 ;
        RECT 717.205 2456.335 717.535 2456.340 ;
        RECT 716.745 2407.700 717.075 2407.705 ;
        RECT 716.745 2407.690 717.330 2407.700 ;
        RECT 716.520 2407.390 717.330 2407.690 ;
        RECT 716.745 2407.380 717.330 2407.390 ;
        RECT 716.745 2407.375 717.075 2407.380 ;
        RECT 716.745 2360.100 717.075 2360.105 ;
        RECT 716.745 2360.090 717.330 2360.100 ;
        RECT 716.745 2359.790 717.530 2360.090 ;
        RECT 716.745 2359.780 717.330 2359.790 ;
        RECT 716.745 2359.775 717.075 2359.780 ;
        RECT 717.205 2359.420 717.535 2359.425 ;
        RECT 716.950 2359.410 717.535 2359.420 ;
        RECT 716.750 2359.110 717.535 2359.410 ;
        RECT 716.950 2359.100 717.535 2359.110 ;
        RECT 717.205 2359.095 717.535 2359.100 ;
        RECT 715.110 2314.530 715.490 2314.540 ;
        RECT 717.205 2314.530 717.535 2314.545 ;
        RECT 715.110 2314.230 717.535 2314.530 ;
        RECT 715.110 2314.220 715.490 2314.230 ;
        RECT 717.205 2314.215 717.535 2314.230 ;
        RECT 717.205 2214.580 717.535 2214.585 ;
        RECT 716.950 2214.570 717.535 2214.580 ;
        RECT 716.750 2214.270 717.535 2214.570 ;
        RECT 716.950 2214.260 717.535 2214.270 ;
        RECT 717.205 2214.255 717.535 2214.260 ;
        RECT 716.285 2128.210 716.615 2128.225 ;
        RECT 716.950 2128.210 717.330 2128.220 ;
        RECT 716.285 2127.910 717.330 2128.210 ;
        RECT 716.285 2127.895 716.615 2127.910 ;
        RECT 716.950 2127.900 717.330 2127.910 ;
        RECT 717.205 2101.020 717.535 2101.025 ;
        RECT 716.950 2101.010 717.535 2101.020 ;
        RECT 716.750 2100.710 717.535 2101.010 ;
        RECT 716.950 2100.700 717.535 2100.710 ;
        RECT 717.205 2100.695 717.535 2100.700 ;
        RECT 717.205 2084.700 717.535 2084.705 ;
        RECT 716.950 2084.690 717.535 2084.700 ;
        RECT 716.750 2084.390 717.535 2084.690 ;
        RECT 716.950 2084.380 717.535 2084.390 ;
        RECT 717.205 2084.375 717.535 2084.380 ;
        RECT 713.985 1945.970 714.315 1945.985 ;
        RECT 716.950 1945.970 717.330 1945.980 ;
        RECT 713.985 1945.670 717.330 1945.970 ;
        RECT 713.985 1945.655 714.315 1945.670 ;
        RECT 716.950 1945.660 717.330 1945.670 ;
        RECT 713.985 1905.170 714.315 1905.185 ;
        RECT 716.950 1905.170 717.330 1905.180 ;
        RECT 713.985 1904.870 717.330 1905.170 ;
        RECT 713.985 1904.855 714.315 1904.870 ;
        RECT 716.950 1904.860 717.330 1904.870 ;
        RECT 716.030 1552.930 716.410 1552.940 ;
        RECT 717.205 1552.930 717.535 1552.945 ;
        RECT 716.030 1552.630 717.535 1552.930 ;
        RECT 716.030 1552.620 716.410 1552.630 ;
        RECT 717.205 1552.615 717.535 1552.630 ;
        RECT 717.205 1546.140 717.535 1546.145 ;
        RECT 716.950 1546.130 717.535 1546.140 ;
        RECT 716.950 1545.830 717.760 1546.130 ;
        RECT 716.950 1545.820 717.535 1545.830 ;
        RECT 717.205 1545.815 717.535 1545.820 ;
        RECT 717.205 1475.420 717.535 1475.425 ;
        RECT 716.950 1475.410 717.535 1475.420 ;
        RECT 716.950 1475.110 717.760 1475.410 ;
        RECT 716.950 1475.100 717.535 1475.110 ;
        RECT 717.205 1475.095 717.535 1475.100 ;
        RECT 716.745 1452.300 717.075 1452.305 ;
        RECT 716.745 1452.290 717.330 1452.300 ;
        RECT 716.745 1451.990 717.530 1452.290 ;
        RECT 716.745 1451.980 717.330 1451.990 ;
        RECT 716.745 1451.975 717.075 1451.980 ;
        RECT 716.950 1426.820 717.330 1427.140 ;
        RECT 716.990 1425.780 717.290 1426.820 ;
        RECT 716.950 1425.460 717.330 1425.780 ;
        RECT 715.110 1402.650 715.490 1402.660 ;
        RECT 716.950 1402.650 717.330 1402.660 ;
        RECT 715.110 1402.350 717.330 1402.650 ;
        RECT 715.110 1402.340 715.490 1402.350 ;
        RECT 716.950 1402.340 717.330 1402.350 ;
        RECT 1294.965 1326.500 1295.295 1326.505 ;
        RECT 1294.710 1326.490 1295.295 1326.500 ;
        RECT 1294.510 1326.190 1295.295 1326.490 ;
        RECT 1294.710 1326.180 1295.295 1326.190 ;
        RECT 1294.965 1326.175 1295.295 1326.180 ;
        RECT 917.510 1325.810 917.890 1325.820 ;
        RECT 957.070 1325.810 957.450 1325.820 ;
        RECT 917.510 1325.510 957.450 1325.810 ;
        RECT 917.510 1325.500 917.890 1325.510 ;
        RECT 957.070 1325.500 957.450 1325.510 ;
      LAYER via3 ;
        RECT 716.980 3501.500 717.300 3501.820 ;
        RECT 716.980 3470.220 717.300 3470.540 ;
        RECT 716.980 3422.620 717.300 3422.940 ;
        RECT 716.980 3373.660 717.300 3373.980 ;
        RECT 716.980 3326.060 717.300 3326.380 ;
        RECT 716.980 3277.100 717.300 3277.420 ;
        RECT 716.980 3229.500 717.300 3229.820 ;
        RECT 716.980 3180.540 717.300 3180.860 ;
        RECT 716.980 3132.940 717.300 3133.260 ;
        RECT 716.980 3083.980 717.300 3084.300 ;
        RECT 716.980 3036.380 717.300 3036.700 ;
        RECT 716.980 2987.420 717.300 2987.740 ;
        RECT 716.980 2939.820 717.300 2940.140 ;
        RECT 716.980 2890.860 717.300 2891.180 ;
        RECT 716.980 2843.260 717.300 2843.580 ;
        RECT 716.980 2794.300 717.300 2794.620 ;
        RECT 716.980 2746.700 717.300 2747.020 ;
        RECT 716.980 2697.060 717.300 2697.380 ;
        RECT 716.980 2649.460 717.300 2649.780 ;
        RECT 716.980 2600.500 717.300 2600.820 ;
        RECT 716.980 2552.900 717.300 2553.220 ;
        RECT 716.980 2503.940 717.300 2504.260 ;
        RECT 716.980 2456.340 717.300 2456.660 ;
        RECT 716.980 2407.380 717.300 2407.700 ;
        RECT 716.980 2359.780 717.300 2360.100 ;
        RECT 716.980 2359.100 717.300 2359.420 ;
        RECT 715.140 2314.220 715.460 2314.540 ;
        RECT 716.980 2214.260 717.300 2214.580 ;
        RECT 716.980 2127.900 717.300 2128.220 ;
        RECT 716.980 2100.700 717.300 2101.020 ;
        RECT 716.980 2084.380 717.300 2084.700 ;
        RECT 716.980 1945.660 717.300 1945.980 ;
        RECT 716.980 1904.860 717.300 1905.180 ;
        RECT 716.060 1552.620 716.380 1552.940 ;
        RECT 716.980 1545.820 717.300 1546.140 ;
        RECT 716.980 1475.100 717.300 1475.420 ;
        RECT 716.980 1451.980 717.300 1452.300 ;
        RECT 716.980 1426.820 717.300 1427.140 ;
        RECT 716.980 1425.460 717.300 1425.780 ;
        RECT 715.140 1402.340 715.460 1402.660 ;
        RECT 716.980 1402.340 717.300 1402.660 ;
        RECT 1294.740 1326.180 1295.060 1326.500 ;
        RECT 917.540 1325.500 917.860 1325.820 ;
        RECT 957.100 1325.500 957.420 1325.820 ;
      LAYER met4 ;
        RECT 716.975 3501.495 717.305 3501.825 ;
        RECT 716.990 3470.545 717.290 3501.495 ;
        RECT 716.975 3470.215 717.305 3470.545 ;
        RECT 716.975 3422.615 717.305 3422.945 ;
        RECT 716.990 3373.985 717.290 3422.615 ;
        RECT 716.975 3373.655 717.305 3373.985 ;
        RECT 716.975 3326.055 717.305 3326.385 ;
        RECT 716.990 3277.425 717.290 3326.055 ;
        RECT 716.975 3277.095 717.305 3277.425 ;
        RECT 716.975 3229.495 717.305 3229.825 ;
        RECT 716.990 3180.865 717.290 3229.495 ;
        RECT 716.975 3180.535 717.305 3180.865 ;
        RECT 716.975 3132.935 717.305 3133.265 ;
        RECT 716.990 3084.305 717.290 3132.935 ;
        RECT 716.975 3083.975 717.305 3084.305 ;
        RECT 716.975 3036.375 717.305 3036.705 ;
        RECT 716.990 2987.745 717.290 3036.375 ;
        RECT 716.975 2987.415 717.305 2987.745 ;
        RECT 716.975 2939.815 717.305 2940.145 ;
        RECT 716.990 2891.185 717.290 2939.815 ;
        RECT 716.975 2890.855 717.305 2891.185 ;
        RECT 716.975 2843.255 717.305 2843.585 ;
        RECT 716.990 2794.625 717.290 2843.255 ;
        RECT 716.975 2794.295 717.305 2794.625 ;
        RECT 716.975 2746.695 717.305 2747.025 ;
        RECT 716.990 2697.385 717.290 2746.695 ;
        RECT 716.975 2697.055 717.305 2697.385 ;
        RECT 716.975 2649.455 717.305 2649.785 ;
        RECT 716.990 2600.825 717.290 2649.455 ;
        RECT 716.975 2600.495 717.305 2600.825 ;
        RECT 716.975 2552.895 717.305 2553.225 ;
        RECT 716.990 2504.265 717.290 2552.895 ;
        RECT 716.975 2503.935 717.305 2504.265 ;
        RECT 716.975 2456.335 717.305 2456.665 ;
        RECT 716.990 2407.705 717.290 2456.335 ;
        RECT 716.975 2407.375 717.305 2407.705 ;
        RECT 716.975 2359.775 717.305 2360.105 ;
        RECT 716.990 2359.425 717.290 2359.775 ;
        RECT 716.975 2359.095 717.305 2359.425 ;
        RECT 715.135 2314.215 715.465 2314.545 ;
        RECT 715.150 2286.650 715.450 2314.215 ;
        RECT 715.150 2286.350 717.290 2286.650 ;
        RECT 716.990 2218.650 717.290 2286.350 ;
        RECT 716.070 2218.350 717.290 2218.650 ;
        RECT 716.070 2215.250 716.370 2218.350 ;
        RECT 716.070 2214.950 717.290 2215.250 ;
        RECT 716.990 2214.585 717.290 2214.950 ;
        RECT 716.975 2214.255 717.305 2214.585 ;
        RECT 716.975 2127.895 717.305 2128.225 ;
        RECT 716.990 2101.025 717.290 2127.895 ;
        RECT 716.975 2100.695 717.305 2101.025 ;
        RECT 716.975 2084.375 717.305 2084.705 ;
        RECT 716.990 1945.985 717.290 2084.375 ;
        RECT 716.975 1945.655 717.305 1945.985 ;
        RECT 716.975 1904.855 717.305 1905.185 ;
        RECT 716.990 1623.650 717.290 1904.855 ;
        RECT 716.070 1623.350 717.290 1623.650 ;
        RECT 716.070 1552.945 716.370 1623.350 ;
        RECT 716.055 1552.615 716.385 1552.945 ;
        RECT 716.975 1545.815 717.305 1546.145 ;
        RECT 716.990 1475.425 717.290 1545.815 ;
        RECT 716.975 1475.095 717.305 1475.425 ;
        RECT 716.975 1451.975 717.305 1452.305 ;
        RECT 716.990 1427.145 717.290 1451.975 ;
        RECT 716.975 1426.815 717.305 1427.145 ;
        RECT 716.975 1425.455 717.305 1425.785 ;
        RECT 716.990 1402.665 717.290 1425.455 ;
        RECT 715.135 1402.335 715.465 1402.665 ;
        RECT 716.975 1402.335 717.305 1402.665 ;
        RECT 715.150 1328.290 715.450 1402.335 ;
        RECT 917.110 1330.510 918.290 1331.690 ;
        RECT 956.670 1330.510 957.850 1331.690 ;
        RECT 1294.310 1330.510 1295.490 1331.690 ;
        RECT 714.710 1327.110 715.890 1328.290 ;
        RECT 917.550 1325.825 917.850 1330.510 ;
        RECT 957.110 1325.825 957.410 1330.510 ;
        RECT 1294.750 1326.505 1295.050 1330.510 ;
        RECT 1294.735 1326.175 1295.065 1326.505 ;
        RECT 917.535 1325.495 917.865 1325.825 ;
        RECT 957.095 1325.495 957.425 1325.825 ;
      LAYER met5 ;
        RECT 727.380 1333.700 918.500 1335.300 ;
        RECT 727.380 1328.500 728.980 1333.700 ;
        RECT 916.900 1330.300 918.500 1333.700 ;
        RECT 956.460 1333.700 1295.700 1335.300 ;
        RECT 956.460 1330.300 958.060 1333.700 ;
        RECT 1294.100 1330.300 1295.700 1333.700 ;
        RECT 714.500 1326.900 728.980 1328.500 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 720.505 2373.625 720.675 2377.875 ;
      LAYER mcon ;
        RECT 720.505 2377.705 720.675 2377.875 ;
      LAYER met1 ;
        RECT 765.970 3498.500 766.290 3498.560 ;
        RECT 770.570 3498.500 770.890 3498.560 ;
        RECT 765.970 3498.360 770.890 3498.500 ;
        RECT 765.970 3498.300 766.290 3498.360 ;
        RECT 770.570 3498.300 770.890 3498.360 ;
        RECT 765.970 2378.200 766.290 2378.260 ;
        RECT 743.060 2378.060 766.290 2378.200 ;
        RECT 720.445 2377.860 720.735 2377.905 ;
        RECT 743.060 2377.860 743.200 2378.060 ;
        RECT 765.970 2378.000 766.290 2378.060 ;
        RECT 720.445 2377.720 743.200 2377.860 ;
        RECT 720.445 2377.675 720.735 2377.720 ;
        RECT 691.450 2373.780 691.770 2373.840 ;
        RECT 720.445 2373.780 720.735 2373.825 ;
        RECT 691.450 2373.640 720.735 2373.780 ;
        RECT 691.450 2373.580 691.770 2373.640 ;
        RECT 720.445 2373.595 720.735 2373.640 ;
        RECT 691.450 1317.740 691.770 1317.800 ;
        RECT 833.590 1317.740 833.910 1317.800 ;
        RECT 691.450 1317.600 833.910 1317.740 ;
        RECT 691.450 1317.540 691.770 1317.600 ;
        RECT 833.590 1317.540 833.910 1317.600 ;
      LAYER via ;
        RECT 766.000 3498.300 766.260 3498.560 ;
        RECT 770.600 3498.300 770.860 3498.560 ;
        RECT 766.000 2378.000 766.260 2378.260 ;
        RECT 691.480 2373.580 691.740 2373.840 ;
        RECT 691.480 1317.540 691.740 1317.800 ;
        RECT 833.620 1317.540 833.880 1317.800 ;
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
        RECT 770.660 3498.590 770.800 3517.600 ;
        RECT 766.000 3498.270 766.260 3498.590 ;
        RECT 770.600 3498.270 770.860 3498.590 ;
        RECT 766.060 2378.290 766.200 3498.270 ;
        RECT 766.000 2377.970 766.260 2378.290 ;
        RECT 691.480 2373.550 691.740 2373.870 ;
        RECT 691.540 1317.830 691.680 2373.550 ;
        RECT 833.660 1323.135 833.940 1327.135 ;
        RECT 833.680 1317.830 833.820 1323.135 ;
        RECT 691.480 1317.510 691.740 1317.830 ;
        RECT 833.620 1317.510 833.880 1317.830 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 445.810 3498.500 446.130 3498.560 ;
        RECT 448.110 3498.500 448.430 3498.560 ;
        RECT 445.810 3498.360 448.430 3498.500 ;
        RECT 445.810 3498.300 446.130 3498.360 ;
        RECT 448.110 3498.300 448.430 3498.360 ;
        RECT 448.110 1321.140 448.430 1321.200 ;
        RECT 961.470 1321.140 961.790 1321.200 ;
        RECT 448.110 1321.000 961.790 1321.140 ;
        RECT 448.110 1320.940 448.430 1321.000 ;
        RECT 961.470 1320.940 961.790 1321.000 ;
      LAYER via ;
        RECT 445.840 3498.300 446.100 3498.560 ;
        RECT 448.140 3498.300 448.400 3498.560 ;
        RECT 448.140 1320.940 448.400 1321.200 ;
        RECT 961.500 1320.940 961.760 1321.200 ;
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
        RECT 445.900 3498.590 446.040 3517.600 ;
        RECT 445.840 3498.270 446.100 3498.590 ;
        RECT 448.140 3498.270 448.400 3498.590 ;
        RECT 448.200 1321.230 448.340 3498.270 ;
        RECT 961.540 1323.135 961.820 1327.135 ;
        RECT 961.560 1321.230 961.700 1323.135 ;
        RECT 448.140 1320.910 448.400 1321.230 ;
        RECT 961.500 1320.910 961.760 1321.230 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 121.510 3498.500 121.830 3498.560 ;
        RECT 123.810 3498.500 124.130 3498.560 ;
        RECT 121.510 3498.360 124.130 3498.500 ;
        RECT 121.510 3498.300 121.830 3498.360 ;
        RECT 123.810 3498.300 124.130 3498.360 ;
        RECT 123.810 1321.480 124.130 1321.540 ;
        RECT 1556.710 1321.480 1557.030 1321.540 ;
        RECT 123.810 1321.340 1557.030 1321.480 ;
        RECT 123.810 1321.280 124.130 1321.340 ;
        RECT 1556.710 1321.280 1557.030 1321.340 ;
      LAYER via ;
        RECT 121.540 3498.300 121.800 3498.560 ;
        RECT 123.840 3498.300 124.100 3498.560 ;
        RECT 123.840 1321.280 124.100 1321.540 ;
        RECT 1556.740 1321.280 1557.000 1321.540 ;
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
        RECT 121.600 3498.590 121.740 3517.600 ;
        RECT 121.540 3498.270 121.800 3498.590 ;
        RECT 123.840 3498.270 124.100 3498.590 ;
        RECT 123.900 1321.570 124.040 3498.270 ;
        RECT 1556.780 1323.135 1557.060 1327.135 ;
        RECT 1556.800 1321.570 1556.940 1323.135 ;
        RECT 123.840 1321.250 124.100 1321.570 ;
        RECT 1556.740 1321.250 1557.000 1321.570 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1753.665 3284.485 1753.835 3313.895 ;
        RECT 1753.665 3236.205 1753.835 3260.175 ;
        RECT 1753.205 3139.645 1753.375 3153.755 ;
        RECT 1752.745 3043.085 1752.915 3057.875 ;
        RECT 1753.205 2994.805 1753.375 3034.075 ;
        RECT 1753.205 2898.245 1753.375 2946.355 ;
      LAYER mcon ;
        RECT 1753.665 3313.725 1753.835 3313.895 ;
        RECT 1753.665 3260.005 1753.835 3260.175 ;
        RECT 1753.205 3153.585 1753.375 3153.755 ;
        RECT 1752.745 3057.705 1752.915 3057.875 ;
        RECT 1753.205 3033.905 1753.375 3034.075 ;
        RECT 1753.205 2946.185 1753.375 2946.355 ;
      LAYER met1 ;
        RECT 17.090 3339.720 17.410 3339.780 ;
        RECT 1752.670 3339.720 1752.990 3339.780 ;
        RECT 17.090 3339.580 1752.990 3339.720 ;
        RECT 17.090 3339.520 17.410 3339.580 ;
        RECT 1752.670 3339.520 1752.990 3339.580 ;
        RECT 1752.670 3313.880 1752.990 3313.940 ;
        RECT 1753.605 3313.880 1753.895 3313.925 ;
        RECT 1752.670 3313.740 1753.895 3313.880 ;
        RECT 1752.670 3313.680 1752.990 3313.740 ;
        RECT 1753.605 3313.695 1753.895 3313.740 ;
        RECT 1753.590 3284.640 1753.910 3284.700 ;
        RECT 1753.395 3284.500 1753.910 3284.640 ;
        RECT 1753.590 3284.440 1753.910 3284.500 ;
        RECT 1753.590 3260.160 1753.910 3260.220 ;
        RECT 1753.395 3260.020 1753.910 3260.160 ;
        RECT 1753.590 3259.960 1753.910 3260.020 ;
        RECT 1753.605 3236.360 1753.895 3236.405 ;
        RECT 1754.050 3236.360 1754.370 3236.420 ;
        RECT 1753.605 3236.220 1754.370 3236.360 ;
        RECT 1753.605 3236.175 1753.895 3236.220 ;
        RECT 1754.050 3236.160 1754.370 3236.220 ;
        RECT 1753.130 3201.680 1753.450 3201.740 ;
        RECT 1754.050 3201.680 1754.370 3201.740 ;
        RECT 1753.130 3201.540 1754.370 3201.680 ;
        RECT 1753.130 3201.480 1753.450 3201.540 ;
        RECT 1754.050 3201.480 1754.370 3201.540 ;
        RECT 1753.130 3153.740 1753.450 3153.800 ;
        RECT 1752.935 3153.600 1753.450 3153.740 ;
        RECT 1753.130 3153.540 1753.450 3153.600 ;
        RECT 1752.670 3139.800 1752.990 3139.860 ;
        RECT 1753.145 3139.800 1753.435 3139.845 ;
        RECT 1752.670 3139.660 1753.435 3139.800 ;
        RECT 1752.670 3139.600 1752.990 3139.660 ;
        RECT 1753.145 3139.615 1753.435 3139.660 ;
        RECT 1752.685 3057.860 1752.975 3057.905 ;
        RECT 1753.130 3057.860 1753.450 3057.920 ;
        RECT 1752.685 3057.720 1753.450 3057.860 ;
        RECT 1752.685 3057.675 1752.975 3057.720 ;
        RECT 1753.130 3057.660 1753.450 3057.720 ;
        RECT 1752.670 3043.240 1752.990 3043.300 ;
        RECT 1752.475 3043.100 1752.990 3043.240 ;
        RECT 1752.670 3043.040 1752.990 3043.100 ;
        RECT 1752.670 3034.060 1752.990 3034.120 ;
        RECT 1753.145 3034.060 1753.435 3034.105 ;
        RECT 1752.670 3033.920 1753.435 3034.060 ;
        RECT 1752.670 3033.860 1752.990 3033.920 ;
        RECT 1753.145 3033.875 1753.435 3033.920 ;
        RECT 1753.130 2994.960 1753.450 2995.020 ;
        RECT 1753.130 2994.820 1753.645 2994.960 ;
        RECT 1753.130 2994.760 1753.450 2994.820 ;
        RECT 1753.130 2960.620 1753.450 2960.680 ;
        RECT 1752.760 2960.480 1753.450 2960.620 ;
        RECT 1752.760 2960.000 1752.900 2960.480 ;
        RECT 1753.130 2960.420 1753.450 2960.480 ;
        RECT 1752.670 2959.740 1752.990 2960.000 ;
        RECT 1752.670 2946.340 1752.990 2946.400 ;
        RECT 1753.145 2946.340 1753.435 2946.385 ;
        RECT 1752.670 2946.200 1753.435 2946.340 ;
        RECT 1752.670 2946.140 1752.990 2946.200 ;
        RECT 1753.145 2946.155 1753.435 2946.200 ;
        RECT 1753.130 2898.400 1753.450 2898.460 ;
        RECT 1753.130 2898.260 1753.645 2898.400 ;
        RECT 1753.130 2898.200 1753.450 2898.260 ;
        RECT 1753.130 2864.060 1753.450 2864.120 ;
        RECT 1752.760 2863.920 1753.450 2864.060 ;
        RECT 1752.760 2863.440 1752.900 2863.920 ;
        RECT 1753.130 2863.860 1753.450 2863.920 ;
        RECT 1752.670 2863.180 1752.990 2863.440 ;
        RECT 1753.130 2767.500 1753.450 2767.560 ;
        RECT 1752.760 2767.360 1753.450 2767.500 ;
        RECT 1752.760 2766.880 1752.900 2767.360 ;
        RECT 1753.130 2767.300 1753.450 2767.360 ;
        RECT 1752.670 2766.620 1752.990 2766.880 ;
        RECT 1752.670 2714.460 1752.990 2714.520 ;
        RECT 1754.050 2714.460 1754.370 2714.520 ;
        RECT 1752.670 2714.320 1754.370 2714.460 ;
        RECT 1752.670 2714.260 1752.990 2714.320 ;
        RECT 1754.050 2714.260 1754.370 2714.320 ;
        RECT 1754.050 2623.340 1754.370 2623.400 ;
        RECT 1753.220 2623.200 1754.370 2623.340 ;
        RECT 1753.220 2622.380 1753.360 2623.200 ;
        RECT 1754.050 2623.140 1754.370 2623.200 ;
        RECT 1753.130 2622.120 1753.450 2622.380 ;
        RECT 1753.130 2573.360 1753.450 2573.420 ;
        RECT 1754.510 2573.360 1754.830 2573.420 ;
        RECT 1753.130 2573.220 1754.830 2573.360 ;
        RECT 1753.130 2573.160 1753.450 2573.220 ;
        RECT 1754.510 2573.160 1754.830 2573.220 ;
        RECT 1754.510 2512.500 1754.830 2512.560 ;
        RECT 1753.220 2512.360 1754.830 2512.500 ;
        RECT 1753.220 2512.220 1753.360 2512.360 ;
        RECT 1754.510 2512.300 1754.830 2512.360 ;
        RECT 1753.130 2511.960 1753.450 2512.220 ;
        RECT 1753.130 2476.940 1753.450 2477.200 ;
        RECT 1753.220 2476.800 1753.360 2476.940 ;
        RECT 1755.430 2476.800 1755.750 2476.860 ;
        RECT 1753.220 2476.660 1755.750 2476.800 ;
        RECT 1755.430 2476.600 1755.750 2476.660 ;
        RECT 1754.510 2042.620 1754.830 2042.680 ;
        RECT 1754.510 2042.480 1755.200 2042.620 ;
        RECT 1754.510 2042.420 1754.830 2042.480 ;
        RECT 1755.060 2041.320 1755.200 2042.480 ;
        RECT 1754.970 2041.060 1755.290 2041.320 ;
        RECT 1754.970 1973.260 1755.290 1973.320 ;
        RECT 1757.270 1973.260 1757.590 1973.320 ;
        RECT 1754.970 1973.120 1757.590 1973.260 ;
        RECT 1754.970 1973.060 1755.290 1973.120 ;
        RECT 1757.270 1973.060 1757.590 1973.120 ;
      LAYER via ;
        RECT 17.120 3339.520 17.380 3339.780 ;
        RECT 1752.700 3339.520 1752.960 3339.780 ;
        RECT 1752.700 3313.680 1752.960 3313.940 ;
        RECT 1753.620 3284.440 1753.880 3284.700 ;
        RECT 1753.620 3259.960 1753.880 3260.220 ;
        RECT 1754.080 3236.160 1754.340 3236.420 ;
        RECT 1753.160 3201.480 1753.420 3201.740 ;
        RECT 1754.080 3201.480 1754.340 3201.740 ;
        RECT 1753.160 3153.540 1753.420 3153.800 ;
        RECT 1752.700 3139.600 1752.960 3139.860 ;
        RECT 1753.160 3057.660 1753.420 3057.920 ;
        RECT 1752.700 3043.040 1752.960 3043.300 ;
        RECT 1752.700 3033.860 1752.960 3034.120 ;
        RECT 1753.160 2994.760 1753.420 2995.020 ;
        RECT 1753.160 2960.420 1753.420 2960.680 ;
        RECT 1752.700 2959.740 1752.960 2960.000 ;
        RECT 1752.700 2946.140 1752.960 2946.400 ;
        RECT 1753.160 2898.200 1753.420 2898.460 ;
        RECT 1753.160 2863.860 1753.420 2864.120 ;
        RECT 1752.700 2863.180 1752.960 2863.440 ;
        RECT 1753.160 2767.300 1753.420 2767.560 ;
        RECT 1752.700 2766.620 1752.960 2766.880 ;
        RECT 1752.700 2714.260 1752.960 2714.520 ;
        RECT 1754.080 2714.260 1754.340 2714.520 ;
        RECT 1754.080 2623.140 1754.340 2623.400 ;
        RECT 1753.160 2622.120 1753.420 2622.380 ;
        RECT 1753.160 2573.160 1753.420 2573.420 ;
        RECT 1754.540 2573.160 1754.800 2573.420 ;
        RECT 1754.540 2512.300 1754.800 2512.560 ;
        RECT 1753.160 2511.960 1753.420 2512.220 ;
        RECT 1753.160 2476.940 1753.420 2477.200 ;
        RECT 1755.460 2476.600 1755.720 2476.860 ;
        RECT 1754.540 2042.420 1754.800 2042.680 ;
        RECT 1755.000 2041.060 1755.260 2041.320 ;
        RECT 1755.000 1973.060 1755.260 1973.320 ;
        RECT 1757.300 1973.060 1757.560 1973.320 ;
      LAYER met2 ;
        RECT 17.110 3339.635 17.390 3340.005 ;
        RECT 17.120 3339.490 17.380 3339.635 ;
        RECT 1752.700 3339.490 1752.960 3339.810 ;
        RECT 1752.760 3313.970 1752.900 3339.490 ;
        RECT 1752.700 3313.650 1752.960 3313.970 ;
        RECT 1753.620 3284.410 1753.880 3284.730 ;
        RECT 1753.680 3260.250 1753.820 3284.410 ;
        RECT 1753.620 3259.930 1753.880 3260.250 ;
        RECT 1754.080 3236.130 1754.340 3236.450 ;
        RECT 1754.140 3201.770 1754.280 3236.130 ;
        RECT 1753.160 3201.450 1753.420 3201.770 ;
        RECT 1754.080 3201.450 1754.340 3201.770 ;
        RECT 1753.220 3153.830 1753.360 3201.450 ;
        RECT 1753.160 3153.510 1753.420 3153.830 ;
        RECT 1752.700 3139.570 1752.960 3139.890 ;
        RECT 1752.760 3105.970 1752.900 3139.570 ;
        RECT 1752.760 3105.830 1753.360 3105.970 ;
        RECT 1753.220 3057.950 1753.360 3105.830 ;
        RECT 1753.160 3057.630 1753.420 3057.950 ;
        RECT 1752.700 3043.010 1752.960 3043.330 ;
        RECT 1752.760 3034.150 1752.900 3043.010 ;
        RECT 1752.700 3033.830 1752.960 3034.150 ;
        RECT 1753.160 2994.730 1753.420 2995.050 ;
        RECT 1753.220 2960.710 1753.360 2994.730 ;
        RECT 1753.160 2960.390 1753.420 2960.710 ;
        RECT 1752.700 2959.710 1752.960 2960.030 ;
        RECT 1752.760 2946.430 1752.900 2959.710 ;
        RECT 1752.700 2946.110 1752.960 2946.430 ;
        RECT 1753.160 2898.170 1753.420 2898.490 ;
        RECT 1753.220 2864.150 1753.360 2898.170 ;
        RECT 1753.160 2863.830 1753.420 2864.150 ;
        RECT 1752.700 2863.150 1752.960 2863.470 ;
        RECT 1752.760 2802.010 1752.900 2863.150 ;
        RECT 1752.760 2801.870 1753.360 2802.010 ;
        RECT 1753.220 2767.590 1753.360 2801.870 ;
        RECT 1753.160 2767.270 1753.420 2767.590 ;
        RECT 1752.700 2766.590 1752.960 2766.910 ;
        RECT 1752.760 2714.550 1752.900 2766.590 ;
        RECT 1752.700 2714.230 1752.960 2714.550 ;
        RECT 1754.080 2714.230 1754.340 2714.550 ;
        RECT 1754.140 2623.430 1754.280 2714.230 ;
        RECT 1754.080 2623.110 1754.340 2623.430 ;
        RECT 1753.160 2622.090 1753.420 2622.410 ;
        RECT 1753.220 2573.450 1753.360 2622.090 ;
        RECT 1753.160 2573.130 1753.420 2573.450 ;
        RECT 1754.540 2573.130 1754.800 2573.450 ;
        RECT 1754.600 2512.590 1754.740 2573.130 ;
        RECT 1754.540 2512.270 1754.800 2512.590 ;
        RECT 1753.160 2511.930 1753.420 2512.250 ;
        RECT 1753.220 2477.230 1753.360 2511.930 ;
        RECT 1753.160 2476.910 1753.420 2477.230 ;
        RECT 1755.460 2476.570 1755.720 2476.890 ;
        RECT 1755.520 2415.205 1755.660 2476.570 ;
        RECT 1755.450 2414.835 1755.730 2415.205 ;
        RECT 1753.610 2414.155 1753.890 2414.525 ;
        RECT 1753.680 2366.245 1753.820 2414.155 ;
        RECT 1752.230 2365.875 1752.510 2366.245 ;
        RECT 1753.610 2365.875 1753.890 2366.245 ;
        RECT 1752.300 2291.330 1752.440 2365.875 ;
        RECT 1752.300 2291.190 1752.900 2291.330 ;
        RECT 1752.760 2285.210 1752.900 2291.190 ;
        RECT 1752.760 2285.070 1753.360 2285.210 ;
        RECT 1753.220 2277.220 1753.360 2285.070 ;
        RECT 1752.300 2277.080 1753.360 2277.220 ;
        RECT 1752.300 2263.450 1752.440 2277.080 ;
        RECT 1752.300 2263.310 1753.360 2263.450 ;
        RECT 1753.220 2197.490 1753.360 2263.310 ;
        RECT 1752.300 2197.350 1753.360 2197.490 ;
        RECT 1752.300 2136.290 1752.440 2197.350 ;
        RECT 1752.300 2136.150 1752.900 2136.290 ;
        RECT 1752.760 2090.730 1752.900 2136.150 ;
        RECT 1752.760 2090.590 1753.360 2090.730 ;
        RECT 1753.220 2043.640 1753.360 2090.590 ;
        RECT 1753.220 2043.500 1754.740 2043.640 ;
        RECT 1754.600 2042.710 1754.740 2043.500 ;
        RECT 1754.540 2042.390 1754.800 2042.710 ;
        RECT 1755.000 2041.030 1755.260 2041.350 ;
        RECT 1755.060 2027.490 1755.200 2041.030 ;
        RECT 1753.220 2027.350 1755.200 2027.490 ;
        RECT 1753.220 2007.770 1753.360 2027.350 ;
        RECT 1753.220 2007.630 1755.200 2007.770 ;
        RECT 1755.060 1973.350 1755.200 2007.630 ;
        RECT 1755.000 1973.030 1755.260 1973.350 ;
        RECT 1757.300 1973.205 1757.560 1973.350 ;
        RECT 1757.290 1972.835 1757.570 1973.205 ;
      LAYER via2 ;
        RECT 17.110 3339.680 17.390 3339.960 ;
        RECT 1755.450 2414.880 1755.730 2415.160 ;
        RECT 1753.610 2414.200 1753.890 2414.480 ;
        RECT 1752.230 2365.920 1752.510 2366.200 ;
        RECT 1753.610 2365.920 1753.890 2366.200 ;
        RECT 1757.290 1972.880 1757.570 1973.160 ;
      LAYER met3 ;
        RECT -4.800 3339.970 2.400 3340.420 ;
        RECT 17.085 3339.970 17.415 3339.985 ;
        RECT -4.800 3339.670 17.415 3339.970 ;
        RECT -4.800 3339.220 2.400 3339.670 ;
        RECT 17.085 3339.655 17.415 3339.670 ;
        RECT 1755.425 2415.170 1755.755 2415.185 ;
        RECT 1753.830 2414.870 1755.755 2415.170 ;
        RECT 1753.830 2414.505 1754.130 2414.870 ;
        RECT 1755.425 2414.855 1755.755 2414.870 ;
        RECT 1753.585 2414.190 1754.130 2414.505 ;
        RECT 1753.585 2414.175 1753.915 2414.190 ;
        RECT 1752.205 2366.210 1752.535 2366.225 ;
        RECT 1753.585 2366.210 1753.915 2366.225 ;
        RECT 1752.205 2365.910 1753.915 2366.210 ;
        RECT 1752.205 2365.895 1752.535 2365.910 ;
        RECT 1753.585 2365.895 1753.915 2365.910 ;
        RECT 1757.265 1973.170 1757.595 1973.185 ;
        RECT 1757.265 1972.855 1757.810 1973.170 ;
        RECT 1757.510 1972.495 1757.810 1972.855 ;
        RECT 1755.835 1971.895 1759.835 1972.495 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 3050.040 16.030 3050.100 ;
        RECT 31.350 3050.040 31.670 3050.100 ;
        RECT 15.710 3049.900 31.670 3050.040 ;
        RECT 15.710 3049.840 16.030 3049.900 ;
        RECT 31.350 3049.840 31.670 3049.900 ;
        RECT 31.350 2125.240 31.670 2125.300 ;
        RECT 706.170 2125.240 706.490 2125.300 ;
        RECT 31.350 2125.100 706.490 2125.240 ;
        RECT 31.350 2125.040 31.670 2125.100 ;
        RECT 706.170 2125.040 706.490 2125.100 ;
      LAYER via ;
        RECT 15.740 3049.840 16.000 3050.100 ;
        RECT 31.380 3049.840 31.640 3050.100 ;
        RECT 31.380 2125.040 31.640 2125.300 ;
        RECT 706.200 2125.040 706.460 2125.300 ;
      LAYER met2 ;
        RECT 15.730 3051.995 16.010 3052.365 ;
        RECT 15.800 3050.130 15.940 3051.995 ;
        RECT 15.740 3049.810 16.000 3050.130 ;
        RECT 31.380 3049.810 31.640 3050.130 ;
        RECT 31.440 2125.330 31.580 3049.810 ;
        RECT 31.380 2125.010 31.640 2125.330 ;
        RECT 706.200 2125.010 706.460 2125.330 ;
        RECT 706.260 2122.125 706.400 2125.010 ;
        RECT 706.190 2121.755 706.470 2122.125 ;
      LAYER via2 ;
        RECT 15.730 3052.040 16.010 3052.320 ;
        RECT 706.190 2121.800 706.470 2122.080 ;
      LAYER met3 ;
        RECT -4.800 3052.330 2.400 3052.780 ;
        RECT 15.705 3052.330 16.035 3052.345 ;
        RECT -4.800 3052.030 16.035 3052.330 ;
        RECT -4.800 3051.580 2.400 3052.030 ;
        RECT 15.705 3052.015 16.035 3052.030 ;
        RECT 706.165 2122.090 706.495 2122.105 ;
        RECT 715.810 2122.090 719.810 2122.095 ;
        RECT 706.165 2121.790 719.810 2122.090 ;
        RECT 706.165 2121.775 706.495 2121.790 ;
        RECT 715.810 2121.495 719.810 2121.790 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.470 1318.080 18.790 1318.140 ;
        RECT 914.550 1318.080 914.870 1318.140 ;
        RECT 18.470 1317.940 914.870 1318.080 ;
        RECT 18.470 1317.880 18.790 1317.940 ;
        RECT 914.550 1317.880 914.870 1317.940 ;
      LAYER via ;
        RECT 18.500 1317.880 18.760 1318.140 ;
        RECT 914.580 1317.880 914.840 1318.140 ;
      LAYER met2 ;
        RECT 18.490 2765.035 18.770 2765.405 ;
        RECT 18.560 1318.170 18.700 2765.035 ;
        RECT 914.620 1323.135 914.900 1327.135 ;
        RECT 914.640 1318.170 914.780 1323.135 ;
        RECT 18.500 1317.850 18.760 1318.170 ;
        RECT 914.580 1317.850 914.840 1318.170 ;
      LAYER via2 ;
        RECT 18.490 2765.080 18.770 2765.360 ;
      LAYER met3 ;
        RECT -4.800 2765.370 2.400 2765.820 ;
        RECT 18.465 2765.370 18.795 2765.385 ;
        RECT -4.800 2765.070 18.795 2765.370 ;
        RECT -4.800 2764.620 2.400 2765.070 ;
        RECT 18.465 2765.055 18.795 2765.070 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 20.310 2477.480 20.630 2477.540 ;
        RECT 993.670 2477.480 993.990 2477.540 ;
        RECT 20.310 2477.340 993.990 2477.480 ;
        RECT 20.310 2477.280 20.630 2477.340 ;
        RECT 993.670 2477.280 993.990 2477.340 ;
      LAYER via ;
        RECT 20.340 2477.280 20.600 2477.540 ;
        RECT 993.700 2477.280 993.960 2477.540 ;
      LAYER met2 ;
        RECT 20.330 2477.395 20.610 2477.765 ;
        RECT 20.340 2477.250 20.600 2477.395 ;
        RECT 993.700 2477.250 993.960 2477.570 ;
        RECT 993.760 2387.890 993.900 2477.250 ;
        RECT 993.760 2387.750 996.660 2387.890 ;
        RECT 996.520 2377.010 996.660 2387.750 ;
        RECT 999.260 2377.010 999.540 2377.880 ;
        RECT 996.520 2376.870 999.540 2377.010 ;
        RECT 999.260 2373.880 999.540 2376.870 ;
      LAYER via2 ;
        RECT 20.330 2477.440 20.610 2477.720 ;
      LAYER met3 ;
        RECT -4.800 2477.730 2.400 2478.180 ;
        RECT 20.305 2477.730 20.635 2477.745 ;
        RECT -4.800 2477.430 20.635 2477.730 ;
        RECT -4.800 2476.980 2.400 2477.430 ;
        RECT 20.305 2477.415 20.635 2477.430 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.930 1318.760 19.250 1318.820 ;
        RECT 937.550 1318.760 937.870 1318.820 ;
        RECT 18.930 1318.620 937.870 1318.760 ;
        RECT 18.930 1318.560 19.250 1318.620 ;
        RECT 937.550 1318.560 937.870 1318.620 ;
      LAYER via ;
        RECT 18.960 1318.560 19.220 1318.820 ;
        RECT 937.580 1318.560 937.840 1318.820 ;
      LAYER met2 ;
        RECT 18.950 2189.755 19.230 2190.125 ;
        RECT 19.020 1318.850 19.160 2189.755 ;
        RECT 937.620 1323.135 937.900 1327.135 ;
        RECT 937.640 1318.850 937.780 1323.135 ;
        RECT 18.960 1318.530 19.220 1318.850 ;
        RECT 937.580 1318.530 937.840 1318.850 ;
      LAYER via2 ;
        RECT 18.950 2189.800 19.230 2190.080 ;
      LAYER met3 ;
        RECT -4.800 2190.090 2.400 2190.540 ;
        RECT 18.925 2190.090 19.255 2190.105 ;
        RECT -4.800 2189.790 19.255 2190.090 ;
        RECT -4.800 2189.340 2.400 2189.790 ;
        RECT 18.925 2189.775 19.255 2189.790 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 19.850 1842.360 20.170 1842.420 ;
        RECT 696.970 1842.360 697.290 1842.420 ;
        RECT 19.850 1842.220 697.290 1842.360 ;
        RECT 19.850 1842.160 20.170 1842.220 ;
        RECT 696.970 1842.160 697.290 1842.220 ;
      LAYER via ;
        RECT 19.880 1842.160 20.140 1842.420 ;
        RECT 697.000 1842.160 697.260 1842.420 ;
      LAYER met2 ;
        RECT 19.870 1902.795 20.150 1903.165 ;
        RECT 19.940 1842.450 20.080 1902.795 ;
        RECT 19.880 1842.130 20.140 1842.450 ;
        RECT 697.000 1842.130 697.260 1842.450 ;
        RECT 697.060 1840.605 697.200 1842.130 ;
        RECT 696.990 1840.235 697.270 1840.605 ;
      LAYER via2 ;
        RECT 19.870 1902.840 20.150 1903.120 ;
        RECT 696.990 1840.280 697.270 1840.560 ;
      LAYER met3 ;
        RECT -4.800 1903.130 2.400 1903.580 ;
        RECT 19.845 1903.130 20.175 1903.145 ;
        RECT -4.800 1902.830 20.175 1903.130 ;
        RECT -4.800 1902.380 2.400 1902.830 ;
        RECT 19.845 1902.815 20.175 1902.830 ;
        RECT 696.965 1840.570 697.295 1840.585 ;
        RECT 715.810 1840.570 719.810 1840.575 ;
        RECT 696.965 1840.270 719.810 1840.570 ;
        RECT 696.965 1840.255 697.295 1840.270 ;
        RECT 715.810 1839.975 719.810 1840.270 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1772.910 2339.440 1773.230 2339.500 ;
        RECT 1797.290 2339.440 1797.610 2339.500 ;
        RECT 1772.910 2339.300 1797.610 2339.440 ;
        RECT 1772.910 2339.240 1773.230 2339.300 ;
        RECT 1797.290 2339.240 1797.610 2339.300 ;
        RECT 1797.290 620.740 1797.610 620.800 ;
        RECT 2900.830 620.740 2901.150 620.800 ;
        RECT 1797.290 620.600 2901.150 620.740 ;
        RECT 1797.290 620.540 1797.610 620.600 ;
        RECT 2900.830 620.540 2901.150 620.600 ;
      LAYER via ;
        RECT 1772.940 2339.240 1773.200 2339.500 ;
        RECT 1797.320 2339.240 1797.580 2339.500 ;
        RECT 1797.320 620.540 1797.580 620.800 ;
        RECT 2900.860 620.540 2901.120 620.800 ;
      LAYER met2 ;
        RECT 1772.930 2339.355 1773.210 2339.725 ;
        RECT 1772.940 2339.210 1773.200 2339.355 ;
        RECT 1797.320 2339.210 1797.580 2339.530 ;
        RECT 1797.380 620.830 1797.520 2339.210 ;
        RECT 1797.320 620.510 1797.580 620.830 ;
        RECT 2900.860 620.510 2901.120 620.830 ;
        RECT 2900.920 615.925 2901.060 620.510 ;
        RECT 2900.850 615.555 2901.130 615.925 ;
      LAYER via2 ;
        RECT 1772.930 2339.400 1773.210 2339.680 ;
        RECT 2900.850 615.600 2901.130 615.880 ;
      LAYER met3 ;
        RECT 1755.835 2339.690 1759.835 2339.695 ;
        RECT 1772.905 2339.690 1773.235 2339.705 ;
        RECT 1755.835 2339.390 1773.235 2339.690 ;
        RECT 1755.835 2339.095 1759.835 2339.390 ;
        RECT 1772.905 2339.375 1773.235 2339.390 ;
        RECT 2900.825 615.890 2901.155 615.905 ;
        RECT 2917.600 615.890 2924.800 616.340 ;
        RECT 2900.825 615.590 2924.800 615.890 ;
        RECT 2900.825 615.575 2901.155 615.590 ;
        RECT 2917.600 615.140 2924.800 615.590 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 688.230 2386.020 688.550 2386.080 ;
        RECT 1196.070 2386.020 1196.390 2386.080 ;
        RECT 688.230 2385.880 1196.390 2386.020 ;
        RECT 688.230 2385.820 688.550 2385.880 ;
        RECT 1196.070 2385.820 1196.390 2385.880 ;
        RECT 16.170 1621.360 16.490 1621.420 ;
        RECT 688.230 1621.360 688.550 1621.420 ;
        RECT 16.170 1621.220 688.550 1621.360 ;
        RECT 16.170 1621.160 16.490 1621.220 ;
        RECT 688.230 1621.160 688.550 1621.220 ;
      LAYER via ;
        RECT 688.260 2385.820 688.520 2386.080 ;
        RECT 1196.100 2385.820 1196.360 2386.080 ;
        RECT 16.200 1621.160 16.460 1621.420 ;
        RECT 688.260 1621.160 688.520 1621.420 ;
      LAYER met2 ;
        RECT 688.260 2385.790 688.520 2386.110 ;
        RECT 1196.100 2385.790 1196.360 2386.110 ;
        RECT 688.320 1621.450 688.460 2385.790 ;
        RECT 1196.160 2377.880 1196.300 2385.790 ;
        RECT 1196.140 2373.880 1196.420 2377.880 ;
        RECT 16.200 1621.130 16.460 1621.450 ;
        RECT 688.260 1621.130 688.520 1621.450 ;
        RECT 16.260 1615.525 16.400 1621.130 ;
        RECT 16.190 1615.155 16.470 1615.525 ;
      LAYER via2 ;
        RECT 16.190 1615.200 16.470 1615.480 ;
      LAYER met3 ;
        RECT -4.800 1615.490 2.400 1615.940 ;
        RECT 16.165 1615.490 16.495 1615.505 ;
        RECT -4.800 1615.190 16.495 1615.490 ;
        RECT -4.800 1614.740 2.400 1615.190 ;
        RECT 16.165 1615.175 16.495 1615.190 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1752.745 1330.165 1752.915 1331.695 ;
        RECT 1756.885 1330.165 1757.055 1331.695 ;
      LAYER mcon ;
        RECT 1752.745 1331.525 1752.915 1331.695 ;
        RECT 1756.885 1331.525 1757.055 1331.695 ;
      LAYER met1 ;
        RECT 1757.270 1343.240 1757.590 1343.300 ;
        RECT 1759.110 1343.240 1759.430 1343.300 ;
        RECT 1757.270 1343.100 1759.430 1343.240 ;
        RECT 1757.270 1343.040 1757.590 1343.100 ;
        RECT 1759.110 1343.040 1759.430 1343.100 ;
        RECT 16.170 1331.680 16.490 1331.740 ;
        RECT 1752.685 1331.680 1752.975 1331.725 ;
        RECT 16.170 1331.540 1752.975 1331.680 ;
        RECT 16.170 1331.480 16.490 1331.540 ;
        RECT 1752.685 1331.495 1752.975 1331.540 ;
        RECT 1756.825 1331.680 1757.115 1331.725 ;
        RECT 1757.270 1331.680 1757.590 1331.740 ;
        RECT 1756.825 1331.540 1757.590 1331.680 ;
        RECT 1756.825 1331.495 1757.115 1331.540 ;
        RECT 1757.270 1331.480 1757.590 1331.540 ;
        RECT 1752.685 1330.320 1752.975 1330.365 ;
        RECT 1756.825 1330.320 1757.115 1330.365 ;
        RECT 1752.685 1330.180 1757.115 1330.320 ;
        RECT 1752.685 1330.135 1752.975 1330.180 ;
        RECT 1756.825 1330.135 1757.115 1330.180 ;
      LAYER via ;
        RECT 1757.300 1343.040 1757.560 1343.300 ;
        RECT 1759.140 1343.040 1759.400 1343.300 ;
        RECT 16.200 1331.480 16.460 1331.740 ;
        RECT 1757.300 1331.480 1757.560 1331.740 ;
      LAYER met2 ;
        RECT 1759.130 1483.915 1759.410 1484.285 ;
        RECT 16.190 1400.275 16.470 1400.645 ;
        RECT 16.260 1331.770 16.400 1400.275 ;
        RECT 1759.200 1343.330 1759.340 1483.915 ;
        RECT 1757.300 1343.010 1757.560 1343.330 ;
        RECT 1759.140 1343.010 1759.400 1343.330 ;
        RECT 1757.360 1331.770 1757.500 1343.010 ;
        RECT 16.200 1331.450 16.460 1331.770 ;
        RECT 1757.300 1331.450 1757.560 1331.770 ;
      LAYER via2 ;
        RECT 1759.130 1483.960 1759.410 1484.240 ;
        RECT 16.190 1400.320 16.470 1400.600 ;
      LAYER met3 ;
        RECT 1755.835 1485.015 1759.835 1485.615 ;
        RECT 1759.350 1484.265 1759.650 1485.015 ;
        RECT 1759.105 1483.950 1759.650 1484.265 ;
        RECT 1759.105 1483.935 1759.435 1483.950 ;
        RECT -4.800 1400.610 2.400 1401.060 ;
        RECT 16.165 1400.610 16.495 1400.625 ;
        RECT -4.800 1400.310 16.495 1400.610 ;
        RECT -4.800 1399.860 2.400 1400.310 ;
        RECT 16.165 1400.295 16.495 1400.310 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 699.270 2385.340 699.590 2385.400 ;
        RECT 1374.550 2385.340 1374.870 2385.400 ;
        RECT 699.270 2385.200 1374.870 2385.340 ;
        RECT 699.270 2385.140 699.590 2385.200 ;
        RECT 1374.550 2385.140 1374.870 2385.200 ;
        RECT 16.170 1186.840 16.490 1186.900 ;
        RECT 699.270 1186.840 699.590 1186.900 ;
        RECT 16.170 1186.700 699.590 1186.840 ;
        RECT 16.170 1186.640 16.490 1186.700 ;
        RECT 699.270 1186.640 699.590 1186.700 ;
      LAYER via ;
        RECT 699.300 2385.140 699.560 2385.400 ;
        RECT 1374.580 2385.140 1374.840 2385.400 ;
        RECT 16.200 1186.640 16.460 1186.900 ;
        RECT 699.300 1186.640 699.560 1186.900 ;
      LAYER met2 ;
        RECT 699.300 2385.110 699.560 2385.430 ;
        RECT 1374.580 2385.110 1374.840 2385.430 ;
        RECT 699.360 1393.845 699.500 2385.110 ;
        RECT 1374.640 2377.880 1374.780 2385.110 ;
        RECT 1374.620 2373.880 1374.900 2377.880 ;
        RECT 699.290 1393.475 699.570 1393.845 ;
        RECT 699.290 1390.755 699.570 1391.125 ;
        RECT 699.360 1186.930 699.500 1390.755 ;
        RECT 16.200 1186.610 16.460 1186.930 ;
        RECT 699.300 1186.610 699.560 1186.930 ;
        RECT 16.260 1185.085 16.400 1186.610 ;
        RECT 16.190 1184.715 16.470 1185.085 ;
      LAYER via2 ;
        RECT 699.290 1393.520 699.570 1393.800 ;
        RECT 699.290 1390.800 699.570 1391.080 ;
        RECT 16.190 1184.760 16.470 1185.040 ;
      LAYER met3 ;
        RECT 699.265 1393.810 699.595 1393.825 ;
        RECT 699.265 1393.495 699.810 1393.810 ;
        RECT 699.510 1391.105 699.810 1393.495 ;
        RECT 699.265 1390.790 699.810 1391.105 ;
        RECT 699.265 1390.775 699.595 1390.790 ;
        RECT -4.800 1185.050 2.400 1185.500 ;
        RECT 16.165 1185.050 16.495 1185.065 ;
        RECT -4.800 1184.750 16.495 1185.050 ;
        RECT -4.800 1184.300 2.400 1184.750 ;
        RECT 16.165 1184.735 16.495 1184.750 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 700.650 2385.680 700.970 2385.740 ;
        RECT 1155.590 2385.680 1155.910 2385.740 ;
        RECT 700.650 2385.540 1155.910 2385.680 ;
        RECT 700.650 2385.480 700.970 2385.540 ;
        RECT 1155.590 2385.480 1155.910 2385.540 ;
        RECT 18.010 972.640 18.330 972.700 ;
        RECT 700.650 972.640 700.970 972.700 ;
        RECT 18.010 972.500 700.970 972.640 ;
        RECT 18.010 972.440 18.330 972.500 ;
        RECT 700.650 972.440 700.970 972.500 ;
      LAYER via ;
        RECT 700.680 2385.480 700.940 2385.740 ;
        RECT 1155.620 2385.480 1155.880 2385.740 ;
        RECT 18.040 972.440 18.300 972.700 ;
        RECT 700.680 972.440 700.940 972.700 ;
      LAYER met2 ;
        RECT 700.680 2385.450 700.940 2385.770 ;
        RECT 1155.620 2385.450 1155.880 2385.770 ;
        RECT 700.740 972.730 700.880 2385.450 ;
        RECT 1155.680 2377.880 1155.820 2385.450 ;
        RECT 1155.660 2373.880 1155.940 2377.880 ;
        RECT 18.040 972.410 18.300 972.730 ;
        RECT 700.680 972.410 700.940 972.730 ;
        RECT 18.100 969.525 18.240 972.410 ;
        RECT 18.030 969.155 18.310 969.525 ;
      LAYER via2 ;
        RECT 18.030 969.200 18.310 969.480 ;
      LAYER met3 ;
        RECT -4.800 969.490 2.400 969.940 ;
        RECT 18.005 969.490 18.335 969.505 ;
        RECT -4.800 969.190 18.335 969.490 ;
        RECT -4.800 968.740 2.400 969.190 ;
        RECT 18.005 969.175 18.335 969.190 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.550 2378.540 17.870 2378.600 ;
        RECT 918.230 2378.540 918.550 2378.600 ;
        RECT 17.550 2378.400 918.550 2378.540 ;
        RECT 17.550 2378.340 17.870 2378.400 ;
        RECT 918.230 2378.340 918.550 2378.400 ;
      LAYER via ;
        RECT 17.580 2378.340 17.840 2378.600 ;
        RECT 918.260 2378.340 918.520 2378.600 ;
      LAYER met2 ;
        RECT 17.580 2378.310 17.840 2378.630 ;
        RECT 918.260 2378.310 918.520 2378.630 ;
        RECT 17.640 753.965 17.780 2378.310 ;
        RECT 918.320 2377.880 918.460 2378.310 ;
        RECT 918.300 2373.880 918.580 2377.880 ;
        RECT 17.570 753.595 17.850 753.965 ;
      LAYER via2 ;
        RECT 17.570 753.640 17.850 753.920 ;
      LAYER met3 ;
        RECT -4.800 753.930 2.400 754.380 ;
        RECT 17.545 753.930 17.875 753.945 ;
        RECT -4.800 753.630 17.875 753.930 ;
        RECT -4.800 753.180 2.400 753.630 ;
        RECT 17.545 753.615 17.875 753.630 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 18.490 1272.435 18.770 1272.805 ;
        RECT 18.560 538.405 18.700 1272.435 ;
        RECT 18.490 538.035 18.770 538.405 ;
      LAYER via2 ;
        RECT 18.490 1272.480 18.770 1272.760 ;
        RECT 18.490 538.080 18.770 538.360 ;
      LAYER met3 ;
        RECT 1755.835 1535.335 1759.835 1535.935 ;
        RECT 1758.430 1533.220 1758.730 1535.335 ;
        RECT 1758.390 1532.900 1758.770 1533.220 ;
        RECT 18.465 1272.770 18.795 1272.785 ;
        RECT 1758.390 1272.770 1758.770 1272.780 ;
        RECT 18.465 1272.470 1758.770 1272.770 ;
        RECT 18.465 1272.455 18.795 1272.470 ;
        RECT 1758.390 1272.460 1758.770 1272.470 ;
        RECT -4.800 538.370 2.400 538.820 ;
        RECT 18.465 538.370 18.795 538.385 ;
        RECT -4.800 538.070 18.795 538.370 ;
        RECT -4.800 537.620 2.400 538.070 ;
        RECT 18.465 538.055 18.795 538.070 ;
      LAYER via3 ;
        RECT 1758.420 1532.900 1758.740 1533.220 ;
        RECT 1758.420 1272.460 1758.740 1272.780 ;
      LAYER met4 ;
        RECT 1758.415 1532.895 1758.745 1533.225 ;
        RECT 1758.430 1272.785 1758.730 1532.895 ;
        RECT 1758.415 1272.455 1758.745 1272.785 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 51.590 1946.060 51.910 1946.120 ;
        RECT 706.170 1946.060 706.490 1946.120 ;
        RECT 51.590 1945.920 706.490 1946.060 ;
        RECT 51.590 1945.860 51.910 1945.920 ;
        RECT 706.170 1945.860 706.490 1945.920 ;
        RECT 17.550 324.260 17.870 324.320 ;
        RECT 51.590 324.260 51.910 324.320 ;
        RECT 17.550 324.120 51.910 324.260 ;
        RECT 17.550 324.060 17.870 324.120 ;
        RECT 51.590 324.060 51.910 324.120 ;
      LAYER via ;
        RECT 51.620 1945.860 51.880 1946.120 ;
        RECT 706.200 1945.860 706.460 1946.120 ;
        RECT 17.580 324.060 17.840 324.320 ;
        RECT 51.620 324.060 51.880 324.320 ;
      LAYER met2 ;
        RECT 706.190 1951.755 706.470 1952.125 ;
        RECT 706.260 1946.150 706.400 1951.755 ;
        RECT 51.620 1945.830 51.880 1946.150 ;
        RECT 706.200 1945.830 706.460 1946.150 ;
        RECT 51.680 324.350 51.820 1945.830 ;
        RECT 17.580 324.030 17.840 324.350 ;
        RECT 51.620 324.030 51.880 324.350 ;
        RECT 17.640 322.845 17.780 324.030 ;
        RECT 17.570 322.475 17.850 322.845 ;
      LAYER via2 ;
        RECT 706.190 1951.800 706.470 1952.080 ;
        RECT 17.570 322.520 17.850 322.800 ;
      LAYER met3 ;
        RECT 706.165 1952.090 706.495 1952.105 ;
        RECT 715.810 1952.090 719.810 1952.095 ;
        RECT 706.165 1951.790 719.810 1952.090 ;
        RECT 706.165 1951.775 706.495 1951.790 ;
        RECT 715.810 1951.495 719.810 1951.790 ;
        RECT -4.800 322.810 2.400 323.260 ;
        RECT 17.545 322.810 17.875 322.825 ;
        RECT -4.800 322.510 17.875 322.810 ;
        RECT -4.800 322.060 2.400 322.510 ;
        RECT 17.545 322.495 17.875 322.510 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1756.370 2320.315 1756.650 2320.685 ;
        RECT 1756.440 1391.125 1756.580 2320.315 ;
        RECT 1756.370 1390.755 1756.650 1391.125 ;
        RECT 1757.750 1299.635 1758.030 1300.005 ;
        RECT 1757.820 1249.005 1757.960 1299.635 ;
        RECT 1757.750 1248.635 1758.030 1249.005 ;
        RECT 1756.830 813.435 1757.110 813.805 ;
        RECT 1756.900 766.885 1757.040 813.435 ;
        RECT 1756.830 766.515 1757.110 766.885 ;
        RECT 1756.370 765.155 1756.650 765.525 ;
        RECT 1756.440 717.925 1756.580 765.155 ;
        RECT 1756.370 717.555 1756.650 717.925 ;
        RECT 1757.750 709.395 1758.030 709.765 ;
        RECT 1757.820 662.845 1757.960 709.395 ;
        RECT 1757.750 662.475 1758.030 662.845 ;
        RECT 1757.290 613.515 1757.570 613.885 ;
        RECT 1757.360 566.965 1757.500 613.515 ;
        RECT 1757.290 566.595 1757.570 566.965 ;
        RECT 1757.750 516.955 1758.030 517.325 ;
        RECT 1757.820 470.405 1757.960 516.955 ;
        RECT 1757.750 470.035 1758.030 470.405 ;
        RECT 1757.750 426.515 1758.030 426.885 ;
        RECT 1757.820 380.645 1757.960 426.515 ;
        RECT 1757.750 380.275 1758.030 380.645 ;
      LAYER via2 ;
        RECT 1756.370 2320.360 1756.650 2320.640 ;
        RECT 1756.370 1390.800 1756.650 1391.080 ;
        RECT 1757.750 1299.680 1758.030 1299.960 ;
        RECT 1757.750 1248.680 1758.030 1248.960 ;
        RECT 1756.830 813.480 1757.110 813.760 ;
        RECT 1756.830 766.560 1757.110 766.840 ;
        RECT 1756.370 765.200 1756.650 765.480 ;
        RECT 1756.370 717.600 1756.650 717.880 ;
        RECT 1757.750 709.440 1758.030 709.720 ;
        RECT 1757.750 662.520 1758.030 662.800 ;
        RECT 1757.290 613.560 1757.570 613.840 ;
        RECT 1757.290 566.640 1757.570 566.920 ;
        RECT 1757.750 517.000 1758.030 517.280 ;
        RECT 1757.750 470.080 1758.030 470.360 ;
        RECT 1757.750 426.560 1758.030 426.840 ;
        RECT 1757.750 380.320 1758.030 380.600 ;
      LAYER met3 ;
        RECT 1755.835 2322.775 1759.835 2323.375 ;
        RECT 1756.590 2320.665 1756.890 2322.775 ;
        RECT 1756.345 2320.350 1756.890 2320.665 ;
        RECT 1756.345 2320.335 1756.675 2320.350 ;
        RECT 1756.345 1391.090 1756.675 1391.105 ;
        RECT 1763.910 1391.090 1764.290 1391.100 ;
        RECT 1756.345 1390.790 1764.290 1391.090 ;
        RECT 1756.345 1390.775 1756.675 1390.790 ;
        RECT 1763.910 1390.780 1764.290 1390.790 ;
        RECT 1763.910 1367.290 1764.290 1367.300 ;
        RECT 1757.510 1366.990 1764.290 1367.290 ;
        RECT 1757.510 1366.620 1757.810 1366.990 ;
        RECT 1763.910 1366.980 1764.290 1366.990 ;
        RECT 1757.470 1366.300 1757.850 1366.620 ;
        RECT 1757.725 1299.980 1758.055 1299.985 ;
        RECT 1757.470 1299.970 1758.055 1299.980 ;
        RECT 1757.270 1299.670 1758.055 1299.970 ;
        RECT 1757.470 1299.660 1758.055 1299.670 ;
        RECT 1757.725 1299.655 1758.055 1299.660 ;
        RECT 1757.725 1248.980 1758.055 1248.985 ;
        RECT 1757.470 1248.970 1758.055 1248.980 ;
        RECT 1757.270 1248.670 1758.055 1248.970 ;
        RECT 1757.470 1248.660 1758.055 1248.670 ;
        RECT 1757.725 1248.655 1758.055 1248.660 ;
        RECT 1756.805 813.770 1757.135 813.785 ;
        RECT 1757.470 813.770 1757.850 813.780 ;
        RECT 1756.805 813.470 1757.850 813.770 ;
        RECT 1756.805 813.455 1757.135 813.470 ;
        RECT 1757.470 813.460 1757.850 813.470 ;
        RECT 1756.805 766.860 1757.135 766.865 ;
        RECT 1756.550 766.850 1757.135 766.860 ;
        RECT 1756.350 766.550 1757.135 766.850 ;
        RECT 1756.550 766.540 1757.135 766.550 ;
        RECT 1756.805 766.535 1757.135 766.540 ;
        RECT 1756.345 765.500 1756.675 765.505 ;
        RECT 1756.345 765.490 1756.930 765.500 ;
        RECT 1756.120 765.190 1756.930 765.490 ;
        RECT 1756.345 765.180 1756.930 765.190 ;
        RECT 1756.345 765.175 1756.675 765.180 ;
        RECT 1756.345 717.900 1756.675 717.905 ;
        RECT 1756.345 717.890 1756.930 717.900 ;
        RECT 1756.345 717.590 1757.130 717.890 ;
        RECT 1756.345 717.580 1756.930 717.590 ;
        RECT 1756.345 717.575 1756.675 717.580 ;
        RECT 1756.550 710.100 1756.930 710.420 ;
        RECT 1756.590 709.730 1756.890 710.100 ;
        RECT 1757.725 709.730 1758.055 709.745 ;
        RECT 1756.590 709.430 1758.055 709.730 ;
        RECT 1757.725 709.415 1758.055 709.430 ;
        RECT 1757.725 662.820 1758.055 662.825 ;
        RECT 1757.470 662.810 1758.055 662.820 ;
        RECT 1757.470 662.510 1758.280 662.810 ;
        RECT 1757.470 662.500 1758.055 662.510 ;
        RECT 1757.725 662.495 1758.055 662.500 ;
        RECT 1757.265 613.860 1757.595 613.865 ;
        RECT 1757.265 613.850 1757.850 613.860 ;
        RECT 1757.040 613.550 1757.850 613.850 ;
        RECT 1757.265 613.540 1757.850 613.550 ;
        RECT 1757.265 613.535 1757.595 613.540 ;
        RECT 1757.265 566.930 1757.595 566.945 ;
        RECT 1757.265 566.615 1757.810 566.930 ;
        RECT 1757.510 566.260 1757.810 566.615 ;
        RECT 1757.470 565.940 1757.850 566.260 ;
        RECT 1757.725 517.300 1758.055 517.305 ;
        RECT 1757.470 517.290 1758.055 517.300 ;
        RECT 1757.470 516.990 1758.280 517.290 ;
        RECT 1757.470 516.980 1758.055 516.990 ;
        RECT 1757.725 516.975 1758.055 516.980 ;
        RECT 1757.725 470.370 1758.055 470.385 ;
        RECT 1757.510 470.055 1758.055 470.370 ;
        RECT 1757.510 469.700 1757.810 470.055 ;
        RECT 1757.470 469.380 1757.850 469.700 ;
        RECT 1757.470 428.890 1757.850 428.900 ;
        RECT 1757.470 428.590 1758.730 428.890 ;
        RECT 1757.470 428.580 1757.850 428.590 ;
        RECT 1757.725 426.850 1758.055 426.865 ;
        RECT 1758.430 426.850 1758.730 428.590 ;
        RECT 1757.725 426.550 1758.730 426.850 ;
        RECT 1757.725 426.535 1758.055 426.550 ;
        RECT 1757.725 380.610 1758.055 380.625 ;
        RECT 1757.510 380.295 1758.055 380.610 ;
        RECT 1757.510 379.940 1757.810 380.295 ;
        RECT 1757.470 379.620 1757.850 379.940 ;
        RECT 1757.470 109.970 1757.850 109.980 ;
        RECT 3.070 109.670 1757.850 109.970 ;
        RECT -4.800 107.250 2.400 107.700 ;
        RECT 3.070 107.250 3.370 109.670 ;
        RECT 1757.470 109.660 1757.850 109.670 ;
        RECT -4.800 106.950 3.370 107.250 ;
        RECT -4.800 106.500 2.400 106.950 ;
      LAYER via3 ;
        RECT 1763.940 1390.780 1764.260 1391.100 ;
        RECT 1763.940 1366.980 1764.260 1367.300 ;
        RECT 1757.500 1366.300 1757.820 1366.620 ;
        RECT 1757.500 1299.660 1757.820 1299.980 ;
        RECT 1757.500 1248.660 1757.820 1248.980 ;
        RECT 1757.500 813.460 1757.820 813.780 ;
        RECT 1756.580 766.540 1756.900 766.860 ;
        RECT 1756.580 765.180 1756.900 765.500 ;
        RECT 1756.580 717.580 1756.900 717.900 ;
        RECT 1756.580 710.100 1756.900 710.420 ;
        RECT 1757.500 662.500 1757.820 662.820 ;
        RECT 1757.500 613.540 1757.820 613.860 ;
        RECT 1757.500 565.940 1757.820 566.260 ;
        RECT 1757.500 516.980 1757.820 517.300 ;
        RECT 1757.500 469.380 1757.820 469.700 ;
        RECT 1757.500 428.580 1757.820 428.900 ;
        RECT 1757.500 379.620 1757.820 379.940 ;
        RECT 1757.500 109.660 1757.820 109.980 ;
      LAYER met4 ;
        RECT 1763.935 1390.775 1764.265 1391.105 ;
        RECT 1763.950 1367.305 1764.250 1390.775 ;
        RECT 1763.935 1366.975 1764.265 1367.305 ;
        RECT 1757.495 1366.295 1757.825 1366.625 ;
        RECT 1757.510 1299.985 1757.810 1366.295 ;
        RECT 1757.495 1299.655 1757.825 1299.985 ;
        RECT 1757.495 1248.655 1757.825 1248.985 ;
        RECT 1757.510 813.785 1757.810 1248.655 ;
        RECT 1757.495 813.455 1757.825 813.785 ;
        RECT 1756.575 766.535 1756.905 766.865 ;
        RECT 1756.590 765.505 1756.890 766.535 ;
        RECT 1756.575 765.175 1756.905 765.505 ;
        RECT 1756.575 717.575 1756.905 717.905 ;
        RECT 1756.590 710.425 1756.890 717.575 ;
        RECT 1756.575 710.095 1756.905 710.425 ;
        RECT 1757.495 662.495 1757.825 662.825 ;
        RECT 1757.510 613.865 1757.810 662.495 ;
        RECT 1757.495 613.535 1757.825 613.865 ;
        RECT 1757.495 565.935 1757.825 566.265 ;
        RECT 1757.510 517.305 1757.810 565.935 ;
        RECT 1757.495 516.975 1757.825 517.305 ;
        RECT 1757.495 469.375 1757.825 469.705 ;
        RECT 1757.510 428.905 1757.810 469.375 ;
        RECT 1757.495 428.575 1757.825 428.905 ;
        RECT 1757.495 379.615 1757.825 379.945 ;
        RECT 1757.510 304.450 1757.810 379.615 ;
        RECT 1757.510 304.150 1758.500 304.450 ;
        RECT 1758.200 303.090 1758.500 304.150 ;
        RECT 1757.510 302.790 1758.500 303.090 ;
        RECT 1757.510 109.985 1757.810 302.790 ;
        RECT 1757.495 109.655 1757.825 109.985 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1392.030 2386.700 1392.350 2386.760 ;
        RECT 1783.950 2386.700 1784.270 2386.760 ;
        RECT 1392.030 2386.560 1784.270 2386.700 ;
        RECT 1392.030 2386.500 1392.350 2386.560 ;
        RECT 1783.950 2386.500 1784.270 2386.560 ;
        RECT 1783.950 855.340 1784.270 855.400 ;
        RECT 2900.830 855.340 2901.150 855.400 ;
        RECT 1783.950 855.200 2901.150 855.340 ;
        RECT 1783.950 855.140 1784.270 855.200 ;
        RECT 2900.830 855.140 2901.150 855.200 ;
      LAYER via ;
        RECT 1392.060 2386.500 1392.320 2386.760 ;
        RECT 1783.980 2386.500 1784.240 2386.760 ;
        RECT 1783.980 855.140 1784.240 855.400 ;
        RECT 2900.860 855.140 2901.120 855.400 ;
      LAYER met2 ;
        RECT 1392.060 2386.470 1392.320 2386.790 ;
        RECT 1783.980 2386.470 1784.240 2386.790 ;
        RECT 1392.120 2377.880 1392.260 2386.470 ;
        RECT 1392.100 2373.880 1392.380 2377.880 ;
        RECT 1784.040 855.430 1784.180 2386.470 ;
        RECT 1783.980 855.110 1784.240 855.430 ;
        RECT 2900.860 855.110 2901.120 855.430 ;
        RECT 2900.920 850.525 2901.060 855.110 ;
        RECT 2900.850 850.155 2901.130 850.525 ;
      LAYER via2 ;
        RECT 2900.850 850.200 2901.130 850.480 ;
      LAYER met3 ;
        RECT 2900.825 850.490 2901.155 850.505 ;
        RECT 2917.600 850.490 2924.800 850.940 ;
        RECT 2900.825 850.190 2924.800 850.490 ;
        RECT 2900.825 850.175 2901.155 850.190 ;
        RECT 2917.600 849.740 2924.800 850.190 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1772.910 1669.980 1773.230 1670.040 ;
        RECT 1778.430 1669.980 1778.750 1670.040 ;
        RECT 1772.910 1669.840 1778.750 1669.980 ;
        RECT 1772.910 1669.780 1773.230 1669.840 ;
        RECT 1778.430 1669.780 1778.750 1669.840 ;
        RECT 1778.430 1089.940 1778.750 1090.000 ;
        RECT 2900.830 1089.940 2901.150 1090.000 ;
        RECT 1778.430 1089.800 2901.150 1089.940 ;
        RECT 1778.430 1089.740 1778.750 1089.800 ;
        RECT 2900.830 1089.740 2901.150 1089.800 ;
      LAYER via ;
        RECT 1772.940 1669.780 1773.200 1670.040 ;
        RECT 1778.460 1669.780 1778.720 1670.040 ;
        RECT 1778.460 1089.740 1778.720 1090.000 ;
        RECT 2900.860 1089.740 2901.120 1090.000 ;
      LAYER met2 ;
        RECT 1772.930 1672.955 1773.210 1673.325 ;
        RECT 1773.000 1670.070 1773.140 1672.955 ;
        RECT 1772.940 1669.750 1773.200 1670.070 ;
        RECT 1778.460 1669.750 1778.720 1670.070 ;
        RECT 1778.520 1090.030 1778.660 1669.750 ;
        RECT 1778.460 1089.710 1778.720 1090.030 ;
        RECT 2900.860 1089.710 2901.120 1090.030 ;
        RECT 2900.920 1085.125 2901.060 1089.710 ;
        RECT 2900.850 1084.755 2901.130 1085.125 ;
      LAYER via2 ;
        RECT 1772.930 1673.000 1773.210 1673.280 ;
        RECT 2900.850 1084.800 2901.130 1085.080 ;
      LAYER met3 ;
        RECT 1755.835 1673.290 1759.835 1673.295 ;
        RECT 1772.905 1673.290 1773.235 1673.305 ;
        RECT 1755.835 1672.990 1773.235 1673.290 ;
        RECT 1755.835 1672.695 1759.835 1672.990 ;
        RECT 1772.905 1672.975 1773.235 1672.990 ;
        RECT 2900.825 1085.090 2901.155 1085.105 ;
        RECT 2917.600 1085.090 2924.800 1085.540 ;
        RECT 2900.825 1084.790 2924.800 1085.090 ;
        RECT 2900.825 1084.775 2901.155 1084.790 ;
        RECT 2917.600 1084.340 2924.800 1084.790 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 690.070 1898.800 690.390 1898.860 ;
        RECT 710.310 1898.800 710.630 1898.860 ;
        RECT 690.070 1898.660 710.630 1898.800 ;
        RECT 690.070 1898.600 690.390 1898.660 ;
        RECT 710.310 1898.600 710.630 1898.660 ;
        RECT 690.070 1324.540 690.390 1324.600 ;
        RECT 2900.830 1324.540 2901.150 1324.600 ;
        RECT 690.070 1324.400 2901.150 1324.540 ;
        RECT 690.070 1324.340 690.390 1324.400 ;
        RECT 2900.830 1324.340 2901.150 1324.400 ;
      LAYER via ;
        RECT 690.100 1898.600 690.360 1898.860 ;
        RECT 710.340 1898.600 710.600 1898.860 ;
        RECT 690.100 1324.340 690.360 1324.600 ;
        RECT 2900.860 1324.340 2901.120 1324.600 ;
      LAYER met2 ;
        RECT 710.330 1900.075 710.610 1900.445 ;
        RECT 710.400 1898.890 710.540 1900.075 ;
        RECT 690.100 1898.570 690.360 1898.890 ;
        RECT 710.340 1898.570 710.600 1898.890 ;
        RECT 690.160 1393.845 690.300 1898.570 ;
        RECT 690.090 1393.475 690.370 1393.845 ;
        RECT 690.090 1390.755 690.370 1391.125 ;
        RECT 690.160 1324.630 690.300 1390.755 ;
        RECT 690.100 1324.310 690.360 1324.630 ;
        RECT 2900.860 1324.310 2901.120 1324.630 ;
        RECT 2900.920 1319.725 2901.060 1324.310 ;
        RECT 2900.850 1319.355 2901.130 1319.725 ;
      LAYER via2 ;
        RECT 710.330 1900.120 710.610 1900.400 ;
        RECT 690.090 1393.520 690.370 1393.800 ;
        RECT 690.090 1390.800 690.370 1391.080 ;
        RECT 2900.850 1319.400 2901.130 1319.680 ;
      LAYER met3 ;
        RECT 710.305 1900.410 710.635 1900.425 ;
        RECT 715.810 1900.410 719.810 1900.415 ;
        RECT 710.305 1900.110 719.810 1900.410 ;
        RECT 710.305 1900.095 710.635 1900.110 ;
        RECT 715.810 1899.815 719.810 1900.110 ;
        RECT 690.065 1393.810 690.395 1393.825 ;
        RECT 690.065 1393.495 690.610 1393.810 ;
        RECT 690.310 1391.105 690.610 1393.495 ;
        RECT 690.065 1390.790 690.610 1391.105 ;
        RECT 690.065 1390.775 690.395 1390.790 ;
        RECT 2900.825 1319.690 2901.155 1319.705 ;
        RECT 2917.600 1319.690 2924.800 1320.140 ;
        RECT 2900.825 1319.390 2924.800 1319.690 ;
        RECT 2900.825 1319.375 2901.155 1319.390 ;
        RECT 2917.600 1318.940 2924.800 1319.390 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1571.430 2380.920 1571.750 2380.980 ;
        RECT 2452.790 2380.920 2453.110 2380.980 ;
        RECT 1571.430 2380.780 2453.110 2380.920 ;
        RECT 1571.430 2380.720 1571.750 2380.780 ;
        RECT 2452.790 2380.720 2453.110 2380.780 ;
        RECT 2452.790 1559.140 2453.110 1559.200 ;
        RECT 2899.910 1559.140 2900.230 1559.200 ;
        RECT 2452.790 1559.000 2900.230 1559.140 ;
        RECT 2452.790 1558.940 2453.110 1559.000 ;
        RECT 2899.910 1558.940 2900.230 1559.000 ;
      LAYER via ;
        RECT 1571.460 2380.720 1571.720 2380.980 ;
        RECT 2452.820 2380.720 2453.080 2380.980 ;
        RECT 2452.820 1558.940 2453.080 1559.200 ;
        RECT 2899.940 1558.940 2900.200 1559.200 ;
      LAYER met2 ;
        RECT 1571.460 2380.690 1571.720 2381.010 ;
        RECT 2452.820 2380.690 2453.080 2381.010 ;
        RECT 1571.520 2377.880 1571.660 2380.690 ;
        RECT 1571.500 2373.880 1571.780 2377.880 ;
        RECT 2452.880 1559.230 2453.020 2380.690 ;
        RECT 2452.820 1558.910 2453.080 1559.230 ;
        RECT 2899.940 1558.910 2900.200 1559.230 ;
        RECT 2900.000 1554.325 2900.140 1558.910 ;
        RECT 2899.930 1553.955 2900.210 1554.325 ;
      LAYER via2 ;
        RECT 2899.930 1554.000 2900.210 1554.280 ;
      LAYER met3 ;
        RECT 2899.905 1554.290 2900.235 1554.305 ;
        RECT 2917.600 1554.290 2924.800 1554.740 ;
        RECT 2899.905 1553.990 2924.800 1554.290 ;
        RECT 2899.905 1553.975 2900.235 1553.990 ;
        RECT 2917.600 1553.540 2924.800 1553.990 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 978.030 1318.760 978.350 1318.820 ;
        RECT 2904.050 1318.760 2904.370 1318.820 ;
        RECT 978.030 1318.620 2904.370 1318.760 ;
        RECT 978.030 1318.560 978.350 1318.620 ;
        RECT 2904.050 1318.560 2904.370 1318.620 ;
      LAYER via ;
        RECT 978.060 1318.560 978.320 1318.820 ;
        RECT 2904.080 1318.560 2904.340 1318.820 ;
      LAYER met2 ;
        RECT 2904.070 1789.235 2904.350 1789.605 ;
        RECT 978.100 1323.135 978.380 1327.135 ;
        RECT 978.120 1318.850 978.260 1323.135 ;
        RECT 2904.140 1318.850 2904.280 1789.235 ;
        RECT 978.060 1318.530 978.320 1318.850 ;
        RECT 2904.080 1318.530 2904.340 1318.850 ;
      LAYER via2 ;
        RECT 2904.070 1789.280 2904.350 1789.560 ;
      LAYER met3 ;
        RECT 2904.045 1789.570 2904.375 1789.585 ;
        RECT 2917.600 1789.570 2924.800 1790.020 ;
        RECT 2904.045 1789.270 2924.800 1789.570 ;
        RECT 2904.045 1789.255 2904.375 1789.270 ;
        RECT 2917.600 1788.820 2924.800 1789.270 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1290.830 1319.780 1291.150 1319.840 ;
        RECT 2903.130 1319.780 2903.450 1319.840 ;
        RECT 1290.830 1319.640 2903.450 1319.780 ;
        RECT 1290.830 1319.580 1291.150 1319.640 ;
        RECT 2903.130 1319.580 2903.450 1319.640 ;
      LAYER via ;
        RECT 1290.860 1319.580 1291.120 1319.840 ;
        RECT 2903.160 1319.580 2903.420 1319.840 ;
      LAYER met2 ;
        RECT 2903.150 2023.835 2903.430 2024.205 ;
        RECT 1290.900 1323.135 1291.180 1327.135 ;
        RECT 1290.920 1319.870 1291.060 1323.135 ;
        RECT 2903.220 1319.870 2903.360 2023.835 ;
        RECT 1290.860 1319.550 1291.120 1319.870 ;
        RECT 2903.160 1319.550 2903.420 1319.870 ;
      LAYER via2 ;
        RECT 2903.150 2023.880 2903.430 2024.160 ;
      LAYER met3 ;
        RECT 2903.125 2024.170 2903.455 2024.185 ;
        RECT 2917.600 2024.170 2924.800 2024.620 ;
        RECT 2903.125 2023.870 2924.800 2024.170 ;
        RECT 2903.125 2023.855 2903.455 2023.870 ;
        RECT 2917.600 2023.420 2924.800 2023.870 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 865.790 2384.320 866.110 2384.380 ;
        RECT 1756.810 2384.320 1757.130 2384.380 ;
        RECT 865.790 2384.180 1757.130 2384.320 ;
        RECT 865.790 2384.120 866.110 2384.180 ;
        RECT 1756.810 2384.120 1757.130 2384.180 ;
        RECT 1757.270 2262.940 1757.590 2263.000 ;
        RECT 2899.910 2262.940 2900.230 2263.000 ;
        RECT 1757.270 2262.800 2900.230 2262.940 ;
        RECT 1757.270 2262.740 1757.590 2262.800 ;
        RECT 2899.910 2262.740 2900.230 2262.800 ;
      LAYER via ;
        RECT 865.820 2384.120 866.080 2384.380 ;
        RECT 1756.840 2384.120 1757.100 2384.380 ;
        RECT 1757.300 2262.740 1757.560 2263.000 ;
        RECT 2899.940 2262.740 2900.200 2263.000 ;
      LAYER met2 ;
        RECT 865.820 2384.090 866.080 2384.410 ;
        RECT 1756.840 2384.090 1757.100 2384.410 ;
        RECT 865.880 2377.880 866.020 2384.090 ;
        RECT 865.860 2373.880 866.140 2377.880 ;
        RECT 1756.900 2308.330 1757.040 2384.090 ;
        RECT 1756.900 2308.190 1757.500 2308.330 ;
        RECT 1757.360 2263.030 1757.500 2308.190 ;
        RECT 1757.300 2262.710 1757.560 2263.030 ;
        RECT 2899.940 2262.710 2900.200 2263.030 ;
        RECT 2900.000 2258.805 2900.140 2262.710 ;
        RECT 2899.930 2258.435 2900.210 2258.805 ;
      LAYER via2 ;
        RECT 2899.930 2258.480 2900.210 2258.760 ;
      LAYER met3 ;
        RECT 2899.905 2258.770 2900.235 2258.785 ;
        RECT 2917.600 2258.770 2924.800 2259.220 ;
        RECT 2899.905 2258.470 2924.800 2258.770 ;
        RECT 2899.905 2258.455 2900.235 2258.470 ;
        RECT 2917.600 2258.020 2924.800 2258.470 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 633.030 45.800 633.350 45.860 ;
        RECT 1214.470 45.800 1214.790 45.860 ;
        RECT 633.030 45.660 1214.790 45.800 ;
        RECT 633.030 45.600 633.350 45.660 ;
        RECT 1214.470 45.600 1214.790 45.660 ;
      LAYER via ;
        RECT 633.060 45.600 633.320 45.860 ;
        RECT 1214.500 45.600 1214.760 45.860 ;
      LAYER met2 ;
        RECT 1215.460 1323.690 1215.740 1327.135 ;
        RECT 1214.560 1323.550 1215.740 1323.690 ;
        RECT 1214.560 45.890 1214.700 1323.550 ;
        RECT 1215.460 1323.135 1215.740 1323.550 ;
        RECT 633.060 45.570 633.320 45.890 ;
        RECT 1214.500 45.570 1214.760 45.890 ;
        RECT 633.120 2.400 633.260 45.570 ;
        RECT 632.910 -4.800 633.470 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1772.910 1456.120 1773.230 1456.180 ;
        RECT 2415.070 1456.120 2415.390 1456.180 ;
        RECT 1772.910 1455.980 2415.390 1456.120 ;
        RECT 1772.910 1455.920 1773.230 1455.980 ;
        RECT 2415.070 1455.920 2415.390 1455.980 ;
        RECT 2415.070 72.660 2415.390 72.720 ;
        RECT 2418.290 72.660 2418.610 72.720 ;
        RECT 2415.070 72.520 2418.610 72.660 ;
        RECT 2415.070 72.460 2415.390 72.520 ;
        RECT 2418.290 72.460 2418.610 72.520 ;
        RECT 2417.370 47.980 2417.690 48.240 ;
        RECT 2417.460 47.560 2417.600 47.980 ;
        RECT 2417.370 47.300 2417.690 47.560 ;
      LAYER via ;
        RECT 1772.940 1455.920 1773.200 1456.180 ;
        RECT 2415.100 1455.920 2415.360 1456.180 ;
        RECT 2415.100 72.460 2415.360 72.720 ;
        RECT 2418.320 72.460 2418.580 72.720 ;
        RECT 2417.400 47.980 2417.660 48.240 ;
        RECT 2417.400 47.300 2417.660 47.560 ;
      LAYER met2 ;
        RECT 1772.930 1459.435 1773.210 1459.805 ;
        RECT 1773.000 1456.210 1773.140 1459.435 ;
        RECT 1772.940 1455.890 1773.200 1456.210 ;
        RECT 2415.100 1455.890 2415.360 1456.210 ;
        RECT 2415.160 72.750 2415.300 1455.890 ;
        RECT 2415.100 72.430 2415.360 72.750 ;
        RECT 2418.320 72.430 2418.580 72.750 ;
        RECT 2418.380 48.805 2418.520 72.430 ;
        RECT 2417.390 48.435 2417.670 48.805 ;
        RECT 2418.310 48.435 2418.590 48.805 ;
        RECT 2417.460 48.270 2417.600 48.435 ;
        RECT 2417.400 47.950 2417.660 48.270 ;
        RECT 2417.400 47.270 2417.660 47.590 ;
        RECT 2417.460 2.400 2417.600 47.270 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
      LAYER via2 ;
        RECT 1772.930 1459.480 1773.210 1459.760 ;
        RECT 2417.390 48.480 2417.670 48.760 ;
        RECT 2418.310 48.480 2418.590 48.760 ;
      LAYER met3 ;
        RECT 1755.835 1459.770 1759.835 1459.775 ;
        RECT 1772.905 1459.770 1773.235 1459.785 ;
        RECT 1755.835 1459.470 1773.235 1459.770 ;
        RECT 1755.835 1459.175 1759.835 1459.470 ;
        RECT 1772.905 1459.455 1773.235 1459.470 ;
        RECT 2417.365 48.770 2417.695 48.785 ;
        RECT 2418.285 48.770 2418.615 48.785 ;
        RECT 2417.365 48.470 2418.615 48.770 ;
        RECT 2417.365 48.455 2417.695 48.470 ;
        RECT 2418.285 48.455 2418.615 48.470 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1738.410 37.980 1738.730 38.040 ;
        RECT 2434.850 37.980 2435.170 38.040 ;
        RECT 1738.410 37.840 2435.170 37.980 ;
        RECT 1738.410 37.780 1738.730 37.840 ;
        RECT 2434.850 37.780 2435.170 37.840 ;
      LAYER via ;
        RECT 1738.440 37.780 1738.700 38.040 ;
        RECT 2434.880 37.780 2435.140 38.040 ;
      LAYER met2 ;
        RECT 1736.180 1323.690 1736.460 1327.135 ;
        RECT 1736.180 1323.550 1738.640 1323.690 ;
        RECT 1736.180 1323.135 1736.460 1323.550 ;
        RECT 1738.500 38.070 1738.640 1323.550 ;
        RECT 1738.440 37.750 1738.700 38.070 ;
        RECT 2434.880 37.750 2435.140 38.070 ;
        RECT 2434.940 2.400 2435.080 37.750 ;
        RECT 2434.730 -4.800 2435.290 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2452.865 2.805 2453.035 20.315 ;
      LAYER mcon ;
        RECT 2452.865 20.145 2453.035 20.315 ;
      LAYER met1 ;
        RECT 1057.150 2381.260 1057.470 2381.320 ;
        RECT 2449.570 2381.260 2449.890 2381.320 ;
        RECT 1057.150 2381.120 2449.890 2381.260 ;
        RECT 1057.150 2381.060 1057.470 2381.120 ;
        RECT 2449.570 2381.060 2449.890 2381.120 ;
        RECT 2449.570 20.300 2449.890 20.360 ;
        RECT 2452.805 20.300 2453.095 20.345 ;
        RECT 2449.570 20.160 2453.095 20.300 ;
        RECT 2449.570 20.100 2449.890 20.160 ;
        RECT 2452.805 20.115 2453.095 20.160 ;
        RECT 2452.790 2.960 2453.110 3.020 ;
        RECT 2452.595 2.820 2453.110 2.960 ;
        RECT 2452.790 2.760 2453.110 2.820 ;
      LAYER via ;
        RECT 1057.180 2381.060 1057.440 2381.320 ;
        RECT 2449.600 2381.060 2449.860 2381.320 ;
        RECT 2449.600 20.100 2449.860 20.360 ;
        RECT 2452.820 2.760 2453.080 3.020 ;
      LAYER met2 ;
        RECT 1057.180 2381.030 1057.440 2381.350 ;
        RECT 2449.600 2381.030 2449.860 2381.350 ;
        RECT 1057.240 2377.880 1057.380 2381.030 ;
        RECT 1057.220 2373.880 1057.500 2377.880 ;
        RECT 2449.660 20.390 2449.800 2381.030 ;
        RECT 2449.600 20.070 2449.860 20.390 ;
        RECT 2452.820 2.730 2453.080 3.050 ;
        RECT 2452.880 2.400 2453.020 2.730 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2470.345 2173.705 2470.515 2221.815 ;
        RECT 2470.345 2077.145 2470.515 2125.255 ;
        RECT 2470.345 1883.685 2470.515 1931.795 ;
        RECT 2470.345 1787.125 2470.515 1835.235 ;
        RECT 2470.345 1690.565 2470.515 1738.675 ;
        RECT 2470.345 1594.005 2470.515 1642.115 ;
        RECT 2470.345 1497.445 2470.515 1545.555 ;
        RECT 2470.345 1400.885 2470.515 1448.995 ;
        RECT 2470.345 1304.325 2470.515 1352.435 ;
        RECT 2470.345 1207.425 2470.515 1255.875 ;
        RECT 2470.345 628.065 2470.515 675.835 ;
        RECT 2470.345 531.505 2470.515 579.615 ;
        RECT 2470.345 434.945 2470.515 483.055 ;
        RECT 2470.345 338.045 2470.515 386.155 ;
        RECT 2470.345 241.485 2470.515 289.595 ;
        RECT 2470.345 144.925 2470.515 193.035 ;
        RECT 2470.345 48.365 2470.515 96.475 ;
        RECT 2470.805 2.805 2470.975 16.915 ;
      LAYER mcon ;
        RECT 2470.345 2221.645 2470.515 2221.815 ;
        RECT 2470.345 2125.085 2470.515 2125.255 ;
        RECT 2470.345 1931.625 2470.515 1931.795 ;
        RECT 2470.345 1835.065 2470.515 1835.235 ;
        RECT 2470.345 1738.505 2470.515 1738.675 ;
        RECT 2470.345 1641.945 2470.515 1642.115 ;
        RECT 2470.345 1545.385 2470.515 1545.555 ;
        RECT 2470.345 1448.825 2470.515 1448.995 ;
        RECT 2470.345 1352.265 2470.515 1352.435 ;
        RECT 2470.345 1255.705 2470.515 1255.875 ;
        RECT 2470.345 675.665 2470.515 675.835 ;
        RECT 2470.345 579.445 2470.515 579.615 ;
        RECT 2470.345 482.885 2470.515 483.055 ;
        RECT 2470.345 385.985 2470.515 386.155 ;
        RECT 2470.345 289.425 2470.515 289.595 ;
        RECT 2470.345 192.865 2470.515 193.035 ;
        RECT 2470.345 96.305 2470.515 96.475 ;
        RECT 2470.805 16.745 2470.975 16.915 ;
      LAYER met1 ;
        RECT 1623.870 2382.620 1624.190 2382.680 ;
        RECT 2465.210 2382.620 2465.530 2382.680 ;
        RECT 1623.870 2382.480 2465.530 2382.620 ;
        RECT 1623.870 2382.420 1624.190 2382.480 ;
        RECT 2465.210 2382.420 2465.530 2382.480 ;
        RECT 2469.350 2318.360 2469.670 2318.420 ;
        RECT 2470.270 2318.360 2470.590 2318.420 ;
        RECT 2469.350 2318.220 2470.590 2318.360 ;
        RECT 2469.350 2318.160 2469.670 2318.220 ;
        RECT 2470.270 2318.160 2470.590 2318.220 ;
        RECT 2470.270 2221.800 2470.590 2221.860 ;
        RECT 2470.075 2221.660 2470.590 2221.800 ;
        RECT 2470.270 2221.600 2470.590 2221.660 ;
        RECT 2470.270 2173.860 2470.590 2173.920 ;
        RECT 2470.075 2173.720 2470.590 2173.860 ;
        RECT 2470.270 2173.660 2470.590 2173.720 ;
        RECT 2470.270 2125.240 2470.590 2125.300 ;
        RECT 2470.075 2125.100 2470.590 2125.240 ;
        RECT 2470.270 2125.040 2470.590 2125.100 ;
        RECT 2470.270 2077.300 2470.590 2077.360 ;
        RECT 2470.075 2077.160 2470.590 2077.300 ;
        RECT 2470.270 2077.100 2470.590 2077.160 ;
        RECT 2470.270 1931.780 2470.590 1931.840 ;
        RECT 2470.075 1931.640 2470.590 1931.780 ;
        RECT 2470.270 1931.580 2470.590 1931.640 ;
        RECT 2470.270 1883.840 2470.590 1883.900 ;
        RECT 2470.075 1883.700 2470.590 1883.840 ;
        RECT 2470.270 1883.640 2470.590 1883.700 ;
        RECT 2470.270 1835.220 2470.590 1835.280 ;
        RECT 2470.075 1835.080 2470.590 1835.220 ;
        RECT 2470.270 1835.020 2470.590 1835.080 ;
        RECT 2470.270 1787.280 2470.590 1787.340 ;
        RECT 2470.075 1787.140 2470.590 1787.280 ;
        RECT 2470.270 1787.080 2470.590 1787.140 ;
        RECT 2470.270 1738.660 2470.590 1738.720 ;
        RECT 2470.075 1738.520 2470.590 1738.660 ;
        RECT 2470.270 1738.460 2470.590 1738.520 ;
        RECT 2470.270 1690.720 2470.590 1690.780 ;
        RECT 2470.075 1690.580 2470.590 1690.720 ;
        RECT 2470.270 1690.520 2470.590 1690.580 ;
        RECT 2470.270 1642.100 2470.590 1642.160 ;
        RECT 2470.075 1641.960 2470.590 1642.100 ;
        RECT 2470.270 1641.900 2470.590 1641.960 ;
        RECT 2470.270 1594.160 2470.590 1594.220 ;
        RECT 2470.075 1594.020 2470.590 1594.160 ;
        RECT 2470.270 1593.960 2470.590 1594.020 ;
        RECT 2470.270 1545.540 2470.590 1545.600 ;
        RECT 2470.075 1545.400 2470.590 1545.540 ;
        RECT 2470.270 1545.340 2470.590 1545.400 ;
        RECT 2470.270 1497.600 2470.590 1497.660 ;
        RECT 2470.075 1497.460 2470.590 1497.600 ;
        RECT 2470.270 1497.400 2470.590 1497.460 ;
        RECT 2470.270 1448.980 2470.590 1449.040 ;
        RECT 2470.075 1448.840 2470.590 1448.980 ;
        RECT 2470.270 1448.780 2470.590 1448.840 ;
        RECT 2470.270 1401.040 2470.590 1401.100 ;
        RECT 2470.075 1400.900 2470.590 1401.040 ;
        RECT 2470.270 1400.840 2470.590 1400.900 ;
        RECT 2470.270 1352.420 2470.590 1352.480 ;
        RECT 2470.075 1352.280 2470.590 1352.420 ;
        RECT 2470.270 1352.220 2470.590 1352.280 ;
        RECT 2470.270 1304.480 2470.590 1304.540 ;
        RECT 2470.075 1304.340 2470.590 1304.480 ;
        RECT 2470.270 1304.280 2470.590 1304.340 ;
        RECT 2470.270 1255.860 2470.590 1255.920 ;
        RECT 2470.075 1255.720 2470.590 1255.860 ;
        RECT 2470.270 1255.660 2470.590 1255.720 ;
        RECT 2470.270 1207.580 2470.590 1207.640 ;
        RECT 2470.075 1207.440 2470.590 1207.580 ;
        RECT 2470.270 1207.380 2470.590 1207.440 ;
        RECT 2470.270 1111.020 2470.590 1111.080 ;
        RECT 2471.190 1111.020 2471.510 1111.080 ;
        RECT 2470.270 1110.880 2471.510 1111.020 ;
        RECT 2470.270 1110.820 2470.590 1110.880 ;
        RECT 2471.190 1110.820 2471.510 1110.880 ;
        RECT 2470.270 1014.460 2470.590 1014.520 ;
        RECT 2471.190 1014.460 2471.510 1014.520 ;
        RECT 2470.270 1014.320 2471.510 1014.460 ;
        RECT 2470.270 1014.260 2470.590 1014.320 ;
        RECT 2471.190 1014.260 2471.510 1014.320 ;
        RECT 2470.270 917.900 2470.590 917.960 ;
        RECT 2471.190 917.900 2471.510 917.960 ;
        RECT 2470.270 917.760 2471.510 917.900 ;
        RECT 2470.270 917.700 2470.590 917.760 ;
        RECT 2471.190 917.700 2471.510 917.760 ;
        RECT 2470.270 772.720 2470.590 772.780 ;
        RECT 2471.190 772.720 2471.510 772.780 ;
        RECT 2470.270 772.580 2471.510 772.720 ;
        RECT 2470.270 772.520 2470.590 772.580 ;
        RECT 2471.190 772.520 2471.510 772.580 ;
        RECT 2470.270 675.820 2470.590 675.880 ;
        RECT 2470.075 675.680 2470.590 675.820 ;
        RECT 2470.270 675.620 2470.590 675.680 ;
        RECT 2470.270 628.220 2470.590 628.280 ;
        RECT 2470.075 628.080 2470.590 628.220 ;
        RECT 2470.270 628.020 2470.590 628.080 ;
        RECT 2470.270 579.600 2470.590 579.660 ;
        RECT 2470.075 579.460 2470.590 579.600 ;
        RECT 2470.270 579.400 2470.590 579.460 ;
        RECT 2470.270 531.660 2470.590 531.720 ;
        RECT 2470.075 531.520 2470.590 531.660 ;
        RECT 2470.270 531.460 2470.590 531.520 ;
        RECT 2470.270 483.040 2470.590 483.100 ;
        RECT 2470.075 482.900 2470.590 483.040 ;
        RECT 2470.270 482.840 2470.590 482.900 ;
        RECT 2470.270 435.100 2470.590 435.160 ;
        RECT 2470.075 434.960 2470.590 435.100 ;
        RECT 2470.270 434.900 2470.590 434.960 ;
        RECT 2470.270 386.140 2470.590 386.200 ;
        RECT 2470.075 386.000 2470.590 386.140 ;
        RECT 2470.270 385.940 2470.590 386.000 ;
        RECT 2470.270 338.200 2470.590 338.260 ;
        RECT 2470.075 338.060 2470.590 338.200 ;
        RECT 2470.270 338.000 2470.590 338.060 ;
        RECT 2470.270 289.580 2470.590 289.640 ;
        RECT 2470.075 289.440 2470.590 289.580 ;
        RECT 2470.270 289.380 2470.590 289.440 ;
        RECT 2470.270 241.640 2470.590 241.700 ;
        RECT 2470.075 241.500 2470.590 241.640 ;
        RECT 2470.270 241.440 2470.590 241.500 ;
        RECT 2470.270 193.020 2470.590 193.080 ;
        RECT 2470.075 192.880 2470.590 193.020 ;
        RECT 2470.270 192.820 2470.590 192.880 ;
        RECT 2470.270 145.080 2470.590 145.140 ;
        RECT 2470.075 144.940 2470.590 145.080 ;
        RECT 2470.270 144.880 2470.590 144.940 ;
        RECT 2470.270 96.460 2470.590 96.520 ;
        RECT 2470.075 96.320 2470.590 96.460 ;
        RECT 2470.270 96.260 2470.590 96.320 ;
        RECT 2470.270 48.520 2470.590 48.580 ;
        RECT 2470.075 48.380 2470.590 48.520 ;
        RECT 2470.270 48.320 2470.590 48.380 ;
        RECT 2470.270 16.900 2470.590 16.960 ;
        RECT 2470.745 16.900 2471.035 16.945 ;
        RECT 2470.270 16.760 2471.035 16.900 ;
        RECT 2470.270 16.700 2470.590 16.760 ;
        RECT 2470.745 16.715 2471.035 16.760 ;
        RECT 2470.730 2.960 2471.050 3.020 ;
        RECT 2470.535 2.820 2471.050 2.960 ;
        RECT 2470.730 2.760 2471.050 2.820 ;
      LAYER via ;
        RECT 1623.900 2382.420 1624.160 2382.680 ;
        RECT 2465.240 2382.420 2465.500 2382.680 ;
        RECT 2469.380 2318.160 2469.640 2318.420 ;
        RECT 2470.300 2318.160 2470.560 2318.420 ;
        RECT 2470.300 2221.600 2470.560 2221.860 ;
        RECT 2470.300 2173.660 2470.560 2173.920 ;
        RECT 2470.300 2125.040 2470.560 2125.300 ;
        RECT 2470.300 2077.100 2470.560 2077.360 ;
        RECT 2470.300 1931.580 2470.560 1931.840 ;
        RECT 2470.300 1883.640 2470.560 1883.900 ;
        RECT 2470.300 1835.020 2470.560 1835.280 ;
        RECT 2470.300 1787.080 2470.560 1787.340 ;
        RECT 2470.300 1738.460 2470.560 1738.720 ;
        RECT 2470.300 1690.520 2470.560 1690.780 ;
        RECT 2470.300 1641.900 2470.560 1642.160 ;
        RECT 2470.300 1593.960 2470.560 1594.220 ;
        RECT 2470.300 1545.340 2470.560 1545.600 ;
        RECT 2470.300 1497.400 2470.560 1497.660 ;
        RECT 2470.300 1448.780 2470.560 1449.040 ;
        RECT 2470.300 1400.840 2470.560 1401.100 ;
        RECT 2470.300 1352.220 2470.560 1352.480 ;
        RECT 2470.300 1304.280 2470.560 1304.540 ;
        RECT 2470.300 1255.660 2470.560 1255.920 ;
        RECT 2470.300 1207.380 2470.560 1207.640 ;
        RECT 2470.300 1110.820 2470.560 1111.080 ;
        RECT 2471.220 1110.820 2471.480 1111.080 ;
        RECT 2470.300 1014.260 2470.560 1014.520 ;
        RECT 2471.220 1014.260 2471.480 1014.520 ;
        RECT 2470.300 917.700 2470.560 917.960 ;
        RECT 2471.220 917.700 2471.480 917.960 ;
        RECT 2470.300 772.520 2470.560 772.780 ;
        RECT 2471.220 772.520 2471.480 772.780 ;
        RECT 2470.300 675.620 2470.560 675.880 ;
        RECT 2470.300 628.020 2470.560 628.280 ;
        RECT 2470.300 579.400 2470.560 579.660 ;
        RECT 2470.300 531.460 2470.560 531.720 ;
        RECT 2470.300 482.840 2470.560 483.100 ;
        RECT 2470.300 434.900 2470.560 435.160 ;
        RECT 2470.300 385.940 2470.560 386.200 ;
        RECT 2470.300 338.000 2470.560 338.260 ;
        RECT 2470.300 289.380 2470.560 289.640 ;
        RECT 2470.300 241.440 2470.560 241.700 ;
        RECT 2470.300 192.820 2470.560 193.080 ;
        RECT 2470.300 144.880 2470.560 145.140 ;
        RECT 2470.300 96.260 2470.560 96.520 ;
        RECT 2470.300 48.320 2470.560 48.580 ;
        RECT 2470.300 16.700 2470.560 16.960 ;
        RECT 2470.760 2.760 2471.020 3.020 ;
      LAYER met2 ;
        RECT 1623.900 2382.390 1624.160 2382.710 ;
        RECT 2465.240 2382.390 2465.500 2382.710 ;
        RECT 1623.960 2377.880 1624.100 2382.390 ;
        RECT 1623.940 2373.880 1624.220 2377.880 ;
        RECT 2465.300 2366.925 2465.440 2382.390 ;
        RECT 2465.230 2366.555 2465.510 2366.925 ;
        RECT 2470.290 2366.555 2470.570 2366.925 ;
        RECT 2470.360 2318.450 2470.500 2366.555 ;
        RECT 2469.380 2318.130 2469.640 2318.450 ;
        RECT 2470.300 2318.130 2470.560 2318.450 ;
        RECT 2469.440 2270.365 2469.580 2318.130 ;
        RECT 2469.370 2269.995 2469.650 2270.365 ;
        RECT 2470.290 2269.995 2470.570 2270.365 ;
        RECT 2470.360 2221.890 2470.500 2269.995 ;
        RECT 2470.300 2221.570 2470.560 2221.890 ;
        RECT 2470.300 2173.630 2470.560 2173.950 ;
        RECT 2470.360 2125.330 2470.500 2173.630 ;
        RECT 2470.300 2125.010 2470.560 2125.330 ;
        RECT 2470.300 2077.070 2470.560 2077.390 ;
        RECT 2470.360 1931.870 2470.500 2077.070 ;
        RECT 2470.300 1931.550 2470.560 1931.870 ;
        RECT 2470.300 1883.610 2470.560 1883.930 ;
        RECT 2470.360 1835.310 2470.500 1883.610 ;
        RECT 2470.300 1834.990 2470.560 1835.310 ;
        RECT 2470.300 1787.050 2470.560 1787.370 ;
        RECT 2470.360 1738.750 2470.500 1787.050 ;
        RECT 2470.300 1738.430 2470.560 1738.750 ;
        RECT 2470.300 1690.490 2470.560 1690.810 ;
        RECT 2470.360 1642.190 2470.500 1690.490 ;
        RECT 2470.300 1641.870 2470.560 1642.190 ;
        RECT 2470.300 1593.930 2470.560 1594.250 ;
        RECT 2470.360 1545.630 2470.500 1593.930 ;
        RECT 2470.300 1545.310 2470.560 1545.630 ;
        RECT 2470.300 1497.370 2470.560 1497.690 ;
        RECT 2470.360 1449.070 2470.500 1497.370 ;
        RECT 2470.300 1448.750 2470.560 1449.070 ;
        RECT 2470.300 1400.810 2470.560 1401.130 ;
        RECT 2470.360 1352.510 2470.500 1400.810 ;
        RECT 2470.300 1352.190 2470.560 1352.510 ;
        RECT 2470.300 1304.250 2470.560 1304.570 ;
        RECT 2470.360 1255.950 2470.500 1304.250 ;
        RECT 2470.300 1255.630 2470.560 1255.950 ;
        RECT 2470.300 1207.350 2470.560 1207.670 ;
        RECT 2470.360 1159.245 2470.500 1207.350 ;
        RECT 2470.290 1158.875 2470.570 1159.245 ;
        RECT 2471.210 1158.875 2471.490 1159.245 ;
        RECT 2471.280 1111.110 2471.420 1158.875 ;
        RECT 2470.300 1110.790 2470.560 1111.110 ;
        RECT 2471.220 1110.790 2471.480 1111.110 ;
        RECT 2470.360 1062.685 2470.500 1110.790 ;
        RECT 2470.290 1062.315 2470.570 1062.685 ;
        RECT 2471.210 1062.315 2471.490 1062.685 ;
        RECT 2471.280 1014.550 2471.420 1062.315 ;
        RECT 2470.300 1014.230 2470.560 1014.550 ;
        RECT 2471.220 1014.230 2471.480 1014.550 ;
        RECT 2470.360 966.125 2470.500 1014.230 ;
        RECT 2470.290 965.755 2470.570 966.125 ;
        RECT 2471.210 965.755 2471.490 966.125 ;
        RECT 2471.280 917.990 2471.420 965.755 ;
        RECT 2470.300 917.670 2470.560 917.990 ;
        RECT 2471.220 917.670 2471.480 917.990 ;
        RECT 2470.360 869.565 2470.500 917.670 ;
        RECT 2470.290 869.195 2470.570 869.565 ;
        RECT 2471.210 869.195 2471.490 869.565 ;
        RECT 2471.280 821.285 2471.420 869.195 ;
        RECT 2470.290 820.915 2470.570 821.285 ;
        RECT 2471.210 820.915 2471.490 821.285 ;
        RECT 2470.360 772.810 2470.500 820.915 ;
        RECT 2470.300 772.490 2470.560 772.810 ;
        RECT 2471.220 772.490 2471.480 772.810 ;
        RECT 2471.280 724.725 2471.420 772.490 ;
        RECT 2470.290 724.355 2470.570 724.725 ;
        RECT 2471.210 724.355 2471.490 724.725 ;
        RECT 2470.360 675.910 2470.500 724.355 ;
        RECT 2470.300 675.590 2470.560 675.910 ;
        RECT 2470.300 627.990 2470.560 628.310 ;
        RECT 2470.360 579.690 2470.500 627.990 ;
        RECT 2470.300 579.370 2470.560 579.690 ;
        RECT 2470.300 531.430 2470.560 531.750 ;
        RECT 2470.360 483.130 2470.500 531.430 ;
        RECT 2470.300 482.810 2470.560 483.130 ;
        RECT 2470.300 434.870 2470.560 435.190 ;
        RECT 2470.360 386.230 2470.500 434.870 ;
        RECT 2470.300 385.910 2470.560 386.230 ;
        RECT 2470.300 337.970 2470.560 338.290 ;
        RECT 2470.360 289.670 2470.500 337.970 ;
        RECT 2470.300 289.350 2470.560 289.670 ;
        RECT 2470.300 241.410 2470.560 241.730 ;
        RECT 2470.360 193.110 2470.500 241.410 ;
        RECT 2470.300 192.790 2470.560 193.110 ;
        RECT 2470.300 144.850 2470.560 145.170 ;
        RECT 2470.360 96.550 2470.500 144.850 ;
        RECT 2470.300 96.230 2470.560 96.550 ;
        RECT 2470.300 48.290 2470.560 48.610 ;
        RECT 2470.360 16.990 2470.500 48.290 ;
        RECT 2470.300 16.670 2470.560 16.990 ;
        RECT 2470.760 2.730 2471.020 3.050 ;
        RECT 2470.820 2.400 2470.960 2.730 ;
        RECT 2470.610 -4.800 2471.170 2.400 ;
      LAYER via2 ;
        RECT 2465.230 2366.600 2465.510 2366.880 ;
        RECT 2470.290 2366.600 2470.570 2366.880 ;
        RECT 2469.370 2270.040 2469.650 2270.320 ;
        RECT 2470.290 2270.040 2470.570 2270.320 ;
        RECT 2470.290 1158.920 2470.570 1159.200 ;
        RECT 2471.210 1158.920 2471.490 1159.200 ;
        RECT 2470.290 1062.360 2470.570 1062.640 ;
        RECT 2471.210 1062.360 2471.490 1062.640 ;
        RECT 2470.290 965.800 2470.570 966.080 ;
        RECT 2471.210 965.800 2471.490 966.080 ;
        RECT 2470.290 869.240 2470.570 869.520 ;
        RECT 2471.210 869.240 2471.490 869.520 ;
        RECT 2470.290 820.960 2470.570 821.240 ;
        RECT 2471.210 820.960 2471.490 821.240 ;
        RECT 2470.290 724.400 2470.570 724.680 ;
        RECT 2471.210 724.400 2471.490 724.680 ;
      LAYER met3 ;
        RECT 2465.205 2366.890 2465.535 2366.905 ;
        RECT 2470.265 2366.890 2470.595 2366.905 ;
        RECT 2465.205 2366.590 2470.595 2366.890 ;
        RECT 2465.205 2366.575 2465.535 2366.590 ;
        RECT 2470.265 2366.575 2470.595 2366.590 ;
        RECT 2469.345 2270.330 2469.675 2270.345 ;
        RECT 2470.265 2270.330 2470.595 2270.345 ;
        RECT 2469.345 2270.030 2470.595 2270.330 ;
        RECT 2469.345 2270.015 2469.675 2270.030 ;
        RECT 2470.265 2270.015 2470.595 2270.030 ;
        RECT 2470.265 1159.210 2470.595 1159.225 ;
        RECT 2471.185 1159.210 2471.515 1159.225 ;
        RECT 2470.265 1158.910 2471.515 1159.210 ;
        RECT 2470.265 1158.895 2470.595 1158.910 ;
        RECT 2471.185 1158.895 2471.515 1158.910 ;
        RECT 2470.265 1062.650 2470.595 1062.665 ;
        RECT 2471.185 1062.650 2471.515 1062.665 ;
        RECT 2470.265 1062.350 2471.515 1062.650 ;
        RECT 2470.265 1062.335 2470.595 1062.350 ;
        RECT 2471.185 1062.335 2471.515 1062.350 ;
        RECT 2470.265 966.090 2470.595 966.105 ;
        RECT 2471.185 966.090 2471.515 966.105 ;
        RECT 2470.265 965.790 2471.515 966.090 ;
        RECT 2470.265 965.775 2470.595 965.790 ;
        RECT 2471.185 965.775 2471.515 965.790 ;
        RECT 2470.265 869.530 2470.595 869.545 ;
        RECT 2471.185 869.530 2471.515 869.545 ;
        RECT 2470.265 869.230 2471.515 869.530 ;
        RECT 2470.265 869.215 2470.595 869.230 ;
        RECT 2471.185 869.215 2471.515 869.230 ;
        RECT 2470.265 821.250 2470.595 821.265 ;
        RECT 2471.185 821.250 2471.515 821.265 ;
        RECT 2470.265 820.950 2471.515 821.250 ;
        RECT 2470.265 820.935 2470.595 820.950 ;
        RECT 2471.185 820.935 2471.515 820.950 ;
        RECT 2470.265 724.690 2470.595 724.705 ;
        RECT 2471.185 724.690 2471.515 724.705 ;
        RECT 2470.265 724.390 2471.515 724.690 ;
        RECT 2470.265 724.375 2470.595 724.390 ;
        RECT 2471.185 724.375 2471.515 724.390 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1409.510 2387.720 1409.830 2387.780 ;
        RECT 1441.710 2387.720 1442.030 2387.780 ;
        RECT 1409.510 2387.580 1442.030 2387.720 ;
        RECT 1409.510 2387.520 1409.830 2387.580 ;
        RECT 1441.710 2387.520 1442.030 2387.580 ;
        RECT 1441.710 2376.840 1442.030 2376.900 ;
        RECT 2484.070 2376.840 2484.390 2376.900 ;
        RECT 1441.710 2376.700 2484.390 2376.840 ;
        RECT 1441.710 2376.640 1442.030 2376.700 ;
        RECT 2484.070 2376.640 2484.390 2376.700 ;
      LAYER via ;
        RECT 1409.540 2387.520 1409.800 2387.780 ;
        RECT 1441.740 2387.520 1442.000 2387.780 ;
        RECT 1441.740 2376.640 1442.000 2376.900 ;
        RECT 2484.100 2376.640 2484.360 2376.900 ;
      LAYER met2 ;
        RECT 1409.540 2387.490 1409.800 2387.810 ;
        RECT 1441.740 2387.490 1442.000 2387.810 ;
        RECT 1409.600 2377.880 1409.740 2387.490 ;
        RECT 1409.580 2373.880 1409.860 2377.880 ;
        RECT 1441.800 2376.930 1441.940 2387.490 ;
        RECT 1441.740 2376.610 1442.000 2376.930 ;
        RECT 2484.100 2376.610 2484.360 2376.930 ;
        RECT 2484.160 24.210 2484.300 2376.610 ;
        RECT 2484.160 24.070 2488.900 24.210 ;
        RECT 2488.760 2.400 2488.900 24.070 ;
        RECT 2488.550 -4.800 2489.110 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1524.510 46.820 1524.830 46.880 ;
        RECT 2506.150 46.820 2506.470 46.880 ;
        RECT 1524.510 46.680 2506.470 46.820 ;
        RECT 1524.510 46.620 1524.830 46.680 ;
        RECT 2506.150 46.620 2506.470 46.680 ;
      LAYER via ;
        RECT 1524.540 46.620 1524.800 46.880 ;
        RECT 2506.180 46.620 2506.440 46.880 ;
      LAYER met2 ;
        RECT 1522.740 1323.690 1523.020 1327.135 ;
        RECT 1522.740 1323.550 1524.740 1323.690 ;
        RECT 1522.740 1323.135 1523.020 1323.550 ;
        RECT 1524.600 46.910 1524.740 1323.550 ;
        RECT 1524.540 46.590 1524.800 46.910 ;
        RECT 2506.180 46.590 2506.440 46.910 ;
        RECT 2506.240 2.400 2506.380 46.590 ;
        RECT 2506.030 -4.800 2506.590 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1283.470 13.500 1283.790 13.560 ;
        RECT 1331.310 13.500 1331.630 13.560 ;
        RECT 1283.470 13.360 1331.630 13.500 ;
        RECT 1283.470 13.300 1283.790 13.360 ;
        RECT 1331.310 13.300 1331.630 13.360 ;
      LAYER via ;
        RECT 1283.500 13.300 1283.760 13.560 ;
        RECT 1331.340 13.300 1331.600 13.560 ;
      LAYER met2 ;
        RECT 2524.110 15.115 2524.390 15.485 ;
        RECT 1331.330 13.755 1331.610 14.125 ;
        RECT 1331.400 13.590 1331.540 13.755 ;
        RECT 1283.500 13.445 1283.760 13.590 ;
        RECT 1283.490 13.075 1283.770 13.445 ;
        RECT 1331.340 13.270 1331.600 13.590 ;
        RECT 2524.180 2.400 2524.320 15.115 ;
        RECT 2523.970 -4.800 2524.530 2.400 ;
      LAYER via2 ;
        RECT 2524.110 15.160 2524.390 15.440 ;
        RECT 1331.330 13.800 1331.610 14.080 ;
        RECT 1283.490 13.120 1283.770 13.400 ;
      LAYER met3 ;
        RECT 694.870 1746.730 695.250 1746.740 ;
        RECT 715.810 1746.730 719.810 1746.735 ;
        RECT 694.870 1746.430 719.810 1746.730 ;
        RECT 694.870 1746.420 695.250 1746.430 ;
        RECT 715.810 1746.135 719.810 1746.430 ;
        RECT 1714.230 20.890 1714.610 20.900 ;
        RECT 1804.390 20.890 1804.770 20.900 ;
        RECT 1714.230 20.590 1804.770 20.890 ;
        RECT 1714.230 20.580 1714.610 20.590 ;
        RECT 1804.390 20.580 1804.770 20.590 ;
        RECT 1852.230 15.450 1852.610 15.460 ;
        RECT 2110.750 15.450 2111.130 15.460 ;
        RECT 1852.230 15.150 2111.130 15.450 ;
        RECT 1852.230 15.140 1852.610 15.150 ;
        RECT 2110.750 15.140 2111.130 15.150 ;
        RECT 2200.910 15.450 2201.290 15.460 ;
        RECT 2248.750 15.450 2249.130 15.460 ;
        RECT 2200.910 15.150 2249.130 15.450 ;
        RECT 2200.910 15.140 2201.290 15.150 ;
        RECT 2248.750 15.140 2249.130 15.150 ;
        RECT 2305.790 15.450 2306.170 15.460 ;
        RECT 2498.070 15.450 2498.450 15.460 ;
        RECT 2305.790 15.150 2498.450 15.450 ;
        RECT 2305.790 15.140 2306.170 15.150 ;
        RECT 2498.070 15.140 2498.450 15.150 ;
        RECT 2509.110 15.450 2509.490 15.460 ;
        RECT 2524.085 15.450 2524.415 15.465 ;
        RECT 2509.110 15.150 2524.415 15.450 ;
        RECT 2509.110 15.140 2509.490 15.150 ;
        RECT 2524.085 15.135 2524.415 15.150 ;
        RECT 741.790 14.090 742.170 14.100 ;
        RECT 785.950 14.090 786.330 14.100 ;
        RECT 741.790 13.790 786.330 14.090 ;
        RECT 741.790 13.780 742.170 13.790 ;
        RECT 785.950 13.780 786.330 13.790 ;
        RECT 1331.305 14.090 1331.635 14.105 ;
        RECT 1355.430 14.090 1355.810 14.100 ;
        RECT 1331.305 13.790 1355.810 14.090 ;
        RECT 1331.305 13.775 1331.635 13.790 ;
        RECT 1355.430 13.780 1355.810 13.790 ;
        RECT 1234.910 13.410 1235.290 13.420 ;
        RECT 1283.465 13.410 1283.795 13.425 ;
        RECT 1234.910 13.110 1283.795 13.410 ;
        RECT 1234.910 13.100 1235.290 13.110 ;
        RECT 1283.465 13.095 1283.795 13.110 ;
        RECT 1055.510 12.050 1055.890 12.060 ;
        RECT 1103.350 12.050 1103.730 12.060 ;
        RECT 1055.510 11.750 1103.730 12.050 ;
        RECT 1055.510 11.740 1055.890 11.750 ;
        RECT 1103.350 11.740 1103.730 11.750 ;
        RECT 820.910 8.650 821.290 8.660 ;
        RECT 868.750 8.650 869.130 8.660 ;
        RECT 820.910 8.350 869.130 8.650 ;
        RECT 820.910 8.340 821.290 8.350 ;
        RECT 868.750 8.340 869.130 8.350 ;
        RECT 1507.230 5.250 1507.610 5.260 ;
        RECT 1511.830 5.250 1512.210 5.260 ;
        RECT 1507.230 4.950 1512.210 5.250 ;
        RECT 1507.230 4.940 1507.610 4.950 ;
        RECT 1511.830 4.940 1512.210 4.950 ;
      LAYER via3 ;
        RECT 694.900 1746.420 695.220 1746.740 ;
        RECT 1714.260 20.580 1714.580 20.900 ;
        RECT 1804.420 20.580 1804.740 20.900 ;
        RECT 1852.260 15.140 1852.580 15.460 ;
        RECT 2110.780 15.140 2111.100 15.460 ;
        RECT 2200.940 15.140 2201.260 15.460 ;
        RECT 2248.780 15.140 2249.100 15.460 ;
        RECT 2305.820 15.140 2306.140 15.460 ;
        RECT 2498.100 15.140 2498.420 15.460 ;
        RECT 2509.140 15.140 2509.460 15.460 ;
        RECT 741.820 13.780 742.140 14.100 ;
        RECT 785.980 13.780 786.300 14.100 ;
        RECT 1355.460 13.780 1355.780 14.100 ;
        RECT 1234.940 13.100 1235.260 13.420 ;
        RECT 1055.540 11.740 1055.860 12.060 ;
        RECT 1103.380 11.740 1103.700 12.060 ;
        RECT 820.940 8.340 821.260 8.660 ;
        RECT 868.780 8.340 869.100 8.660 ;
        RECT 1507.260 4.940 1507.580 5.260 ;
        RECT 1511.860 4.940 1512.180 5.260 ;
      LAYER met4 ;
        RECT 694.895 1746.415 695.225 1746.745 ;
        RECT 694.910 15.890 695.210 1746.415 ;
        RECT 1714.255 20.575 1714.585 20.905 ;
        RECT 1804.415 20.575 1804.745 20.905 ;
        RECT 1234.510 18.110 1235.690 19.290 ;
        RECT 694.470 14.710 695.650 15.890 ;
        RECT 741.390 14.710 742.570 15.890 ;
        RECT 868.350 14.710 869.530 15.890 ;
        RECT 1102.950 14.710 1104.130 15.890 ;
        RECT 1112.150 15.450 1113.330 15.890 ;
        RECT 1112.150 15.150 1114.730 15.450 ;
        RECT 1112.150 14.710 1113.330 15.150 ;
        RECT 741.830 14.105 742.130 14.710 ;
        RECT 741.815 13.775 742.145 14.105 ;
        RECT 785.975 13.775 786.305 14.105 ;
        RECT 785.990 12.490 786.290 13.775 ;
        RECT 785.550 11.310 786.730 12.490 ;
        RECT 820.510 7.910 821.690 9.090 ;
        RECT 868.790 8.665 869.090 14.710 ;
        RECT 1055.110 11.310 1056.290 12.490 ;
        RECT 1103.390 12.065 1103.690 14.710 ;
        RECT 1114.430 12.490 1114.730 15.150 ;
        RECT 1234.950 13.425 1235.250 18.110 ;
        RECT 1714.270 15.890 1714.570 20.575 ;
        RECT 1675.190 15.450 1676.370 15.890 ;
        RECT 1673.790 15.150 1676.370 15.450 ;
        RECT 1355.455 13.775 1355.785 14.105 ;
        RECT 1234.935 13.095 1235.265 13.425 ;
        RECT 1355.470 12.490 1355.770 13.775 ;
        RECT 1673.790 12.490 1674.090 15.150 ;
        RECT 1675.190 14.710 1676.370 15.150 ;
        RECT 1713.830 14.710 1715.010 15.890 ;
        RECT 1103.375 11.735 1103.705 12.065 ;
        RECT 1113.990 11.310 1115.170 12.490 ;
        RECT 1355.030 11.310 1356.210 12.490 ;
        RECT 1673.350 11.310 1674.530 12.490 ;
        RECT 1804.430 9.090 1804.730 20.575 ;
        RECT 1852.255 15.135 1852.585 15.465 ;
        RECT 2110.775 15.135 2111.105 15.465 ;
        RECT 2200.935 15.135 2201.265 15.465 ;
        RECT 1852.270 9.090 1852.570 15.135 ;
        RECT 2110.790 12.490 2111.090 15.135 ;
        RECT 2200.950 12.490 2201.250 15.135 ;
        RECT 2248.350 14.710 2249.530 15.890 ;
        RECT 2305.390 14.710 2306.570 15.890 ;
        RECT 2497.670 14.710 2498.850 15.890 ;
        RECT 2508.710 14.710 2509.890 15.890 ;
        RECT 2110.350 11.310 2111.530 12.490 ;
        RECT 2200.510 11.310 2201.690 12.490 ;
        RECT 868.775 8.335 869.105 8.665 ;
        RECT 1803.990 7.910 1805.170 9.090 ;
        RECT 1851.830 7.910 1853.010 9.090 ;
        RECT 1506.830 4.510 1508.010 5.690 ;
        RECT 1511.430 4.510 1512.610 5.690 ;
      LAYER met5 ;
        RECT 939.900 17.900 974.620 19.500 ;
        RECT 694.260 14.500 742.780 16.100 ;
        RECT 868.140 14.500 904.700 16.100 ;
        RECT 785.340 11.100 820.980 12.700 ;
        RECT 819.380 9.300 820.980 11.100 ;
        RECT 903.100 9.300 904.700 14.500 ;
        RECT 939.900 9.300 941.500 17.900 ;
        RECT 973.020 12.700 974.620 17.900 ;
        RECT 1216.820 17.900 1235.900 19.500 ;
        RECT 1102.740 14.500 1113.540 16.100 ;
        RECT 1216.820 12.700 1218.420 17.900 ;
        RECT 1674.980 14.500 1715.220 16.100 ;
        RECT 2110.140 14.500 2201.900 16.100 ;
        RECT 2248.140 14.500 2306.780 16.100 ;
        RECT 2497.460 14.500 2510.100 16.100 ;
        RECT 973.020 11.100 1007.740 12.700 ;
        RECT 819.380 7.700 822.680 9.300 ;
        RECT 903.100 7.700 941.500 9.300 ;
        RECT 1006.140 9.300 1007.740 11.100 ;
        RECT 1023.620 11.100 1056.500 12.700 ;
        RECT 1113.780 11.100 1218.420 12.700 ;
        RECT 1354.820 11.100 1429.100 12.700 ;
        RECT 1023.620 9.300 1025.220 11.100 ;
        RECT 1006.140 7.700 1025.220 9.300 ;
        RECT 1427.500 9.300 1429.100 11.100 ;
        RECT 1558.140 11.100 1674.740 12.700 ;
        RECT 2110.140 11.100 2111.740 14.500 ;
        RECT 2200.300 11.100 2201.900 14.500 ;
        RECT 1427.500 7.700 1476.940 9.300 ;
        RECT 1475.340 5.900 1476.940 7.700 ;
        RECT 1558.140 5.900 1559.740 11.100 ;
        RECT 1803.780 7.700 1853.220 9.300 ;
        RECT 1475.340 4.300 1508.220 5.900 ;
        RECT 1511.220 4.300 1559.740 5.900 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2539.345 1538.925 2539.515 1587.035 ;
        RECT 2539.345 1442.025 2539.515 1490.475 ;
        RECT 2539.345 910.945 2539.515 959.055 ;
        RECT 2539.805 814.385 2539.975 862.495 ;
        RECT 2539.345 766.105 2539.515 814.215 ;
        RECT 2539.805 717.825 2539.975 765.595 ;
        RECT 2539.345 669.545 2539.515 717.655 ;
        RECT 2539.345 620.925 2539.515 669.035 ;
        RECT 2539.345 476.425 2539.515 524.195 ;
        RECT 2539.345 427.805 2539.515 475.915 ;
        RECT 2539.345 283.305 2539.515 331.075 ;
        RECT 2539.345 186.745 2539.515 234.515 ;
        RECT 2539.345 138.465 2539.515 186.235 ;
        RECT 2539.345 90.185 2539.515 137.955 ;
      LAYER mcon ;
        RECT 2539.345 1586.865 2539.515 1587.035 ;
        RECT 2539.345 1490.305 2539.515 1490.475 ;
        RECT 2539.345 958.885 2539.515 959.055 ;
        RECT 2539.805 862.325 2539.975 862.495 ;
        RECT 2539.345 814.045 2539.515 814.215 ;
        RECT 2539.805 765.425 2539.975 765.595 ;
        RECT 2539.345 717.485 2539.515 717.655 ;
        RECT 2539.345 668.865 2539.515 669.035 ;
        RECT 2539.345 524.025 2539.515 524.195 ;
        RECT 2539.345 475.745 2539.515 475.915 ;
        RECT 2539.345 330.905 2539.515 331.075 ;
        RECT 2539.345 234.345 2539.515 234.515 ;
        RECT 2539.345 186.065 2539.515 186.235 ;
        RECT 2539.345 137.785 2539.515 137.955 ;
      LAYER met1 ;
        RECT 1772.910 1600.960 1773.230 1601.020 ;
        RECT 2539.270 1600.960 2539.590 1601.020 ;
        RECT 1772.910 1600.820 2539.590 1600.960 ;
        RECT 1772.910 1600.760 1773.230 1600.820 ;
        RECT 2539.270 1600.760 2539.590 1600.820 ;
        RECT 2539.270 1587.020 2539.590 1587.080 ;
        RECT 2539.075 1586.880 2539.590 1587.020 ;
        RECT 2539.270 1586.820 2539.590 1586.880 ;
        RECT 2539.270 1539.080 2539.590 1539.140 ;
        RECT 2539.075 1538.940 2539.590 1539.080 ;
        RECT 2539.270 1538.880 2539.590 1538.940 ;
        RECT 2539.270 1490.460 2539.590 1490.520 ;
        RECT 2539.075 1490.320 2539.590 1490.460 ;
        RECT 2539.270 1490.260 2539.590 1490.320 ;
        RECT 2539.270 1442.180 2539.590 1442.240 ;
        RECT 2539.075 1442.040 2539.590 1442.180 ;
        RECT 2539.270 1441.980 2539.590 1442.040 ;
        RECT 2539.270 1345.620 2539.590 1345.680 ;
        RECT 2540.190 1345.620 2540.510 1345.680 ;
        RECT 2539.270 1345.480 2540.510 1345.620 ;
        RECT 2539.270 1345.420 2539.590 1345.480 ;
        RECT 2540.190 1345.420 2540.510 1345.480 ;
        RECT 2539.270 1249.060 2539.590 1249.120 ;
        RECT 2540.190 1249.060 2540.510 1249.120 ;
        RECT 2539.270 1248.920 2540.510 1249.060 ;
        RECT 2539.270 1248.860 2539.590 1248.920 ;
        RECT 2540.190 1248.860 2540.510 1248.920 ;
        RECT 2537.890 1055.600 2538.210 1055.660 ;
        RECT 2538.810 1055.600 2539.130 1055.660 ;
        RECT 2537.890 1055.460 2539.130 1055.600 ;
        RECT 2537.890 1055.400 2538.210 1055.460 ;
        RECT 2538.810 1055.400 2539.130 1055.460 ;
        RECT 2537.890 1007.320 2538.210 1007.380 ;
        RECT 2539.270 1007.320 2539.590 1007.380 ;
        RECT 2537.890 1007.180 2539.590 1007.320 ;
        RECT 2537.890 1007.120 2538.210 1007.180 ;
        RECT 2539.270 1007.120 2539.590 1007.180 ;
        RECT 2539.270 959.040 2539.590 959.100 ;
        RECT 2539.075 958.900 2539.590 959.040 ;
        RECT 2539.270 958.840 2539.590 958.900 ;
        RECT 2539.270 911.100 2539.590 911.160 ;
        RECT 2539.075 910.960 2539.590 911.100 ;
        RECT 2539.270 910.900 2539.590 910.960 ;
        RECT 2537.890 910.420 2538.210 910.480 ;
        RECT 2539.270 910.420 2539.590 910.480 ;
        RECT 2537.890 910.280 2539.590 910.420 ;
        RECT 2537.890 910.220 2538.210 910.280 ;
        RECT 2539.270 910.220 2539.590 910.280 ;
        RECT 2539.270 862.480 2539.590 862.540 ;
        RECT 2539.745 862.480 2540.035 862.525 ;
        RECT 2539.270 862.340 2540.035 862.480 ;
        RECT 2539.270 862.280 2539.590 862.340 ;
        RECT 2539.745 862.295 2540.035 862.340 ;
        RECT 2539.730 814.540 2540.050 814.600 ;
        RECT 2539.535 814.400 2540.050 814.540 ;
        RECT 2539.730 814.340 2540.050 814.400 ;
        RECT 2539.270 814.200 2539.590 814.260 ;
        RECT 2539.075 814.060 2539.590 814.200 ;
        RECT 2539.270 814.000 2539.590 814.060 ;
        RECT 2539.285 766.260 2539.575 766.305 ;
        RECT 2539.730 766.260 2540.050 766.320 ;
        RECT 2539.285 766.120 2540.050 766.260 ;
        RECT 2539.285 766.075 2539.575 766.120 ;
        RECT 2539.730 766.060 2540.050 766.120 ;
        RECT 2539.270 765.580 2539.590 765.640 ;
        RECT 2539.745 765.580 2540.035 765.625 ;
        RECT 2539.270 765.440 2540.035 765.580 ;
        RECT 2539.270 765.380 2539.590 765.440 ;
        RECT 2539.745 765.395 2540.035 765.440 ;
        RECT 2539.730 717.980 2540.050 718.040 ;
        RECT 2539.535 717.840 2540.050 717.980 ;
        RECT 2539.730 717.780 2540.050 717.840 ;
        RECT 2539.270 717.640 2539.590 717.700 ;
        RECT 2539.075 717.500 2539.590 717.640 ;
        RECT 2539.270 717.440 2539.590 717.500 ;
        RECT 2538.810 669.700 2539.130 669.760 ;
        RECT 2539.285 669.700 2539.575 669.745 ;
        RECT 2538.810 669.560 2539.575 669.700 ;
        RECT 2538.810 669.500 2539.130 669.560 ;
        RECT 2539.285 669.515 2539.575 669.560 ;
        RECT 2539.270 669.020 2539.590 669.080 ;
        RECT 2539.075 668.880 2539.590 669.020 ;
        RECT 2539.270 668.820 2539.590 668.880 ;
        RECT 2539.270 621.080 2539.590 621.140 ;
        RECT 2539.075 620.940 2539.590 621.080 ;
        RECT 2539.270 620.880 2539.590 620.940 ;
        RECT 2538.350 572.460 2538.670 572.520 ;
        RECT 2539.270 572.460 2539.590 572.520 ;
        RECT 2538.350 572.320 2539.590 572.460 ;
        RECT 2538.350 572.260 2538.670 572.320 ;
        RECT 2539.270 572.260 2539.590 572.320 ;
        RECT 2539.270 524.180 2539.590 524.240 ;
        RECT 2539.075 524.040 2539.590 524.180 ;
        RECT 2539.270 523.980 2539.590 524.040 ;
        RECT 2539.285 476.580 2539.575 476.625 ;
        RECT 2539.730 476.580 2540.050 476.640 ;
        RECT 2539.285 476.440 2540.050 476.580 ;
        RECT 2539.285 476.395 2539.575 476.440 ;
        RECT 2539.730 476.380 2540.050 476.440 ;
        RECT 2539.270 475.900 2539.590 475.960 ;
        RECT 2539.075 475.760 2539.590 475.900 ;
        RECT 2539.270 475.700 2539.590 475.760 ;
        RECT 2539.270 427.960 2539.590 428.020 ;
        RECT 2539.075 427.820 2539.590 427.960 ;
        RECT 2539.270 427.760 2539.590 427.820 ;
        RECT 2538.350 379.340 2538.670 379.400 ;
        RECT 2539.270 379.340 2539.590 379.400 ;
        RECT 2538.350 379.200 2539.590 379.340 ;
        RECT 2538.350 379.140 2538.670 379.200 ;
        RECT 2539.270 379.140 2539.590 379.200 ;
        RECT 2539.270 331.060 2539.590 331.120 ;
        RECT 2539.075 330.920 2539.590 331.060 ;
        RECT 2539.270 330.860 2539.590 330.920 ;
        RECT 2539.285 283.460 2539.575 283.505 ;
        RECT 2539.730 283.460 2540.050 283.520 ;
        RECT 2539.285 283.320 2540.050 283.460 ;
        RECT 2539.285 283.275 2539.575 283.320 ;
        RECT 2539.730 283.260 2540.050 283.320 ;
        RECT 2538.350 282.780 2538.670 282.840 ;
        RECT 2539.270 282.780 2539.590 282.840 ;
        RECT 2538.350 282.640 2539.590 282.780 ;
        RECT 2538.350 282.580 2538.670 282.640 ;
        RECT 2539.270 282.580 2539.590 282.640 ;
        RECT 2539.270 234.500 2539.590 234.560 ;
        RECT 2539.075 234.360 2539.590 234.500 ;
        RECT 2539.270 234.300 2539.590 234.360 ;
        RECT 2539.285 186.900 2539.575 186.945 ;
        RECT 2539.730 186.900 2540.050 186.960 ;
        RECT 2539.285 186.760 2540.050 186.900 ;
        RECT 2539.285 186.715 2539.575 186.760 ;
        RECT 2539.730 186.700 2540.050 186.760 ;
        RECT 2539.270 186.220 2539.590 186.280 ;
        RECT 2539.075 186.080 2539.590 186.220 ;
        RECT 2539.270 186.020 2539.590 186.080 ;
        RECT 2539.270 138.620 2539.590 138.680 ;
        RECT 2539.075 138.480 2539.590 138.620 ;
        RECT 2539.270 138.420 2539.590 138.480 ;
        RECT 2539.270 137.940 2539.590 138.000 ;
        RECT 2539.075 137.800 2539.590 137.940 ;
        RECT 2539.270 137.740 2539.590 137.800 ;
        RECT 2539.285 90.340 2539.575 90.385 ;
        RECT 2539.730 90.340 2540.050 90.400 ;
        RECT 2539.285 90.200 2540.050 90.340 ;
        RECT 2539.285 90.155 2539.575 90.200 ;
        RECT 2539.730 90.140 2540.050 90.200 ;
        RECT 2539.270 89.660 2539.590 89.720 ;
        RECT 2541.110 89.660 2541.430 89.720 ;
        RECT 2539.270 89.520 2541.430 89.660 ;
        RECT 2539.270 89.460 2539.590 89.520 ;
        RECT 2541.110 89.460 2541.430 89.520 ;
        RECT 2541.110 2.960 2541.430 3.020 ;
        RECT 2542.030 2.960 2542.350 3.020 ;
        RECT 2541.110 2.820 2542.350 2.960 ;
        RECT 2541.110 2.760 2541.430 2.820 ;
        RECT 2542.030 2.760 2542.350 2.820 ;
      LAYER via ;
        RECT 1772.940 1600.760 1773.200 1601.020 ;
        RECT 2539.300 1600.760 2539.560 1601.020 ;
        RECT 2539.300 1586.820 2539.560 1587.080 ;
        RECT 2539.300 1538.880 2539.560 1539.140 ;
        RECT 2539.300 1490.260 2539.560 1490.520 ;
        RECT 2539.300 1441.980 2539.560 1442.240 ;
        RECT 2539.300 1345.420 2539.560 1345.680 ;
        RECT 2540.220 1345.420 2540.480 1345.680 ;
        RECT 2539.300 1248.860 2539.560 1249.120 ;
        RECT 2540.220 1248.860 2540.480 1249.120 ;
        RECT 2537.920 1055.400 2538.180 1055.660 ;
        RECT 2538.840 1055.400 2539.100 1055.660 ;
        RECT 2537.920 1007.120 2538.180 1007.380 ;
        RECT 2539.300 1007.120 2539.560 1007.380 ;
        RECT 2539.300 958.840 2539.560 959.100 ;
        RECT 2539.300 910.900 2539.560 911.160 ;
        RECT 2537.920 910.220 2538.180 910.480 ;
        RECT 2539.300 910.220 2539.560 910.480 ;
        RECT 2539.300 862.280 2539.560 862.540 ;
        RECT 2539.760 814.340 2540.020 814.600 ;
        RECT 2539.300 814.000 2539.560 814.260 ;
        RECT 2539.760 766.060 2540.020 766.320 ;
        RECT 2539.300 765.380 2539.560 765.640 ;
        RECT 2539.760 717.780 2540.020 718.040 ;
        RECT 2539.300 717.440 2539.560 717.700 ;
        RECT 2538.840 669.500 2539.100 669.760 ;
        RECT 2539.300 668.820 2539.560 669.080 ;
        RECT 2539.300 620.880 2539.560 621.140 ;
        RECT 2538.380 572.260 2538.640 572.520 ;
        RECT 2539.300 572.260 2539.560 572.520 ;
        RECT 2539.300 523.980 2539.560 524.240 ;
        RECT 2539.760 476.380 2540.020 476.640 ;
        RECT 2539.300 475.700 2539.560 475.960 ;
        RECT 2539.300 427.760 2539.560 428.020 ;
        RECT 2538.380 379.140 2538.640 379.400 ;
        RECT 2539.300 379.140 2539.560 379.400 ;
        RECT 2539.300 330.860 2539.560 331.120 ;
        RECT 2539.760 283.260 2540.020 283.520 ;
        RECT 2538.380 282.580 2538.640 282.840 ;
        RECT 2539.300 282.580 2539.560 282.840 ;
        RECT 2539.300 234.300 2539.560 234.560 ;
        RECT 2539.760 186.700 2540.020 186.960 ;
        RECT 2539.300 186.020 2539.560 186.280 ;
        RECT 2539.300 138.420 2539.560 138.680 ;
        RECT 2539.300 137.740 2539.560 138.000 ;
        RECT 2539.760 90.140 2540.020 90.400 ;
        RECT 2539.300 89.460 2539.560 89.720 ;
        RECT 2541.140 89.460 2541.400 89.720 ;
        RECT 2541.140 2.760 2541.400 3.020 ;
        RECT 2542.060 2.760 2542.320 3.020 ;
      LAYER met2 ;
        RECT 1772.930 1604.955 1773.210 1605.325 ;
        RECT 1773.000 1601.050 1773.140 1604.955 ;
        RECT 1772.940 1600.730 1773.200 1601.050 ;
        RECT 2539.300 1600.730 2539.560 1601.050 ;
        RECT 2539.360 1587.110 2539.500 1600.730 ;
        RECT 2539.300 1586.790 2539.560 1587.110 ;
        RECT 2539.300 1538.850 2539.560 1539.170 ;
        RECT 2539.360 1490.550 2539.500 1538.850 ;
        RECT 2539.300 1490.230 2539.560 1490.550 ;
        RECT 2539.300 1441.950 2539.560 1442.270 ;
        RECT 2539.360 1393.845 2539.500 1441.950 ;
        RECT 2539.290 1393.475 2539.570 1393.845 ;
        RECT 2540.210 1393.475 2540.490 1393.845 ;
        RECT 2540.280 1345.710 2540.420 1393.475 ;
        RECT 2539.300 1345.390 2539.560 1345.710 ;
        RECT 2540.220 1345.390 2540.480 1345.710 ;
        RECT 2539.360 1297.285 2539.500 1345.390 ;
        RECT 2539.290 1296.915 2539.570 1297.285 ;
        RECT 2540.210 1296.915 2540.490 1297.285 ;
        RECT 2540.280 1249.150 2540.420 1296.915 ;
        RECT 2539.300 1248.830 2539.560 1249.150 ;
        RECT 2540.220 1248.830 2540.480 1249.150 ;
        RECT 2539.360 1208.885 2539.500 1248.830 ;
        RECT 2539.290 1208.515 2539.570 1208.885 ;
        RECT 2539.290 1207.835 2539.570 1208.205 ;
        RECT 2539.360 1104.165 2539.500 1207.835 ;
        RECT 2537.910 1103.795 2538.190 1104.165 ;
        RECT 2539.290 1103.795 2539.570 1104.165 ;
        RECT 2537.980 1055.885 2538.120 1103.795 ;
        RECT 2537.910 1055.515 2538.190 1055.885 ;
        RECT 2538.830 1055.515 2539.110 1055.885 ;
        RECT 2537.920 1055.370 2538.180 1055.515 ;
        RECT 2538.840 1055.370 2539.100 1055.515 ;
        RECT 2537.980 1007.605 2538.120 1055.370 ;
        RECT 2537.910 1007.235 2538.190 1007.605 ;
        RECT 2539.290 1007.235 2539.570 1007.605 ;
        RECT 2537.920 1007.090 2538.180 1007.235 ;
        RECT 2539.300 1007.090 2539.560 1007.235 ;
        RECT 2537.980 959.325 2538.120 1007.090 ;
        RECT 2537.910 958.955 2538.190 959.325 ;
        RECT 2538.830 959.210 2539.110 959.325 ;
        RECT 2538.830 959.130 2539.500 959.210 ;
        RECT 2538.830 959.070 2539.560 959.130 ;
        RECT 2538.830 958.955 2539.110 959.070 ;
        RECT 2539.300 958.810 2539.560 959.070 ;
        RECT 2539.360 958.655 2539.500 958.810 ;
        RECT 2539.300 910.870 2539.560 911.190 ;
        RECT 2539.360 910.510 2539.500 910.870 ;
        RECT 2537.920 910.190 2538.180 910.510 ;
        RECT 2539.300 910.190 2539.560 910.510 ;
        RECT 2537.980 862.765 2538.120 910.190 ;
        RECT 2537.910 862.395 2538.190 862.765 ;
        RECT 2538.830 862.650 2539.110 862.765 ;
        RECT 2538.830 862.570 2539.500 862.650 ;
        RECT 2538.830 862.510 2539.560 862.570 ;
        RECT 2538.830 862.395 2539.110 862.510 ;
        RECT 2539.300 862.250 2539.560 862.510 ;
        RECT 2539.360 862.095 2539.500 862.250 ;
        RECT 2539.760 814.370 2540.020 814.630 ;
        RECT 2539.360 814.310 2540.020 814.370 ;
        RECT 2539.360 814.290 2539.960 814.310 ;
        RECT 2539.300 814.230 2539.960 814.290 ;
        RECT 2539.300 813.970 2539.560 814.230 ;
        RECT 2539.760 766.090 2540.020 766.350 ;
        RECT 2539.360 766.030 2540.020 766.090 ;
        RECT 2539.360 765.950 2539.960 766.030 ;
        RECT 2539.360 765.670 2539.500 765.950 ;
        RECT 2539.300 765.350 2539.560 765.670 ;
        RECT 2539.760 717.810 2540.020 718.070 ;
        RECT 2539.360 717.750 2540.020 717.810 ;
        RECT 2539.360 717.730 2539.960 717.750 ;
        RECT 2539.300 717.670 2539.960 717.730 ;
        RECT 2539.300 717.410 2539.560 717.670 ;
        RECT 2538.840 669.530 2539.100 669.790 ;
        RECT 2538.840 669.470 2539.500 669.530 ;
        RECT 2538.900 669.390 2539.500 669.470 ;
        RECT 2539.360 669.110 2539.500 669.390 ;
        RECT 2539.300 668.790 2539.560 669.110 ;
        RECT 2539.300 620.850 2539.560 621.170 ;
        RECT 2539.360 620.685 2539.500 620.850 ;
        RECT 2539.290 620.315 2539.570 620.685 ;
        RECT 2540.670 619.635 2540.950 620.005 ;
        RECT 2540.740 573.085 2540.880 619.635 ;
        RECT 2539.750 572.970 2540.030 573.085 ;
        RECT 2539.360 572.830 2540.030 572.970 ;
        RECT 2539.360 572.550 2539.500 572.830 ;
        RECT 2539.750 572.715 2540.030 572.830 ;
        RECT 2540.670 572.715 2540.950 573.085 ;
        RECT 2538.380 572.230 2538.640 572.550 ;
        RECT 2539.300 572.230 2539.560 572.550 ;
        RECT 2538.440 524.805 2538.580 572.230 ;
        RECT 2538.370 524.435 2538.650 524.805 ;
        RECT 2539.290 524.435 2539.570 524.805 ;
        RECT 2539.360 524.270 2539.500 524.435 ;
        RECT 2539.300 523.950 2539.560 524.270 ;
        RECT 2539.760 476.410 2540.020 476.670 ;
        RECT 2539.360 476.350 2540.020 476.410 ;
        RECT 2539.360 476.270 2539.960 476.350 ;
        RECT 2539.360 475.990 2539.500 476.270 ;
        RECT 2539.300 475.670 2539.560 475.990 ;
        RECT 2539.300 427.730 2539.560 428.050 ;
        RECT 2539.360 379.430 2539.500 427.730 ;
        RECT 2538.380 379.110 2538.640 379.430 ;
        RECT 2539.300 379.110 2539.560 379.430 ;
        RECT 2538.440 331.685 2538.580 379.110 ;
        RECT 2538.370 331.315 2538.650 331.685 ;
        RECT 2539.290 331.315 2539.570 331.685 ;
        RECT 2539.360 331.150 2539.500 331.315 ;
        RECT 2539.300 330.830 2539.560 331.150 ;
        RECT 2539.760 283.290 2540.020 283.550 ;
        RECT 2539.360 283.230 2540.020 283.290 ;
        RECT 2539.360 283.150 2539.960 283.230 ;
        RECT 2539.360 282.870 2539.500 283.150 ;
        RECT 2538.380 282.550 2538.640 282.870 ;
        RECT 2539.300 282.550 2539.560 282.870 ;
        RECT 2538.440 235.125 2538.580 282.550 ;
        RECT 2538.370 234.755 2538.650 235.125 ;
        RECT 2539.290 234.755 2539.570 235.125 ;
        RECT 2539.360 234.590 2539.500 234.755 ;
        RECT 2539.300 234.270 2539.560 234.590 ;
        RECT 2539.760 186.730 2540.020 186.990 ;
        RECT 2539.360 186.670 2540.020 186.730 ;
        RECT 2539.360 186.590 2539.960 186.670 ;
        RECT 2539.360 186.310 2539.500 186.590 ;
        RECT 2539.300 185.990 2539.560 186.310 ;
        RECT 2539.300 138.390 2539.560 138.710 ;
        RECT 2539.360 138.030 2539.500 138.390 ;
        RECT 2539.300 137.710 2539.560 138.030 ;
        RECT 2539.760 90.170 2540.020 90.430 ;
        RECT 2539.360 90.110 2540.020 90.170 ;
        RECT 2539.360 90.030 2539.960 90.110 ;
        RECT 2539.360 89.750 2539.500 90.030 ;
        RECT 2539.300 89.430 2539.560 89.750 ;
        RECT 2541.140 89.430 2541.400 89.750 ;
        RECT 2541.200 3.050 2541.340 89.430 ;
        RECT 2541.140 2.730 2541.400 3.050 ;
        RECT 2542.060 2.730 2542.320 3.050 ;
        RECT 2542.120 2.400 2542.260 2.730 ;
        RECT 2541.910 -4.800 2542.470 2.400 ;
      LAYER via2 ;
        RECT 1772.930 1605.000 1773.210 1605.280 ;
        RECT 2539.290 1393.520 2539.570 1393.800 ;
        RECT 2540.210 1393.520 2540.490 1393.800 ;
        RECT 2539.290 1296.960 2539.570 1297.240 ;
        RECT 2540.210 1296.960 2540.490 1297.240 ;
        RECT 2539.290 1208.560 2539.570 1208.840 ;
        RECT 2539.290 1207.880 2539.570 1208.160 ;
        RECT 2537.910 1103.840 2538.190 1104.120 ;
        RECT 2539.290 1103.840 2539.570 1104.120 ;
        RECT 2537.910 1055.560 2538.190 1055.840 ;
        RECT 2538.830 1055.560 2539.110 1055.840 ;
        RECT 2537.910 1007.280 2538.190 1007.560 ;
        RECT 2539.290 1007.280 2539.570 1007.560 ;
        RECT 2537.910 959.000 2538.190 959.280 ;
        RECT 2538.830 959.000 2539.110 959.280 ;
        RECT 2537.910 862.440 2538.190 862.720 ;
        RECT 2538.830 862.440 2539.110 862.720 ;
        RECT 2539.290 620.360 2539.570 620.640 ;
        RECT 2540.670 619.680 2540.950 619.960 ;
        RECT 2539.750 572.760 2540.030 573.040 ;
        RECT 2540.670 572.760 2540.950 573.040 ;
        RECT 2538.370 524.480 2538.650 524.760 ;
        RECT 2539.290 524.480 2539.570 524.760 ;
        RECT 2538.370 331.360 2538.650 331.640 ;
        RECT 2539.290 331.360 2539.570 331.640 ;
        RECT 2538.370 234.800 2538.650 235.080 ;
        RECT 2539.290 234.800 2539.570 235.080 ;
      LAYER met3 ;
        RECT 1755.835 1605.290 1759.835 1605.295 ;
        RECT 1772.905 1605.290 1773.235 1605.305 ;
        RECT 1755.835 1604.990 1773.235 1605.290 ;
        RECT 1755.835 1604.695 1759.835 1604.990 ;
        RECT 1772.905 1604.975 1773.235 1604.990 ;
        RECT 2539.265 1393.810 2539.595 1393.825 ;
        RECT 2540.185 1393.810 2540.515 1393.825 ;
        RECT 2539.265 1393.510 2540.515 1393.810 ;
        RECT 2539.265 1393.495 2539.595 1393.510 ;
        RECT 2540.185 1393.495 2540.515 1393.510 ;
        RECT 2539.265 1297.250 2539.595 1297.265 ;
        RECT 2540.185 1297.250 2540.515 1297.265 ;
        RECT 2539.265 1296.950 2540.515 1297.250 ;
        RECT 2539.265 1296.935 2539.595 1296.950 ;
        RECT 2540.185 1296.935 2540.515 1296.950 ;
        RECT 2539.265 1208.850 2539.595 1208.865 ;
        RECT 2538.590 1208.550 2539.595 1208.850 ;
        RECT 2538.590 1208.170 2538.890 1208.550 ;
        RECT 2539.265 1208.535 2539.595 1208.550 ;
        RECT 2539.265 1208.170 2539.595 1208.185 ;
        RECT 2538.590 1207.870 2539.595 1208.170 ;
        RECT 2539.265 1207.855 2539.595 1207.870 ;
        RECT 2537.885 1104.130 2538.215 1104.145 ;
        RECT 2539.265 1104.130 2539.595 1104.145 ;
        RECT 2537.885 1103.830 2539.595 1104.130 ;
        RECT 2537.885 1103.815 2538.215 1103.830 ;
        RECT 2539.265 1103.815 2539.595 1103.830 ;
        RECT 2537.885 1055.850 2538.215 1055.865 ;
        RECT 2538.805 1055.850 2539.135 1055.865 ;
        RECT 2537.885 1055.550 2539.135 1055.850 ;
        RECT 2537.885 1055.535 2538.215 1055.550 ;
        RECT 2538.805 1055.535 2539.135 1055.550 ;
        RECT 2537.885 1007.570 2538.215 1007.585 ;
        RECT 2539.265 1007.570 2539.595 1007.585 ;
        RECT 2537.885 1007.270 2539.595 1007.570 ;
        RECT 2537.885 1007.255 2538.215 1007.270 ;
        RECT 2539.265 1007.255 2539.595 1007.270 ;
        RECT 2537.885 959.290 2538.215 959.305 ;
        RECT 2538.805 959.290 2539.135 959.305 ;
        RECT 2537.885 958.990 2539.135 959.290 ;
        RECT 2537.885 958.975 2538.215 958.990 ;
        RECT 2538.805 958.975 2539.135 958.990 ;
        RECT 2537.885 862.730 2538.215 862.745 ;
        RECT 2538.805 862.730 2539.135 862.745 ;
        RECT 2537.885 862.430 2539.135 862.730 ;
        RECT 2537.885 862.415 2538.215 862.430 ;
        RECT 2538.805 862.415 2539.135 862.430 ;
        RECT 2539.265 620.650 2539.595 620.665 ;
        RECT 2538.590 620.350 2539.595 620.650 ;
        RECT 2538.590 619.970 2538.890 620.350 ;
        RECT 2539.265 620.335 2539.595 620.350 ;
        RECT 2540.645 619.970 2540.975 619.985 ;
        RECT 2538.590 619.670 2540.975 619.970 ;
        RECT 2540.645 619.655 2540.975 619.670 ;
        RECT 2539.725 573.050 2540.055 573.065 ;
        RECT 2540.645 573.050 2540.975 573.065 ;
        RECT 2539.725 572.750 2540.975 573.050 ;
        RECT 2539.725 572.735 2540.055 572.750 ;
        RECT 2540.645 572.735 2540.975 572.750 ;
        RECT 2538.345 524.770 2538.675 524.785 ;
        RECT 2539.265 524.770 2539.595 524.785 ;
        RECT 2538.345 524.470 2539.595 524.770 ;
        RECT 2538.345 524.455 2538.675 524.470 ;
        RECT 2539.265 524.455 2539.595 524.470 ;
        RECT 2538.345 331.650 2538.675 331.665 ;
        RECT 2539.265 331.650 2539.595 331.665 ;
        RECT 2538.345 331.350 2539.595 331.650 ;
        RECT 2538.345 331.335 2538.675 331.350 ;
        RECT 2539.265 331.335 2539.595 331.350 ;
        RECT 2538.345 235.090 2538.675 235.105 ;
        RECT 2539.265 235.090 2539.595 235.105 ;
        RECT 2538.345 234.790 2539.595 235.090 ;
        RECT 2538.345 234.775 2538.675 234.790 ;
        RECT 2539.265 234.775 2539.595 234.790 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1681.830 2380.240 1682.150 2380.300 ;
        RECT 2559.970 2380.240 2560.290 2380.300 ;
        RECT 1681.830 2380.100 2560.290 2380.240 ;
        RECT 1681.830 2380.040 1682.150 2380.100 ;
        RECT 2559.970 2380.040 2560.290 2380.100 ;
      LAYER via ;
        RECT 1681.860 2380.040 1682.120 2380.300 ;
        RECT 2560.000 2380.040 2560.260 2380.300 ;
      LAYER met2 ;
        RECT 1681.860 2380.010 1682.120 2380.330 ;
        RECT 2560.000 2380.010 2560.260 2380.330 ;
        RECT 1681.920 2377.880 1682.060 2380.010 ;
        RECT 1681.900 2373.880 1682.180 2377.880 ;
        RECT 2560.060 2.400 2560.200 2380.010 ;
        RECT 2559.850 -4.800 2560.410 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2577.930 16.475 2578.210 16.845 ;
        RECT 2578.000 2.400 2578.140 16.475 ;
        RECT 2577.790 -4.800 2578.350 2.400 ;
      LAYER via2 ;
        RECT 2577.930 16.520 2578.210 16.800 ;
      LAYER met3 ;
        RECT 693.950 1677.370 694.330 1677.380 ;
        RECT 715.810 1677.370 719.810 1677.375 ;
        RECT 693.950 1677.070 719.810 1677.370 ;
        RECT 693.950 1677.060 694.330 1677.070 ;
        RECT 715.810 1676.775 719.810 1677.070 ;
        RECT 693.950 16.810 694.330 16.820 ;
        RECT 2577.905 16.810 2578.235 16.825 ;
        RECT 693.950 16.510 2578.235 16.810 ;
        RECT 693.950 16.500 694.330 16.510 ;
        RECT 2577.905 16.495 2578.235 16.510 ;
      LAYER via3 ;
        RECT 693.980 1677.060 694.300 1677.380 ;
        RECT 693.980 16.500 694.300 16.820 ;
      LAYER met4 ;
        RECT 693.975 1677.055 694.305 1677.385 ;
        RECT 693.990 16.825 694.290 1677.055 ;
        RECT 693.975 16.495 694.305 16.825 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 706.705 1427.745 706.875 1430.295 ;
      LAYER mcon ;
        RECT 706.705 1430.125 706.875 1430.295 ;
      LAYER met1 ;
        RECT 706.630 1430.280 706.950 1430.340 ;
        RECT 706.435 1430.140 706.950 1430.280 ;
        RECT 706.630 1430.080 706.950 1430.140 ;
        RECT 706.630 1427.900 706.950 1427.960 ;
        RECT 706.435 1427.760 706.950 1427.900 ;
        RECT 706.630 1427.700 706.950 1427.760 ;
        RECT 688.230 1421.100 688.550 1421.160 ;
        RECT 706.630 1421.100 706.950 1421.160 ;
        RECT 688.230 1420.960 706.950 1421.100 ;
        RECT 688.230 1420.900 688.550 1420.960 ;
        RECT 706.630 1420.900 706.950 1420.960 ;
        RECT 688.230 30.840 688.550 30.900 ;
        RECT 811.510 30.840 811.830 30.900 ;
        RECT 688.230 30.700 811.830 30.840 ;
        RECT 688.230 30.640 688.550 30.700 ;
        RECT 811.510 30.640 811.830 30.700 ;
      LAYER via ;
        RECT 706.660 1430.080 706.920 1430.340 ;
        RECT 706.660 1427.700 706.920 1427.960 ;
        RECT 688.260 1420.900 688.520 1421.160 ;
        RECT 706.660 1420.900 706.920 1421.160 ;
        RECT 688.260 30.640 688.520 30.900 ;
        RECT 811.540 30.640 811.800 30.900 ;
      LAYER met2 ;
        RECT 706.650 2095.915 706.930 2096.285 ;
        RECT 706.720 1430.370 706.860 2095.915 ;
        RECT 706.660 1430.050 706.920 1430.370 ;
        RECT 706.660 1427.670 706.920 1427.990 ;
        RECT 706.720 1421.190 706.860 1427.670 ;
        RECT 688.260 1420.870 688.520 1421.190 ;
        RECT 706.660 1420.870 706.920 1421.190 ;
        RECT 688.320 1393.845 688.460 1420.870 ;
        RECT 688.250 1393.475 688.530 1393.845 ;
        RECT 688.250 1390.755 688.530 1391.125 ;
        RECT 688.320 30.930 688.460 1390.755 ;
        RECT 688.260 30.610 688.520 30.930 ;
        RECT 811.540 30.610 811.800 30.930 ;
        RECT 811.600 2.400 811.740 30.610 ;
        RECT 811.390 -4.800 811.950 2.400 ;
      LAYER via2 ;
        RECT 706.650 2095.960 706.930 2096.240 ;
        RECT 688.250 1393.520 688.530 1393.800 ;
        RECT 688.250 1390.800 688.530 1391.080 ;
      LAYER met3 ;
        RECT 706.625 2096.250 706.955 2096.265 ;
        RECT 715.810 2096.250 719.810 2096.255 ;
        RECT 706.625 2095.950 719.810 2096.250 ;
        RECT 706.625 2095.935 706.955 2095.950 ;
        RECT 715.810 2095.655 719.810 2095.950 ;
        RECT 688.225 1393.810 688.555 1393.825 ;
        RECT 688.225 1393.495 688.770 1393.810 ;
        RECT 688.470 1391.105 688.770 1393.495 ;
        RECT 688.225 1390.790 688.770 1391.105 ;
        RECT 688.225 1390.775 688.555 1390.790 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 737.910 45.120 738.230 45.180 ;
        RECT 2595.390 45.120 2595.710 45.180 ;
        RECT 737.910 44.980 2595.710 45.120 ;
        RECT 737.910 44.920 738.230 44.980 ;
        RECT 2595.390 44.920 2595.710 44.980 ;
      LAYER via ;
        RECT 737.940 44.920 738.200 45.180 ;
        RECT 2595.420 44.920 2595.680 45.180 ;
      LAYER met2 ;
        RECT 735.220 1323.690 735.500 1327.135 ;
        RECT 735.220 1323.550 738.140 1323.690 ;
        RECT 735.220 1323.135 735.500 1323.550 ;
        RECT 738.000 45.210 738.140 1323.550 ;
        RECT 737.940 44.890 738.200 45.210 ;
        RECT 2595.420 44.890 2595.680 45.210 ;
        RECT 2595.480 2.400 2595.620 44.890 ;
        RECT 2595.270 -4.800 2595.830 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 713.070 410.620 713.390 410.680 ;
        RECT 2608.270 410.620 2608.590 410.680 ;
        RECT 713.070 410.480 2608.590 410.620 ;
        RECT 713.070 410.420 713.390 410.480 ;
        RECT 2608.270 410.420 2608.590 410.480 ;
        RECT 2608.270 14.180 2608.590 14.240 ;
        RECT 2608.270 14.040 2613.560 14.180 ;
        RECT 2608.270 13.980 2608.590 14.040 ;
        RECT 2613.420 13.900 2613.560 14.040 ;
        RECT 2613.330 13.640 2613.650 13.900 ;
      LAYER via ;
        RECT 713.100 410.420 713.360 410.680 ;
        RECT 2608.300 410.420 2608.560 410.680 ;
        RECT 2608.300 13.980 2608.560 14.240 ;
        RECT 2613.360 13.640 2613.620 13.900 ;
      LAYER met2 ;
        RECT 713.090 1668.875 713.370 1669.245 ;
        RECT 713.160 410.710 713.300 1668.875 ;
        RECT 713.100 410.390 713.360 410.710 ;
        RECT 2608.300 410.390 2608.560 410.710 ;
        RECT 2608.360 14.270 2608.500 410.390 ;
        RECT 2608.300 13.950 2608.560 14.270 ;
        RECT 2613.360 13.610 2613.620 13.930 ;
        RECT 2613.420 2.400 2613.560 13.610 ;
        RECT 2613.210 -4.800 2613.770 2.400 ;
      LAYER via2 ;
        RECT 713.090 1668.920 713.370 1669.200 ;
      LAYER met3 ;
        RECT 713.065 1669.210 713.395 1669.225 ;
        RECT 715.810 1669.210 719.810 1669.215 ;
        RECT 713.065 1668.910 719.810 1669.210 ;
        RECT 713.065 1668.895 713.395 1668.910 ;
        RECT 715.810 1668.615 719.810 1668.910 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1574.190 1311.280 1574.510 1311.340 ;
        RECT 1579.710 1311.280 1580.030 1311.340 ;
        RECT 1574.190 1311.140 1580.030 1311.280 ;
        RECT 1574.190 1311.080 1574.510 1311.140 ;
        RECT 1579.710 1311.080 1580.030 1311.140 ;
        RECT 1579.710 46.140 1580.030 46.200 ;
        RECT 2631.270 46.140 2631.590 46.200 ;
        RECT 1579.710 46.000 2631.590 46.140 ;
        RECT 1579.710 45.940 1580.030 46.000 ;
        RECT 2631.270 45.940 2631.590 46.000 ;
      LAYER via ;
        RECT 1574.220 1311.080 1574.480 1311.340 ;
        RECT 1579.740 1311.080 1580.000 1311.340 ;
        RECT 1579.740 45.940 1580.000 46.200 ;
        RECT 2631.300 45.940 2631.560 46.200 ;
      LAYER met2 ;
        RECT 1574.260 1323.135 1574.540 1327.135 ;
        RECT 1574.280 1311.370 1574.420 1323.135 ;
        RECT 1574.220 1311.050 1574.480 1311.370 ;
        RECT 1579.740 1311.050 1580.000 1311.370 ;
        RECT 1579.800 46.230 1579.940 1311.050 ;
        RECT 1579.740 45.910 1580.000 46.230 ;
        RECT 2631.300 45.910 2631.560 46.230 ;
        RECT 2631.360 2.400 2631.500 45.910 ;
        RECT 2631.150 -4.800 2631.710 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1634.450 46.480 1634.770 46.540 ;
        RECT 2649.210 46.480 2649.530 46.540 ;
        RECT 1634.450 46.340 2649.530 46.480 ;
        RECT 1634.450 46.280 1634.770 46.340 ;
        RECT 2649.210 46.280 2649.530 46.340 ;
      LAYER via ;
        RECT 1634.480 46.280 1634.740 46.540 ;
        RECT 2649.240 46.280 2649.500 46.540 ;
      LAYER met2 ;
        RECT 1632.220 1323.690 1632.500 1327.135 ;
        RECT 1632.220 1323.550 1634.680 1323.690 ;
        RECT 1632.220 1323.135 1632.500 1323.550 ;
        RECT 1634.540 46.570 1634.680 1323.550 ;
        RECT 1634.480 46.250 1634.740 46.570 ;
        RECT 2649.240 46.250 2649.500 46.570 ;
        RECT 2649.300 2.400 2649.440 46.250 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2663.545 2311.745 2663.715 2359.855 ;
        RECT 2663.545 2214.845 2663.715 2262.615 ;
        RECT 2663.545 2118.285 2663.715 2166.395 ;
        RECT 2663.545 2021.725 2663.715 2069.835 ;
        RECT 2663.545 1925.165 2663.715 1973.275 ;
        RECT 2663.545 1828.605 2663.715 1876.715 ;
        RECT 2663.545 1732.045 2663.715 1780.155 ;
        RECT 2663.545 1635.485 2663.715 1683.595 ;
        RECT 2663.545 1538.925 2663.715 1587.035 ;
        RECT 2663.545 1442.025 2663.715 1490.475 ;
        RECT 2663.545 862.665 2663.715 910.435 ;
        RECT 2663.545 766.105 2663.715 814.215 ;
        RECT 2663.545 669.545 2663.715 717.655 ;
        RECT 2663.545 572.645 2663.715 620.415 ;
        RECT 2663.545 476.085 2663.715 524.195 ;
        RECT 2663.545 379.525 2663.715 427.635 ;
        RECT 2663.545 282.965 2663.715 331.075 ;
        RECT 2663.545 186.405 2663.715 234.515 ;
        RECT 2663.545 89.845 2663.715 137.955 ;
      LAYER mcon ;
        RECT 2663.545 2359.685 2663.715 2359.855 ;
        RECT 2663.545 2262.445 2663.715 2262.615 ;
        RECT 2663.545 2166.225 2663.715 2166.395 ;
        RECT 2663.545 2069.665 2663.715 2069.835 ;
        RECT 2663.545 1973.105 2663.715 1973.275 ;
        RECT 2663.545 1876.545 2663.715 1876.715 ;
        RECT 2663.545 1779.985 2663.715 1780.155 ;
        RECT 2663.545 1683.425 2663.715 1683.595 ;
        RECT 2663.545 1586.865 2663.715 1587.035 ;
        RECT 2663.545 1490.305 2663.715 1490.475 ;
        RECT 2663.545 910.265 2663.715 910.435 ;
        RECT 2663.545 814.045 2663.715 814.215 ;
        RECT 2663.545 717.485 2663.715 717.655 ;
        RECT 2663.545 620.245 2663.715 620.415 ;
        RECT 2663.545 524.025 2663.715 524.195 ;
        RECT 2663.545 427.465 2663.715 427.635 ;
        RECT 2663.545 330.905 2663.715 331.075 ;
        RECT 2663.545 234.345 2663.715 234.515 ;
        RECT 2663.545 137.785 2663.715 137.955 ;
      LAYER met1 ;
        RECT 2663.470 2359.840 2663.790 2359.900 ;
        RECT 2663.275 2359.700 2663.790 2359.840 ;
        RECT 2663.470 2359.640 2663.790 2359.700 ;
        RECT 2663.470 2311.900 2663.790 2311.960 ;
        RECT 2663.275 2311.760 2663.790 2311.900 ;
        RECT 2663.470 2311.700 2663.790 2311.760 ;
        RECT 2663.470 2262.600 2663.790 2262.660 ;
        RECT 2663.275 2262.460 2663.790 2262.600 ;
        RECT 2663.470 2262.400 2663.790 2262.460 ;
        RECT 2663.470 2215.000 2663.790 2215.060 ;
        RECT 2663.275 2214.860 2663.790 2215.000 ;
        RECT 2663.470 2214.800 2663.790 2214.860 ;
        RECT 2663.470 2166.380 2663.790 2166.440 ;
        RECT 2663.275 2166.240 2663.790 2166.380 ;
        RECT 2663.470 2166.180 2663.790 2166.240 ;
        RECT 2663.470 2118.440 2663.790 2118.500 ;
        RECT 2663.275 2118.300 2663.790 2118.440 ;
        RECT 2663.470 2118.240 2663.790 2118.300 ;
        RECT 2663.470 2069.820 2663.790 2069.880 ;
        RECT 2663.275 2069.680 2663.790 2069.820 ;
        RECT 2663.470 2069.620 2663.790 2069.680 ;
        RECT 2663.470 2021.880 2663.790 2021.940 ;
        RECT 2663.275 2021.740 2663.790 2021.880 ;
        RECT 2663.470 2021.680 2663.790 2021.740 ;
        RECT 2663.470 1973.260 2663.790 1973.320 ;
        RECT 2663.275 1973.120 2663.790 1973.260 ;
        RECT 2663.470 1973.060 2663.790 1973.120 ;
        RECT 2663.470 1925.320 2663.790 1925.380 ;
        RECT 2663.275 1925.180 2663.790 1925.320 ;
        RECT 2663.470 1925.120 2663.790 1925.180 ;
        RECT 2663.470 1876.700 2663.790 1876.760 ;
        RECT 2663.275 1876.560 2663.790 1876.700 ;
        RECT 2663.470 1876.500 2663.790 1876.560 ;
        RECT 2663.470 1828.760 2663.790 1828.820 ;
        RECT 2663.275 1828.620 2663.790 1828.760 ;
        RECT 2663.470 1828.560 2663.790 1828.620 ;
        RECT 2663.470 1780.140 2663.790 1780.200 ;
        RECT 2663.275 1780.000 2663.790 1780.140 ;
        RECT 2663.470 1779.940 2663.790 1780.000 ;
        RECT 2663.470 1732.200 2663.790 1732.260 ;
        RECT 2663.275 1732.060 2663.790 1732.200 ;
        RECT 2663.470 1732.000 2663.790 1732.060 ;
        RECT 2663.470 1683.580 2663.790 1683.640 ;
        RECT 2663.275 1683.440 2663.790 1683.580 ;
        RECT 2663.470 1683.380 2663.790 1683.440 ;
        RECT 2663.470 1635.640 2663.790 1635.700 ;
        RECT 2663.275 1635.500 2663.790 1635.640 ;
        RECT 2663.470 1635.440 2663.790 1635.500 ;
        RECT 2663.470 1587.020 2663.790 1587.080 ;
        RECT 2663.275 1586.880 2663.790 1587.020 ;
        RECT 2663.470 1586.820 2663.790 1586.880 ;
        RECT 2663.470 1539.080 2663.790 1539.140 ;
        RECT 2663.275 1538.940 2663.790 1539.080 ;
        RECT 2663.470 1538.880 2663.790 1538.940 ;
        RECT 2663.470 1490.460 2663.790 1490.520 ;
        RECT 2663.275 1490.320 2663.790 1490.460 ;
        RECT 2663.470 1490.260 2663.790 1490.320 ;
        RECT 2663.470 1442.180 2663.790 1442.240 ;
        RECT 2663.275 1442.040 2663.790 1442.180 ;
        RECT 2663.470 1441.980 2663.790 1442.040 ;
        RECT 2663.470 1345.620 2663.790 1345.680 ;
        RECT 2664.390 1345.620 2664.710 1345.680 ;
        RECT 2663.470 1345.480 2664.710 1345.620 ;
        RECT 2663.470 1345.420 2663.790 1345.480 ;
        RECT 2664.390 1345.420 2664.710 1345.480 ;
        RECT 2663.470 1249.060 2663.790 1249.120 ;
        RECT 2664.390 1249.060 2664.710 1249.120 ;
        RECT 2663.470 1248.920 2664.710 1249.060 ;
        RECT 2663.470 1248.860 2663.790 1248.920 ;
        RECT 2664.390 1248.860 2664.710 1248.920 ;
        RECT 2663.470 1152.500 2663.790 1152.560 ;
        RECT 2664.390 1152.500 2664.710 1152.560 ;
        RECT 2663.470 1152.360 2664.710 1152.500 ;
        RECT 2663.470 1152.300 2663.790 1152.360 ;
        RECT 2664.390 1152.300 2664.710 1152.360 ;
        RECT 2663.470 1007.320 2663.790 1007.380 ;
        RECT 2664.390 1007.320 2664.710 1007.380 ;
        RECT 2663.470 1007.180 2664.710 1007.320 ;
        RECT 2663.470 1007.120 2663.790 1007.180 ;
        RECT 2664.390 1007.120 2664.710 1007.180 ;
        RECT 2663.470 910.420 2663.790 910.480 ;
        RECT 2663.275 910.280 2663.790 910.420 ;
        RECT 2663.470 910.220 2663.790 910.280 ;
        RECT 2663.470 862.820 2663.790 862.880 ;
        RECT 2663.275 862.680 2663.790 862.820 ;
        RECT 2663.470 862.620 2663.790 862.680 ;
        RECT 2663.470 814.200 2663.790 814.260 ;
        RECT 2663.275 814.060 2663.790 814.200 ;
        RECT 2663.470 814.000 2663.790 814.060 ;
        RECT 2663.470 766.260 2663.790 766.320 ;
        RECT 2663.275 766.120 2663.790 766.260 ;
        RECT 2663.470 766.060 2663.790 766.120 ;
        RECT 2663.470 717.640 2663.790 717.700 ;
        RECT 2663.275 717.500 2663.790 717.640 ;
        RECT 2663.470 717.440 2663.790 717.500 ;
        RECT 2663.470 669.700 2663.790 669.760 ;
        RECT 2663.275 669.560 2663.790 669.700 ;
        RECT 2663.470 669.500 2663.790 669.560 ;
        RECT 2663.470 620.400 2663.790 620.460 ;
        RECT 2663.275 620.260 2663.790 620.400 ;
        RECT 2663.470 620.200 2663.790 620.260 ;
        RECT 2663.470 572.800 2663.790 572.860 ;
        RECT 2663.275 572.660 2663.790 572.800 ;
        RECT 2663.470 572.600 2663.790 572.660 ;
        RECT 2663.470 524.180 2663.790 524.240 ;
        RECT 2663.275 524.040 2663.790 524.180 ;
        RECT 2663.470 523.980 2663.790 524.040 ;
        RECT 2663.470 476.240 2663.790 476.300 ;
        RECT 2663.275 476.100 2663.790 476.240 ;
        RECT 2663.470 476.040 2663.790 476.100 ;
        RECT 2663.470 427.620 2663.790 427.680 ;
        RECT 2663.275 427.480 2663.790 427.620 ;
        RECT 2663.470 427.420 2663.790 427.480 ;
        RECT 2663.470 379.680 2663.790 379.740 ;
        RECT 2663.275 379.540 2663.790 379.680 ;
        RECT 2663.470 379.480 2663.790 379.540 ;
        RECT 2663.470 331.060 2663.790 331.120 ;
        RECT 2663.275 330.920 2663.790 331.060 ;
        RECT 2663.470 330.860 2663.790 330.920 ;
        RECT 2663.470 283.120 2663.790 283.180 ;
        RECT 2663.275 282.980 2663.790 283.120 ;
        RECT 2663.470 282.920 2663.790 282.980 ;
        RECT 2663.470 234.500 2663.790 234.560 ;
        RECT 2663.275 234.360 2663.790 234.500 ;
        RECT 2663.470 234.300 2663.790 234.360 ;
        RECT 2663.470 186.560 2663.790 186.620 ;
        RECT 2663.275 186.420 2663.790 186.560 ;
        RECT 2663.470 186.360 2663.790 186.420 ;
        RECT 2663.470 137.940 2663.790 138.000 ;
        RECT 2663.275 137.800 2663.790 137.940 ;
        RECT 2663.470 137.740 2663.790 137.800 ;
        RECT 2663.470 90.000 2663.790 90.060 ;
        RECT 2663.275 89.860 2663.790 90.000 ;
        RECT 2663.470 89.800 2663.790 89.860 ;
        RECT 2663.470 62.260 2663.790 62.520 ;
        RECT 2663.560 61.780 2663.700 62.260 ;
        RECT 2667.150 61.780 2667.470 61.840 ;
        RECT 2663.560 61.640 2667.470 61.780 ;
        RECT 2667.150 61.580 2667.470 61.640 ;
        RECT 2667.150 47.980 2667.470 48.240 ;
        RECT 2667.240 47.560 2667.380 47.980 ;
        RECT 2667.150 47.300 2667.470 47.560 ;
      LAYER via ;
        RECT 2663.500 2359.640 2663.760 2359.900 ;
        RECT 2663.500 2311.700 2663.760 2311.960 ;
        RECT 2663.500 2262.400 2663.760 2262.660 ;
        RECT 2663.500 2214.800 2663.760 2215.060 ;
        RECT 2663.500 2166.180 2663.760 2166.440 ;
        RECT 2663.500 2118.240 2663.760 2118.500 ;
        RECT 2663.500 2069.620 2663.760 2069.880 ;
        RECT 2663.500 2021.680 2663.760 2021.940 ;
        RECT 2663.500 1973.060 2663.760 1973.320 ;
        RECT 2663.500 1925.120 2663.760 1925.380 ;
        RECT 2663.500 1876.500 2663.760 1876.760 ;
        RECT 2663.500 1828.560 2663.760 1828.820 ;
        RECT 2663.500 1779.940 2663.760 1780.200 ;
        RECT 2663.500 1732.000 2663.760 1732.260 ;
        RECT 2663.500 1683.380 2663.760 1683.640 ;
        RECT 2663.500 1635.440 2663.760 1635.700 ;
        RECT 2663.500 1586.820 2663.760 1587.080 ;
        RECT 2663.500 1538.880 2663.760 1539.140 ;
        RECT 2663.500 1490.260 2663.760 1490.520 ;
        RECT 2663.500 1441.980 2663.760 1442.240 ;
        RECT 2663.500 1345.420 2663.760 1345.680 ;
        RECT 2664.420 1345.420 2664.680 1345.680 ;
        RECT 2663.500 1248.860 2663.760 1249.120 ;
        RECT 2664.420 1248.860 2664.680 1249.120 ;
        RECT 2663.500 1152.300 2663.760 1152.560 ;
        RECT 2664.420 1152.300 2664.680 1152.560 ;
        RECT 2663.500 1007.120 2663.760 1007.380 ;
        RECT 2664.420 1007.120 2664.680 1007.380 ;
        RECT 2663.500 910.220 2663.760 910.480 ;
        RECT 2663.500 862.620 2663.760 862.880 ;
        RECT 2663.500 814.000 2663.760 814.260 ;
        RECT 2663.500 766.060 2663.760 766.320 ;
        RECT 2663.500 717.440 2663.760 717.700 ;
        RECT 2663.500 669.500 2663.760 669.760 ;
        RECT 2663.500 620.200 2663.760 620.460 ;
        RECT 2663.500 572.600 2663.760 572.860 ;
        RECT 2663.500 523.980 2663.760 524.240 ;
        RECT 2663.500 476.040 2663.760 476.300 ;
        RECT 2663.500 427.420 2663.760 427.680 ;
        RECT 2663.500 379.480 2663.760 379.740 ;
        RECT 2663.500 330.860 2663.760 331.120 ;
        RECT 2663.500 282.920 2663.760 283.180 ;
        RECT 2663.500 234.300 2663.760 234.560 ;
        RECT 2663.500 186.360 2663.760 186.620 ;
        RECT 2663.500 137.740 2663.760 138.000 ;
        RECT 2663.500 89.800 2663.760 90.060 ;
        RECT 2663.500 62.260 2663.760 62.520 ;
        RECT 2667.180 61.580 2667.440 61.840 ;
        RECT 2667.180 47.980 2667.440 48.240 ;
        RECT 2667.180 47.300 2667.440 47.560 ;
      LAYER met2 ;
        RECT 1068.260 2374.970 1068.540 2377.880 ;
        RECT 1069.130 2374.970 1069.410 2375.085 ;
        RECT 1068.260 2374.830 1069.410 2374.970 ;
        RECT 1068.260 2373.880 1068.540 2374.830 ;
        RECT 1069.130 2374.715 1069.410 2374.830 ;
        RECT 2663.490 2374.715 2663.770 2375.085 ;
        RECT 2663.560 2359.930 2663.700 2374.715 ;
        RECT 2663.500 2359.610 2663.760 2359.930 ;
        RECT 2663.500 2311.670 2663.760 2311.990 ;
        RECT 2663.560 2262.690 2663.700 2311.670 ;
        RECT 2663.500 2262.370 2663.760 2262.690 ;
        RECT 2663.500 2214.770 2663.760 2215.090 ;
        RECT 2663.560 2166.470 2663.700 2214.770 ;
        RECT 2663.500 2166.150 2663.760 2166.470 ;
        RECT 2663.500 2118.210 2663.760 2118.530 ;
        RECT 2663.560 2069.910 2663.700 2118.210 ;
        RECT 2663.500 2069.590 2663.760 2069.910 ;
        RECT 2663.500 2021.650 2663.760 2021.970 ;
        RECT 2663.560 1973.350 2663.700 2021.650 ;
        RECT 2663.500 1973.030 2663.760 1973.350 ;
        RECT 2663.500 1925.090 2663.760 1925.410 ;
        RECT 2663.560 1876.790 2663.700 1925.090 ;
        RECT 2663.500 1876.470 2663.760 1876.790 ;
        RECT 2663.500 1828.530 2663.760 1828.850 ;
        RECT 2663.560 1780.230 2663.700 1828.530 ;
        RECT 2663.500 1779.910 2663.760 1780.230 ;
        RECT 2663.500 1731.970 2663.760 1732.290 ;
        RECT 2663.560 1683.670 2663.700 1731.970 ;
        RECT 2663.500 1683.350 2663.760 1683.670 ;
        RECT 2663.500 1635.410 2663.760 1635.730 ;
        RECT 2663.560 1587.110 2663.700 1635.410 ;
        RECT 2663.500 1586.790 2663.760 1587.110 ;
        RECT 2663.500 1538.850 2663.760 1539.170 ;
        RECT 2663.560 1490.550 2663.700 1538.850 ;
        RECT 2663.500 1490.230 2663.760 1490.550 ;
        RECT 2663.500 1441.950 2663.760 1442.270 ;
        RECT 2663.560 1393.845 2663.700 1441.950 ;
        RECT 2663.490 1393.475 2663.770 1393.845 ;
        RECT 2664.410 1393.475 2664.690 1393.845 ;
        RECT 2664.480 1345.710 2664.620 1393.475 ;
        RECT 2663.500 1345.390 2663.760 1345.710 ;
        RECT 2664.420 1345.390 2664.680 1345.710 ;
        RECT 2663.560 1297.285 2663.700 1345.390 ;
        RECT 2663.490 1296.915 2663.770 1297.285 ;
        RECT 2664.410 1296.915 2664.690 1297.285 ;
        RECT 2664.480 1249.150 2664.620 1296.915 ;
        RECT 2663.500 1248.830 2663.760 1249.150 ;
        RECT 2664.420 1248.830 2664.680 1249.150 ;
        RECT 2663.560 1200.725 2663.700 1248.830 ;
        RECT 2663.490 1200.355 2663.770 1200.725 ;
        RECT 2664.410 1200.355 2664.690 1200.725 ;
        RECT 2664.480 1152.590 2664.620 1200.355 ;
        RECT 2663.500 1152.270 2663.760 1152.590 ;
        RECT 2664.420 1152.270 2664.680 1152.590 ;
        RECT 2663.560 1104.165 2663.700 1152.270 ;
        RECT 2663.490 1103.795 2663.770 1104.165 ;
        RECT 2664.410 1103.795 2664.690 1104.165 ;
        RECT 2664.480 1055.885 2664.620 1103.795 ;
        RECT 2663.490 1055.515 2663.770 1055.885 ;
        RECT 2664.410 1055.515 2664.690 1055.885 ;
        RECT 2663.560 1007.410 2663.700 1055.515 ;
        RECT 2663.500 1007.090 2663.760 1007.410 ;
        RECT 2664.420 1007.090 2664.680 1007.410 ;
        RECT 2664.480 959.325 2664.620 1007.090 ;
        RECT 2663.490 958.955 2663.770 959.325 ;
        RECT 2664.410 958.955 2664.690 959.325 ;
        RECT 2663.560 910.510 2663.700 958.955 ;
        RECT 2663.500 910.190 2663.760 910.510 ;
        RECT 2663.500 862.590 2663.760 862.910 ;
        RECT 2663.560 814.290 2663.700 862.590 ;
        RECT 2663.500 813.970 2663.760 814.290 ;
        RECT 2663.500 766.030 2663.760 766.350 ;
        RECT 2663.560 717.730 2663.700 766.030 ;
        RECT 2663.500 717.410 2663.760 717.730 ;
        RECT 2663.500 669.470 2663.760 669.790 ;
        RECT 2663.560 620.490 2663.700 669.470 ;
        RECT 2663.500 620.170 2663.760 620.490 ;
        RECT 2663.500 572.570 2663.760 572.890 ;
        RECT 2663.560 524.270 2663.700 572.570 ;
        RECT 2663.500 523.950 2663.760 524.270 ;
        RECT 2663.500 476.010 2663.760 476.330 ;
        RECT 2663.560 427.710 2663.700 476.010 ;
        RECT 2663.500 427.390 2663.760 427.710 ;
        RECT 2663.500 379.450 2663.760 379.770 ;
        RECT 2663.560 331.150 2663.700 379.450 ;
        RECT 2663.500 330.830 2663.760 331.150 ;
        RECT 2663.500 282.890 2663.760 283.210 ;
        RECT 2663.560 234.590 2663.700 282.890 ;
        RECT 2663.500 234.270 2663.760 234.590 ;
        RECT 2663.500 186.330 2663.760 186.650 ;
        RECT 2663.560 138.030 2663.700 186.330 ;
        RECT 2663.500 137.710 2663.760 138.030 ;
        RECT 2663.500 89.770 2663.760 90.090 ;
        RECT 2663.560 62.550 2663.700 89.770 ;
        RECT 2663.500 62.230 2663.760 62.550 ;
        RECT 2667.180 61.550 2667.440 61.870 ;
        RECT 2667.240 48.270 2667.380 61.550 ;
        RECT 2667.180 47.950 2667.440 48.270 ;
        RECT 2667.180 47.270 2667.440 47.590 ;
        RECT 2667.240 2.400 2667.380 47.270 ;
        RECT 2667.030 -4.800 2667.590 2.400 ;
      LAYER via2 ;
        RECT 1069.130 2374.760 1069.410 2375.040 ;
        RECT 2663.490 2374.760 2663.770 2375.040 ;
        RECT 2663.490 1393.520 2663.770 1393.800 ;
        RECT 2664.410 1393.520 2664.690 1393.800 ;
        RECT 2663.490 1296.960 2663.770 1297.240 ;
        RECT 2664.410 1296.960 2664.690 1297.240 ;
        RECT 2663.490 1200.400 2663.770 1200.680 ;
        RECT 2664.410 1200.400 2664.690 1200.680 ;
        RECT 2663.490 1103.840 2663.770 1104.120 ;
        RECT 2664.410 1103.840 2664.690 1104.120 ;
        RECT 2663.490 1055.560 2663.770 1055.840 ;
        RECT 2664.410 1055.560 2664.690 1055.840 ;
        RECT 2663.490 959.000 2663.770 959.280 ;
        RECT 2664.410 959.000 2664.690 959.280 ;
      LAYER met3 ;
        RECT 1069.105 2375.050 1069.435 2375.065 ;
        RECT 2663.465 2375.050 2663.795 2375.065 ;
        RECT 1069.105 2374.750 2663.795 2375.050 ;
        RECT 1069.105 2374.735 1069.435 2374.750 ;
        RECT 2663.465 2374.735 2663.795 2374.750 ;
        RECT 2663.465 1393.810 2663.795 1393.825 ;
        RECT 2664.385 1393.810 2664.715 1393.825 ;
        RECT 2663.465 1393.510 2664.715 1393.810 ;
        RECT 2663.465 1393.495 2663.795 1393.510 ;
        RECT 2664.385 1393.495 2664.715 1393.510 ;
        RECT 2663.465 1297.250 2663.795 1297.265 ;
        RECT 2664.385 1297.250 2664.715 1297.265 ;
        RECT 2663.465 1296.950 2664.715 1297.250 ;
        RECT 2663.465 1296.935 2663.795 1296.950 ;
        RECT 2664.385 1296.935 2664.715 1296.950 ;
        RECT 2663.465 1200.690 2663.795 1200.705 ;
        RECT 2664.385 1200.690 2664.715 1200.705 ;
        RECT 2663.465 1200.390 2664.715 1200.690 ;
        RECT 2663.465 1200.375 2663.795 1200.390 ;
        RECT 2664.385 1200.375 2664.715 1200.390 ;
        RECT 2663.465 1104.130 2663.795 1104.145 ;
        RECT 2664.385 1104.130 2664.715 1104.145 ;
        RECT 2663.465 1103.830 2664.715 1104.130 ;
        RECT 2663.465 1103.815 2663.795 1103.830 ;
        RECT 2664.385 1103.815 2664.715 1103.830 ;
        RECT 2663.465 1055.850 2663.795 1055.865 ;
        RECT 2664.385 1055.850 2664.715 1055.865 ;
        RECT 2663.465 1055.550 2664.715 1055.850 ;
        RECT 2663.465 1055.535 2663.795 1055.550 ;
        RECT 2664.385 1055.535 2664.715 1055.550 ;
        RECT 2663.465 959.290 2663.795 959.305 ;
        RECT 2664.385 959.290 2664.715 959.305 ;
        RECT 2663.465 958.990 2664.715 959.290 ;
        RECT 2663.465 958.975 2663.795 958.990 ;
        RECT 2664.385 958.975 2664.715 958.990 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2684.650 15.115 2684.930 15.485 ;
        RECT 2684.720 2.400 2684.860 15.115 ;
        RECT 2684.510 -4.800 2685.070 2.400 ;
      LAYER via2 ;
        RECT 2684.650 15.160 2684.930 15.440 ;
      LAYER met3 ;
        RECT 712.350 1695.050 712.730 1695.060 ;
        RECT 715.810 1695.050 719.810 1695.055 ;
        RECT 712.350 1694.750 719.810 1695.050 ;
        RECT 712.350 1694.740 712.730 1694.750 ;
        RECT 715.810 1694.455 719.810 1694.750 ;
        RECT 958.910 25.650 959.290 25.660 ;
        RECT 969.030 25.650 969.410 25.660 ;
        RECT 958.910 25.350 969.410 25.650 ;
        RECT 958.910 25.340 959.290 25.350 ;
        RECT 969.030 25.340 969.410 25.350 ;
        RECT 2412.510 25.650 2412.890 25.660 ;
        RECT 2418.030 25.650 2418.410 25.660 ;
        RECT 2412.510 25.350 2418.410 25.650 ;
        RECT 2412.510 25.340 2412.890 25.350 ;
        RECT 2418.030 25.340 2418.410 25.350 ;
        RECT 1007.670 22.250 1008.050 22.260 ;
        RECT 1054.590 22.250 1054.970 22.260 ;
        RECT 1007.670 21.950 1054.970 22.250 ;
        RECT 1007.670 21.940 1008.050 21.950 ;
        RECT 1054.590 21.940 1054.970 21.950 ;
        RECT 1628.670 22.250 1629.050 22.260 ;
        RECT 1659.950 22.250 1660.330 22.260 ;
        RECT 1628.670 21.950 1660.330 22.250 ;
        RECT 1628.670 21.940 1629.050 21.950 ;
        RECT 1659.950 21.940 1660.330 21.950 ;
        RECT 1766.670 22.250 1767.050 22.260 ;
        RECT 1813.590 22.250 1813.970 22.260 ;
        RECT 1766.670 21.950 1813.970 22.250 ;
        RECT 1766.670 21.940 1767.050 21.950 ;
        RECT 1813.590 21.940 1813.970 21.950 ;
        RECT 1997.590 22.250 1997.970 22.260 ;
        RECT 2027.950 22.250 2028.330 22.260 ;
        RECT 1997.590 21.950 2028.330 22.250 ;
        RECT 1997.590 21.940 1997.970 21.950 ;
        RECT 2027.950 21.940 2028.330 21.950 ;
        RECT 2200.910 22.250 2201.290 22.260 ;
        RECT 2248.750 22.250 2249.130 22.260 ;
        RECT 2200.910 21.950 2249.130 22.250 ;
        RECT 2200.910 21.940 2201.290 21.950 ;
        RECT 2248.750 21.940 2249.130 21.950 ;
        RECT 2360.990 22.250 2361.370 22.260 ;
        RECT 2369.270 22.250 2369.650 22.260 ;
        RECT 2360.990 21.950 2369.650 22.250 ;
        RECT 2360.990 21.940 2361.370 21.950 ;
        RECT 2369.270 21.940 2369.650 21.950 ;
        RECT 2456.670 22.250 2457.050 22.260 ;
        RECT 2503.590 22.250 2503.970 22.260 ;
        RECT 2456.670 21.950 2503.970 22.250 ;
        RECT 2456.670 21.940 2457.050 21.950 ;
        RECT 2503.590 21.940 2503.970 21.950 ;
        RECT 1690.310 21.570 1690.690 21.580 ;
        RECT 1753.790 21.570 1754.170 21.580 ;
        RECT 1690.310 21.270 1754.170 21.570 ;
        RECT 1690.310 21.260 1690.690 21.270 ;
        RECT 1753.790 21.260 1754.170 21.270 ;
        RECT 862.310 20.890 862.690 20.900 ;
        RECT 910.150 20.890 910.530 20.900 ;
        RECT 862.310 20.590 910.530 20.890 ;
        RECT 862.310 20.580 862.690 20.590 ;
        RECT 910.150 20.580 910.530 20.590 ;
        RECT 773.070 20.210 773.450 20.220 ;
        RECT 786.870 20.210 787.250 20.220 ;
        RECT 773.070 19.910 787.250 20.210 ;
        RECT 773.070 19.900 773.450 19.910 ;
        RECT 786.870 19.900 787.250 19.910 ;
        RECT 2570.750 15.450 2571.130 15.460 ;
        RECT 2648.950 15.450 2649.330 15.460 ;
        RECT 2570.750 15.150 2649.330 15.450 ;
        RECT 2570.750 15.140 2571.130 15.150 ;
        RECT 2648.950 15.140 2649.330 15.150 ;
        RECT 2660.910 15.450 2661.290 15.460 ;
        RECT 2684.625 15.450 2684.955 15.465 ;
        RECT 2660.910 15.150 2684.955 15.450 ;
        RECT 2660.910 15.140 2661.290 15.150 ;
        RECT 2684.625 15.135 2684.955 15.150 ;
        RECT 820.910 14.090 821.290 14.100 ;
        RECT 837.470 14.090 837.850 14.100 ;
        RECT 820.910 13.790 837.850 14.090 ;
        RECT 820.910 13.780 821.290 13.790 ;
        RECT 837.470 13.780 837.850 13.790 ;
      LAYER via3 ;
        RECT 712.380 1694.740 712.700 1695.060 ;
        RECT 958.940 25.340 959.260 25.660 ;
        RECT 969.060 25.340 969.380 25.660 ;
        RECT 2412.540 25.340 2412.860 25.660 ;
        RECT 2418.060 25.340 2418.380 25.660 ;
        RECT 1007.700 21.940 1008.020 22.260 ;
        RECT 1054.620 21.940 1054.940 22.260 ;
        RECT 1628.700 21.940 1629.020 22.260 ;
        RECT 1659.980 21.940 1660.300 22.260 ;
        RECT 1766.700 21.940 1767.020 22.260 ;
        RECT 1813.620 21.940 1813.940 22.260 ;
        RECT 1997.620 21.940 1997.940 22.260 ;
        RECT 2027.980 21.940 2028.300 22.260 ;
        RECT 2200.940 21.940 2201.260 22.260 ;
        RECT 2248.780 21.940 2249.100 22.260 ;
        RECT 2361.020 21.940 2361.340 22.260 ;
        RECT 2369.300 21.940 2369.620 22.260 ;
        RECT 2456.700 21.940 2457.020 22.260 ;
        RECT 2503.620 21.940 2503.940 22.260 ;
        RECT 1690.340 21.260 1690.660 21.580 ;
        RECT 1753.820 21.260 1754.140 21.580 ;
        RECT 862.340 20.580 862.660 20.900 ;
        RECT 910.180 20.580 910.500 20.900 ;
        RECT 773.100 19.900 773.420 20.220 ;
        RECT 786.900 19.900 787.220 20.220 ;
        RECT 2570.780 15.140 2571.100 15.460 ;
        RECT 2648.980 15.140 2649.300 15.460 ;
        RECT 2660.940 15.140 2661.260 15.460 ;
        RECT 820.940 13.780 821.260 14.100 ;
        RECT 837.500 13.780 837.820 14.100 ;
      LAYER met4 ;
        RECT 712.375 1694.735 712.705 1695.065 ;
        RECT 712.390 19.290 712.690 1694.735 ;
        RECT 958.510 24.910 959.690 26.090 ;
        RECT 969.055 25.335 969.385 25.665 ;
        RECT 969.070 22.690 969.370 25.335 ;
        RECT 2368.870 24.910 2370.050 26.090 ;
        RECT 2412.110 24.910 2413.290 26.090 ;
        RECT 2418.055 25.335 2418.385 25.665 ;
        RECT 968.630 21.510 969.810 22.690 ;
        RECT 1007.270 21.510 1008.450 22.690 ;
        RECT 1054.190 21.510 1055.370 22.690 ;
        RECT 1628.270 21.510 1629.450 22.690 ;
        RECT 1659.975 21.935 1660.305 22.265 ;
        RECT 862.335 20.575 862.665 20.905 ;
        RECT 910.175 20.575 910.505 20.905 ;
        RECT 773.095 19.895 773.425 20.225 ;
        RECT 786.895 19.895 787.225 20.225 ;
        RECT 773.110 19.290 773.410 19.895 ;
        RECT 711.950 18.110 713.130 19.290 ;
        RECT 772.670 18.110 773.850 19.290 ;
        RECT 786.910 15.890 787.210 19.895 ;
        RECT 862.350 19.290 862.650 20.575 ;
        RECT 910.190 19.290 910.490 20.575 ;
        RECT 1659.990 19.290 1660.290 21.935 ;
        RECT 1690.335 21.255 1690.665 21.585 ;
        RECT 1753.390 21.510 1754.570 22.690 ;
        RECT 1766.270 21.510 1767.450 22.690 ;
        RECT 1813.190 21.510 1814.370 22.690 ;
        RECT 1997.190 21.510 1998.370 22.690 ;
        RECT 2027.975 21.935 2028.305 22.265 ;
        RECT 1753.815 21.255 1754.145 21.510 ;
        RECT 1690.350 19.290 1690.650 21.255 ;
        RECT 2027.990 19.290 2028.290 21.935 ;
        RECT 2200.510 21.510 2201.690 22.690 ;
        RECT 2248.775 21.935 2249.105 22.265 ;
        RECT 2248.790 19.290 2249.090 21.935 ;
        RECT 2307.230 21.510 2308.410 22.690 ;
        RECT 2360.590 21.510 2361.770 22.690 ;
        RECT 2369.310 22.265 2369.610 24.910 ;
        RECT 2418.070 22.690 2418.370 25.335 ;
        RECT 2369.295 21.935 2369.625 22.265 ;
        RECT 2417.630 21.510 2418.810 22.690 ;
        RECT 2456.270 21.510 2457.450 22.690 ;
        RECT 2503.615 21.935 2503.945 22.265 ;
        RECT 837.070 18.110 838.250 19.290 ;
        RECT 861.910 18.110 863.090 19.290 ;
        RECT 909.750 18.110 910.930 19.290 ;
        RECT 1659.550 18.110 1660.730 19.290 ;
        RECT 1689.910 18.110 1691.090 19.290 ;
        RECT 2027.550 18.110 2028.730 19.290 ;
        RECT 2248.350 18.110 2249.530 19.290 ;
        RECT 2305.390 18.850 2306.570 19.290 ;
        RECT 2307.670 18.850 2307.970 21.510 ;
        RECT 2305.390 18.550 2307.970 18.850 ;
        RECT 2305.390 18.110 2306.570 18.550 ;
        RECT 786.470 14.710 787.650 15.890 ;
        RECT 820.510 14.710 821.690 15.890 ;
        RECT 820.950 14.105 821.250 14.710 ;
        RECT 837.510 14.105 837.810 18.110 ;
        RECT 820.935 13.775 821.265 14.105 ;
        RECT 837.495 13.775 837.825 14.105 ;
        RECT 2503.630 12.490 2503.930 21.935 ;
        RECT 2648.550 21.510 2649.730 22.690 ;
        RECT 2570.350 14.710 2571.530 15.890 ;
        RECT 2648.990 15.465 2649.290 21.510 ;
        RECT 2648.975 15.135 2649.305 15.465 ;
        RECT 2660.510 14.710 2661.690 15.890 ;
        RECT 2503.190 11.310 2504.370 12.490 ;
      LAYER via4 ;
        RECT 1753.390 21.510 1754.570 22.690 ;
      LAYER met5 ;
        RECT 916.900 24.700 959.900 26.300 ;
        RECT 1812.980 24.700 1853.220 26.300 ;
        RECT 916.900 19.500 918.500 24.700 ;
        RECT 968.420 21.300 1008.660 22.900 ;
        RECT 1053.980 21.300 1080.420 22.900 ;
        RECT 711.740 17.900 774.060 19.500 ;
        RECT 836.860 17.900 863.300 19.500 ;
        RECT 909.540 17.900 918.500 19.500 ;
        RECT 1078.820 19.500 1080.420 21.300 ;
        RECT 1121.140 21.300 1629.660 22.900 ;
        RECT 1753.180 21.300 1767.660 22.900 ;
        RECT 1812.980 21.300 1814.580 24.700 ;
        RECT 1851.620 22.900 1853.220 24.700 ;
        RECT 2064.140 24.700 2109.900 26.300 ;
        RECT 2368.660 24.700 2413.500 26.300 ;
        RECT 1851.620 21.300 1998.580 22.900 ;
        RECT 1121.140 19.500 1122.740 21.300 ;
        RECT 2064.140 19.500 2065.740 24.700 ;
        RECT 1078.820 17.900 1122.740 19.500 ;
        RECT 1659.340 17.900 1691.300 19.500 ;
        RECT 2027.340 17.900 2065.740 19.500 ;
        RECT 2108.300 19.500 2109.900 24.700 ;
        RECT 2200.300 19.500 2201.900 22.900 ;
        RECT 2307.020 21.300 2361.980 22.900 ;
        RECT 2417.420 21.300 2457.660 22.900 ;
        RECT 2648.340 21.300 2656.380 22.900 ;
        RECT 2108.300 17.900 2201.900 19.500 ;
        RECT 2248.140 17.900 2306.780 19.500 ;
        RECT 2654.780 16.100 2656.380 21.300 ;
        RECT 786.260 14.500 821.900 16.100 ;
        RECT 2527.820 14.500 2571.740 16.100 ;
        RECT 2654.780 14.500 2661.900 16.100 ;
        RECT 2527.820 12.700 2529.420 14.500 ;
        RECT 2502.980 11.100 2529.420 12.700 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 882.810 45.460 883.130 45.520 ;
        RECT 2702.570 45.460 2702.890 45.520 ;
        RECT 882.810 45.320 2702.890 45.460 ;
        RECT 882.810 45.260 883.130 45.320 ;
        RECT 2702.570 45.260 2702.890 45.320 ;
      LAYER via ;
        RECT 882.840 45.260 883.100 45.520 ;
        RECT 2702.600 45.260 2702.860 45.520 ;
      LAYER met2 ;
        RECT 880.580 1323.690 880.860 1327.135 ;
        RECT 880.580 1323.550 883.040 1323.690 ;
        RECT 880.580 1323.135 880.860 1323.550 ;
        RECT 882.900 45.550 883.040 1323.550 ;
        RECT 882.840 45.230 883.100 45.550 ;
        RECT 2702.600 45.230 2702.860 45.550 ;
        RECT 2702.660 2.400 2702.800 45.230 ;
        RECT 2702.450 -4.800 2703.010 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1486.330 2374.460 1486.650 2374.520 ;
        RECT 2718.670 2374.460 2718.990 2374.520 ;
        RECT 1486.330 2374.320 2718.990 2374.460 ;
        RECT 1486.330 2374.260 1486.650 2374.320 ;
        RECT 2718.670 2374.260 2718.990 2374.320 ;
        RECT 2718.670 2.960 2718.990 3.020 ;
        RECT 2720.510 2.960 2720.830 3.020 ;
        RECT 2718.670 2.820 2720.830 2.960 ;
        RECT 2718.670 2.760 2718.990 2.820 ;
        RECT 2720.510 2.760 2720.830 2.820 ;
      LAYER via ;
        RECT 1486.360 2374.260 1486.620 2374.520 ;
        RECT 2718.700 2374.260 2718.960 2374.520 ;
        RECT 2718.700 2.760 2718.960 3.020 ;
        RECT 2720.540 2.760 2720.800 3.020 ;
      LAYER met2 ;
        RECT 1485.020 2374.290 1485.300 2377.880 ;
        RECT 1486.360 2374.290 1486.620 2374.550 ;
        RECT 1485.020 2374.230 1486.620 2374.290 ;
        RECT 2718.700 2374.230 2718.960 2374.550 ;
        RECT 1485.020 2374.150 1486.560 2374.230 ;
        RECT 1485.020 2373.880 1485.300 2374.150 ;
        RECT 2718.760 3.050 2718.900 2374.230 ;
        RECT 2718.700 2.730 2718.960 3.050 ;
        RECT 2720.540 2.730 2720.800 3.050 ;
        RECT 2720.600 2.400 2720.740 2.730 ;
        RECT 2720.390 -4.800 2720.950 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1379.150 1255.660 1379.470 1255.920 ;
        RECT 1379.240 1255.240 1379.380 1255.660 ;
        RECT 1379.150 1254.980 1379.470 1255.240 ;
        RECT 1379.150 45.800 1379.470 45.860 ;
        RECT 2738.450 45.800 2738.770 45.860 ;
        RECT 1379.150 45.660 2738.770 45.800 ;
        RECT 1379.150 45.600 1379.470 45.660 ;
        RECT 2738.450 45.600 2738.770 45.660 ;
      LAYER via ;
        RECT 1379.180 1255.660 1379.440 1255.920 ;
        RECT 1379.180 1254.980 1379.440 1255.240 ;
        RECT 1379.180 45.600 1379.440 45.860 ;
        RECT 2738.480 45.600 2738.740 45.860 ;
      LAYER met2 ;
        RECT 1377.380 1323.690 1377.660 1327.135 ;
        RECT 1377.380 1323.550 1379.380 1323.690 ;
        RECT 1377.380 1323.135 1377.660 1323.550 ;
        RECT 1379.240 1255.950 1379.380 1323.550 ;
        RECT 1379.180 1255.630 1379.440 1255.950 ;
        RECT 1379.180 1254.950 1379.440 1255.270 ;
        RECT 1379.240 45.890 1379.380 1254.950 ;
        RECT 1379.180 45.570 1379.440 45.890 ;
        RECT 2738.480 45.570 2738.740 45.890 ;
        RECT 2738.540 2.400 2738.680 45.570 ;
        RECT 2738.330 -4.800 2738.890 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 782.070 1311.620 782.390 1311.680 ;
        RECT 786.210 1311.620 786.530 1311.680 ;
        RECT 782.070 1311.480 786.530 1311.620 ;
        RECT 782.070 1311.420 782.390 1311.480 ;
        RECT 786.210 1311.420 786.530 1311.480 ;
        RECT 786.210 44.780 786.530 44.840 ;
        RECT 2755.930 44.780 2756.250 44.840 ;
        RECT 786.210 44.640 2756.250 44.780 ;
        RECT 786.210 44.580 786.530 44.640 ;
        RECT 2755.930 44.580 2756.250 44.640 ;
      LAYER via ;
        RECT 782.100 1311.420 782.360 1311.680 ;
        RECT 786.240 1311.420 786.500 1311.680 ;
        RECT 786.240 44.580 786.500 44.840 ;
        RECT 2755.960 44.580 2756.220 44.840 ;
      LAYER met2 ;
        RECT 782.140 1323.135 782.420 1327.135 ;
        RECT 782.160 1311.710 782.300 1323.135 ;
        RECT 782.100 1311.390 782.360 1311.710 ;
        RECT 786.240 1311.390 786.500 1311.710 ;
        RECT 786.300 44.870 786.440 1311.390 ;
        RECT 786.240 44.550 786.500 44.870 ;
        RECT 2755.960 44.550 2756.220 44.870 ;
        RECT 2756.020 2.400 2756.160 44.550 ;
        RECT 2755.810 -4.800 2756.370 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 748.030 2374.260 748.350 2374.520 ;
        RECT 696.510 2374.120 696.830 2374.180 ;
        RECT 748.120 2374.120 748.260 2374.260 ;
        RECT 696.510 2373.980 748.260 2374.120 ;
        RECT 696.510 2373.920 696.830 2373.980 ;
        RECT 696.510 15.540 696.830 15.600 ;
        RECT 829.450 15.540 829.770 15.600 ;
        RECT 696.510 15.400 829.770 15.540 ;
        RECT 696.510 15.340 696.830 15.400 ;
        RECT 829.450 15.340 829.770 15.400 ;
      LAYER via ;
        RECT 748.060 2374.260 748.320 2374.520 ;
        RECT 696.540 2373.920 696.800 2374.180 ;
        RECT 696.540 15.340 696.800 15.600 ;
        RECT 829.480 15.340 829.740 15.600 ;
      LAYER met2 ;
        RECT 748.060 2374.290 748.320 2374.550 ;
        RECT 749.940 2374.290 750.220 2377.880 ;
        RECT 748.060 2374.230 750.220 2374.290 ;
        RECT 696.540 2373.890 696.800 2374.210 ;
        RECT 748.120 2374.150 750.220 2374.230 ;
        RECT 696.600 1393.845 696.740 2373.890 ;
        RECT 749.940 2373.880 750.220 2374.150 ;
        RECT 696.530 1393.475 696.810 1393.845 ;
        RECT 696.530 1392.115 696.810 1392.485 ;
        RECT 696.600 15.630 696.740 1392.115 ;
        RECT 696.540 15.310 696.800 15.630 ;
        RECT 829.480 15.310 829.740 15.630 ;
        RECT 829.540 2.400 829.680 15.310 ;
        RECT 829.330 -4.800 829.890 2.400 ;
      LAYER via2 ;
        RECT 696.530 1393.520 696.810 1393.800 ;
        RECT 696.530 1392.160 696.810 1392.440 ;
      LAYER met3 ;
        RECT 696.505 1393.810 696.835 1393.825 ;
        RECT 696.505 1393.495 697.050 1393.810 ;
        RECT 696.750 1392.465 697.050 1393.495 ;
        RECT 696.505 1392.150 697.050 1392.465 ;
        RECT 696.505 1392.135 696.835 1392.150 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 712.150 86.260 712.470 86.320 ;
        RECT 2774.330 86.260 2774.650 86.320 ;
        RECT 712.150 86.120 2774.650 86.260 ;
        RECT 712.150 86.060 712.470 86.120 ;
        RECT 2774.330 86.060 2774.650 86.120 ;
      LAYER via ;
        RECT 712.180 86.060 712.440 86.320 ;
        RECT 2774.360 86.060 2774.620 86.320 ;
      LAYER met2 ;
        RECT 712.170 1583.195 712.450 1583.565 ;
        RECT 712.240 86.350 712.380 1583.195 ;
        RECT 712.180 86.030 712.440 86.350 ;
        RECT 2774.360 86.030 2774.620 86.350 ;
        RECT 2774.420 17.410 2774.560 86.030 ;
        RECT 2773.960 17.270 2774.560 17.410 ;
        RECT 2773.960 2.400 2774.100 17.270 ;
        RECT 2773.750 -4.800 2774.310 2.400 ;
      LAYER via2 ;
        RECT 712.170 1583.240 712.450 1583.520 ;
      LAYER met3 ;
        RECT 712.145 1583.530 712.475 1583.545 ;
        RECT 715.810 1583.530 719.810 1583.535 ;
        RECT 712.145 1583.230 719.810 1583.530 ;
        RECT 712.145 1583.215 712.475 1583.230 ;
        RECT 715.810 1582.935 719.810 1583.230 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 712.610 1500.660 712.930 1500.720 ;
        RECT 716.750 1500.660 717.070 1500.720 ;
        RECT 712.610 1500.520 717.070 1500.660 ;
        RECT 712.610 1500.460 712.930 1500.520 ;
        RECT 716.750 1500.460 717.070 1500.520 ;
      LAYER via ;
        RECT 712.640 1500.460 712.900 1500.720 ;
        RECT 716.780 1500.460 717.040 1500.720 ;
      LAYER met2 ;
        RECT 716.770 2196.555 717.050 2196.925 ;
        RECT 716.840 1500.750 716.980 2196.555 ;
        RECT 712.640 1500.430 712.900 1500.750 ;
        RECT 716.780 1500.430 717.040 1500.750 ;
        RECT 712.700 1452.325 712.840 1500.430 ;
        RECT 712.630 1451.955 712.910 1452.325 ;
        RECT 716.310 1328.875 716.590 1329.245 ;
        RECT 716.380 1293.885 716.520 1328.875 ;
        RECT 716.310 1293.515 716.590 1293.885 ;
        RECT 2787.690 1293.515 2787.970 1293.885 ;
        RECT 2787.760 17.410 2787.900 1293.515 ;
        RECT 2787.760 17.270 2792.040 17.410 ;
        RECT 2791.900 2.400 2792.040 17.270 ;
        RECT 2791.690 -4.800 2792.250 2.400 ;
      LAYER via2 ;
        RECT 716.770 2196.600 717.050 2196.880 ;
        RECT 712.630 1452.000 712.910 1452.280 ;
        RECT 716.310 1328.920 716.590 1329.200 ;
        RECT 716.310 1293.560 716.590 1293.840 ;
        RECT 2787.690 1293.560 2787.970 1293.840 ;
      LAYER met3 ;
        RECT 715.810 2199.015 719.810 2199.615 ;
        RECT 716.990 2196.905 717.290 2199.015 ;
        RECT 716.745 2196.590 717.290 2196.905 ;
        RECT 716.745 2196.575 717.075 2196.590 ;
        RECT 712.605 1452.290 712.935 1452.305 ;
        RECT 716.030 1452.290 716.410 1452.300 ;
        RECT 712.605 1451.990 716.410 1452.290 ;
        RECT 712.605 1451.975 712.935 1451.990 ;
        RECT 716.030 1451.980 716.410 1451.990 ;
        RECT 716.030 1426.820 716.410 1427.140 ;
        RECT 716.070 1425.780 716.370 1426.820 ;
        RECT 716.030 1425.460 716.410 1425.780 ;
        RECT 716.285 1329.220 716.615 1329.225 ;
        RECT 716.030 1329.210 716.615 1329.220 ;
        RECT 715.830 1328.910 716.615 1329.210 ;
        RECT 716.030 1328.900 716.615 1328.910 ;
        RECT 716.285 1328.895 716.615 1328.900 ;
        RECT 716.285 1293.850 716.615 1293.865 ;
        RECT 2787.665 1293.850 2787.995 1293.865 ;
        RECT 716.285 1293.550 2787.995 1293.850 ;
        RECT 716.285 1293.535 716.615 1293.550 ;
        RECT 2787.665 1293.535 2787.995 1293.550 ;
      LAYER via3 ;
        RECT 716.060 1451.980 716.380 1452.300 ;
        RECT 716.060 1426.820 716.380 1427.140 ;
        RECT 716.060 1425.460 716.380 1425.780 ;
        RECT 716.060 1328.900 716.380 1329.220 ;
      LAYER met4 ;
        RECT 716.055 1451.975 716.385 1452.305 ;
        RECT 716.070 1427.145 716.370 1451.975 ;
        RECT 716.055 1426.815 716.385 1427.145 ;
        RECT 716.055 1425.455 716.385 1425.785 ;
        RECT 716.070 1329.225 716.370 1425.455 ;
        RECT 716.055 1328.895 716.385 1329.225 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2808.390 85.835 2808.670 86.205 ;
        RECT 2808.460 17.410 2808.600 85.835 ;
        RECT 2808.460 17.270 2809.980 17.410 ;
        RECT 2809.840 2.400 2809.980 17.270 ;
        RECT 2809.630 -4.800 2810.190 2.400 ;
      LAYER via2 ;
        RECT 2808.390 85.880 2808.670 86.160 ;
      LAYER met3 ;
        RECT 711.430 2156.090 711.810 2156.100 ;
        RECT 715.810 2156.090 719.810 2156.095 ;
        RECT 711.430 2155.790 719.810 2156.090 ;
        RECT 711.430 2155.780 711.810 2155.790 ;
        RECT 715.810 2155.495 719.810 2155.790 ;
        RECT 711.430 86.170 711.810 86.180 ;
        RECT 2808.365 86.170 2808.695 86.185 ;
        RECT 711.430 85.870 2808.695 86.170 ;
        RECT 711.430 85.860 711.810 85.870 ;
        RECT 2808.365 85.855 2808.695 85.870 ;
      LAYER via3 ;
        RECT 711.460 2155.780 711.780 2156.100 ;
        RECT 711.460 85.860 711.780 86.180 ;
      LAYER met4 ;
        RECT 711.455 2155.775 711.785 2156.105 ;
        RECT 711.470 86.185 711.770 2155.775 ;
        RECT 711.455 85.855 711.785 86.185 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2614.785 1738.845 2615.875 1739.015 ;
      LAYER mcon ;
        RECT 2615.705 1738.845 2615.875 1739.015 ;
      LAYER met1 ;
        RECT 1772.910 1739.000 1773.230 1739.060 ;
        RECT 2614.725 1739.000 2615.015 1739.045 ;
        RECT 1772.910 1738.860 2615.015 1739.000 ;
        RECT 1772.910 1738.800 1773.230 1738.860 ;
        RECT 2614.725 1738.815 2615.015 1738.860 ;
        RECT 2615.645 1739.000 2615.935 1739.045 ;
        RECT 2818.950 1739.000 2819.270 1739.060 ;
        RECT 2615.645 1738.860 2819.270 1739.000 ;
        RECT 2615.645 1738.815 2615.935 1738.860 ;
        RECT 2818.950 1738.800 2819.270 1738.860 ;
        RECT 2818.950 16.900 2819.270 16.960 ;
        RECT 2827.690 16.900 2828.010 16.960 ;
        RECT 2818.950 16.760 2828.010 16.900 ;
        RECT 2818.950 16.700 2819.270 16.760 ;
        RECT 2827.690 16.700 2828.010 16.760 ;
      LAYER via ;
        RECT 1772.940 1738.800 1773.200 1739.060 ;
        RECT 2818.980 1738.800 2819.240 1739.060 ;
        RECT 2818.980 16.700 2819.240 16.960 ;
        RECT 2827.720 16.700 2827.980 16.960 ;
      LAYER met2 ;
        RECT 1772.930 1740.955 1773.210 1741.325 ;
        RECT 1773.000 1739.090 1773.140 1740.955 ;
        RECT 1772.940 1738.770 1773.200 1739.090 ;
        RECT 2818.980 1738.770 2819.240 1739.090 ;
        RECT 2819.040 16.990 2819.180 1738.770 ;
        RECT 2818.980 16.670 2819.240 16.990 ;
        RECT 2827.720 16.670 2827.980 16.990 ;
        RECT 2827.780 2.400 2827.920 16.670 ;
        RECT 2827.570 -4.800 2828.130 2.400 ;
      LAYER via2 ;
        RECT 1772.930 1741.000 1773.210 1741.280 ;
      LAYER met3 ;
        RECT 1755.835 1741.290 1759.835 1741.295 ;
        RECT 1772.905 1741.290 1773.235 1741.305 ;
        RECT 1755.835 1740.990 1773.235 1741.290 ;
        RECT 1755.835 1740.695 1759.835 1740.990 ;
        RECT 1772.905 1740.975 1773.235 1740.990 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2842.890 1307.115 2843.170 1307.485 ;
        RECT 2842.960 6.530 2843.100 1307.115 ;
        RECT 2842.960 6.390 2845.400 6.530 ;
        RECT 2845.260 2.400 2845.400 6.390 ;
        RECT 2845.050 -4.800 2845.610 2.400 ;
      LAYER via2 ;
        RECT 2842.890 1307.160 2843.170 1307.440 ;
      LAYER met3 ;
        RECT 714.190 1609.370 714.570 1609.380 ;
        RECT 715.810 1609.370 719.810 1609.375 ;
        RECT 714.190 1609.070 719.810 1609.370 ;
        RECT 714.190 1609.060 714.570 1609.070 ;
        RECT 715.810 1608.775 719.810 1609.070 ;
        RECT 714.190 1338.730 714.570 1338.740 ;
        RECT 716.950 1338.730 717.330 1338.740 ;
        RECT 714.190 1338.430 717.330 1338.730 ;
        RECT 714.190 1338.420 714.570 1338.430 ;
        RECT 716.950 1338.420 717.330 1338.430 ;
        RECT 716.950 1308.810 717.330 1308.820 ;
        RECT 716.950 1308.510 729.250 1308.810 ;
        RECT 716.950 1308.500 717.330 1308.510 ;
        RECT 728.950 1307.450 729.250 1308.510 ;
        RECT 2842.865 1307.450 2843.195 1307.465 ;
        RECT 728.950 1307.150 2843.195 1307.450 ;
        RECT 2842.865 1307.135 2843.195 1307.150 ;
      LAYER via3 ;
        RECT 714.220 1609.060 714.540 1609.380 ;
        RECT 714.220 1338.420 714.540 1338.740 ;
        RECT 716.980 1338.420 717.300 1338.740 ;
        RECT 716.980 1308.500 717.300 1308.820 ;
      LAYER met4 ;
        RECT 714.215 1609.055 714.545 1609.385 ;
        RECT 714.230 1338.745 714.530 1609.055 ;
        RECT 714.215 1338.415 714.545 1338.745 ;
        RECT 716.975 1338.415 717.305 1338.745 ;
        RECT 716.990 1308.825 717.290 1338.415 ;
        RECT 716.975 1308.495 717.305 1308.825 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1710.810 24.040 1711.130 24.100 ;
        RECT 2863.110 24.040 2863.430 24.100 ;
        RECT 1710.810 23.900 2863.430 24.040 ;
        RECT 1710.810 23.840 1711.130 23.900 ;
        RECT 2863.110 23.840 2863.430 23.900 ;
      LAYER via ;
        RECT 1710.840 23.840 1711.100 24.100 ;
        RECT 2863.140 23.840 2863.400 24.100 ;
      LAYER met2 ;
        RECT 1707.660 1323.690 1707.940 1327.135 ;
        RECT 1707.660 1323.550 1711.040 1323.690 ;
        RECT 1707.660 1323.135 1707.940 1323.550 ;
        RECT 1710.900 24.130 1711.040 1323.550 ;
        RECT 1710.840 23.810 1711.100 24.130 ;
        RECT 2863.140 23.810 2863.400 24.130 ;
        RECT 2863.200 2.400 2863.340 23.810 ;
        RECT 2862.990 -4.800 2863.550 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1770.610 2139.180 1770.930 2139.240 ;
        RECT 2818.490 2139.180 2818.810 2139.240 ;
        RECT 1770.610 2139.040 2818.810 2139.180 ;
        RECT 1770.610 2138.980 1770.930 2139.040 ;
        RECT 2818.490 2138.980 2818.810 2139.040 ;
        RECT 2818.490 18.260 2818.810 18.320 ;
        RECT 2881.050 18.260 2881.370 18.320 ;
        RECT 2818.490 18.120 2881.370 18.260 ;
        RECT 2818.490 18.060 2818.810 18.120 ;
        RECT 2881.050 18.060 2881.370 18.120 ;
      LAYER via ;
        RECT 1770.640 2138.980 1770.900 2139.240 ;
        RECT 2818.520 2138.980 2818.780 2139.240 ;
        RECT 2818.520 18.060 2818.780 18.320 ;
        RECT 2881.080 18.060 2881.340 18.320 ;
      LAYER met2 ;
        RECT 1770.630 2143.515 1770.910 2143.885 ;
        RECT 1770.700 2139.270 1770.840 2143.515 ;
        RECT 1770.640 2138.950 1770.900 2139.270 ;
        RECT 2818.520 2138.950 2818.780 2139.270 ;
        RECT 2818.580 18.350 2818.720 2138.950 ;
        RECT 2818.520 18.030 2818.780 18.350 ;
        RECT 2881.080 18.030 2881.340 18.350 ;
        RECT 2881.140 2.400 2881.280 18.030 ;
        RECT 2880.930 -4.800 2881.490 2.400 ;
      LAYER via2 ;
        RECT 1770.630 2143.560 1770.910 2143.840 ;
      LAYER met3 ;
        RECT 1755.835 2143.850 1759.835 2143.855 ;
        RECT 1770.605 2143.850 1770.935 2143.865 ;
        RECT 1755.835 2143.550 1770.935 2143.850 ;
        RECT 1755.835 2143.255 1759.835 2143.550 ;
        RECT 1770.605 2143.535 1770.935 2143.550 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 779.770 2376.500 780.090 2376.560 ;
        RECT 1559.470 2376.500 1559.790 2376.560 ;
        RECT 779.770 2376.360 1559.790 2376.500 ;
        RECT 779.770 2376.300 780.090 2376.360 ;
        RECT 1559.470 2376.300 1559.790 2376.360 ;
        RECT 2898.070 2.960 2898.390 3.020 ;
        RECT 2898.990 2.960 2899.310 3.020 ;
        RECT 2898.070 2.820 2899.310 2.960 ;
        RECT 2898.070 2.760 2898.390 2.820 ;
        RECT 2898.990 2.760 2899.310 2.820 ;
      LAYER via ;
        RECT 779.800 2376.300 780.060 2376.560 ;
        RECT 1559.500 2376.300 1559.760 2376.560 ;
        RECT 2898.100 2.760 2898.360 3.020 ;
        RECT 2899.020 2.760 2899.280 3.020 ;
      LAYER met2 ;
        RECT 779.380 2376.330 779.660 2377.880 ;
        RECT 1559.490 2377.435 1559.770 2377.805 ;
        RECT 2898.090 2377.435 2898.370 2377.805 ;
        RECT 1559.560 2376.590 1559.700 2377.435 ;
        RECT 779.800 2376.330 780.060 2376.590 ;
        RECT 779.380 2376.270 780.060 2376.330 ;
        RECT 1559.500 2376.270 1559.760 2376.590 ;
        RECT 779.380 2376.190 780.000 2376.270 ;
        RECT 779.380 2373.880 779.660 2376.190 ;
        RECT 2898.160 3.050 2898.300 2377.435 ;
        RECT 2898.100 2.730 2898.360 3.050 ;
        RECT 2899.020 2.730 2899.280 3.050 ;
        RECT 2899.080 2.400 2899.220 2.730 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
      LAYER via2 ;
        RECT 1559.490 2377.480 1559.770 2377.760 ;
        RECT 2898.090 2377.480 2898.370 2377.760 ;
      LAYER met3 ;
        RECT 1559.465 2377.770 1559.795 2377.785 ;
        RECT 2898.065 2377.770 2898.395 2377.785 ;
        RECT 1559.465 2377.470 2898.395 2377.770 ;
        RECT 1559.465 2377.455 1559.795 2377.470 ;
        RECT 2898.065 2377.455 2898.395 2377.470 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1739.860 2374.290 1740.140 2377.880 ;
        RECT 1741.190 2374.290 1741.470 2374.405 ;
        RECT 1739.860 2374.150 1741.470 2374.290 ;
        RECT 1739.860 2373.880 1740.140 2374.150 ;
        RECT 1741.190 2374.035 1741.470 2374.150 ;
        RECT 846.950 19.875 847.230 20.245 ;
        RECT 847.020 2.400 847.160 19.875 ;
        RECT 846.810 -4.800 847.370 2.400 ;
      LAYER via2 ;
        RECT 1741.190 2374.080 1741.470 2374.360 ;
        RECT 846.950 19.920 847.230 20.200 ;
      LAYER met3 ;
        RECT 1741.165 2374.370 1741.495 2374.385 ;
        RECT 1742.750 2374.370 1743.130 2374.380 ;
        RECT 1741.165 2374.070 1743.130 2374.370 ;
        RECT 1741.165 2374.055 1741.495 2374.070 ;
        RECT 1742.750 2374.060 1743.130 2374.070 ;
        RECT 846.925 20.210 847.255 20.225 ;
        RECT 1742.750 20.210 1743.130 20.220 ;
        RECT 846.925 19.910 1743.130 20.210 ;
        RECT 846.925 19.895 847.255 19.910 ;
        RECT 1742.750 19.900 1743.130 19.910 ;
      LAYER via3 ;
        RECT 1742.780 2374.060 1743.100 2374.380 ;
        RECT 1742.780 19.900 1743.100 20.220 ;
      LAYER met4 ;
        RECT 1742.775 2374.055 1743.105 2374.385 ;
        RECT 1742.790 20.225 1743.090 2374.055 ;
        RECT 1742.775 19.895 1743.105 20.225 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 864.870 25.400 865.190 25.460 ;
        RECT 980.330 25.400 980.650 25.460 ;
        RECT 864.870 25.260 980.650 25.400 ;
        RECT 864.870 25.200 865.190 25.260 ;
        RECT 980.330 25.200 980.650 25.260 ;
      LAYER via ;
        RECT 864.900 25.200 865.160 25.460 ;
        RECT 980.360 25.200 980.620 25.460 ;
      LAYER met2 ;
        RECT 984.540 1323.690 984.820 1327.135 ;
        RECT 980.420 1323.550 984.820 1323.690 ;
        RECT 980.420 25.490 980.560 1323.550 ;
        RECT 984.540 1323.135 984.820 1323.550 ;
        RECT 864.900 25.170 865.160 25.490 ;
        RECT 980.360 25.170 980.620 25.490 ;
        RECT 864.960 2.400 865.100 25.170 ;
        RECT 864.750 -4.800 865.310 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 882.810 25.740 883.130 25.800 ;
        RECT 966.070 25.740 966.390 25.800 ;
        RECT 882.810 25.600 966.390 25.740 ;
        RECT 882.810 25.540 883.130 25.600 ;
        RECT 966.070 25.540 966.390 25.600 ;
      LAYER via ;
        RECT 882.840 25.540 883.100 25.800 ;
        RECT 966.100 25.540 966.360 25.800 ;
      LAYER met2 ;
        RECT 967.060 1323.690 967.340 1327.135 ;
        RECT 966.160 1323.550 967.340 1323.690 ;
        RECT 966.160 25.830 966.300 1323.550 ;
        RECT 967.060 1323.135 967.340 1323.550 ;
        RECT 882.840 25.510 883.100 25.830 ;
        RECT 966.100 25.510 966.360 25.830 ;
        RECT 882.900 2.400 883.040 25.510 ;
        RECT 882.690 -4.800 883.250 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 713.145 1905.785 713.315 1912.415 ;
        RECT 713.605 1832.005 713.775 1860.055 ;
        RECT 712.225 1747.345 712.395 1769.955 ;
        RECT 712.225 1637.865 712.395 1661.495 ;
        RECT 717.285 1631.745 717.455 1657.755 ;
        RECT 730.625 1326.085 730.795 1332.715 ;
        RECT 1148.305 1326.425 1148.475 1332.715 ;
      LAYER mcon ;
        RECT 713.145 1912.245 713.315 1912.415 ;
        RECT 713.605 1859.885 713.775 1860.055 ;
        RECT 712.225 1769.785 712.395 1769.955 ;
        RECT 712.225 1661.325 712.395 1661.495 ;
        RECT 717.285 1657.585 717.455 1657.755 ;
        RECT 730.625 1332.545 730.795 1332.715 ;
        RECT 1148.305 1332.545 1148.475 1332.715 ;
      LAYER met1 ;
        RECT 975.270 2388.060 975.590 2388.120 ;
        RECT 979.870 2388.060 980.190 2388.120 ;
        RECT 975.270 2387.920 980.190 2388.060 ;
        RECT 975.270 2387.860 975.590 2387.920 ;
        RECT 979.870 2387.860 980.190 2387.920 ;
        RECT 713.070 1936.200 713.390 1936.260 ;
        RECT 717.670 1936.200 717.990 1936.260 ;
        RECT 713.070 1936.060 717.990 1936.200 ;
        RECT 713.070 1936.000 713.390 1936.060 ;
        RECT 717.670 1936.000 717.990 1936.060 ;
        RECT 713.070 1912.400 713.390 1912.460 ;
        RECT 712.875 1912.260 713.390 1912.400 ;
        RECT 713.070 1912.200 713.390 1912.260 ;
        RECT 713.070 1905.940 713.390 1906.000 ;
        RECT 712.875 1905.800 713.390 1905.940 ;
        RECT 713.070 1905.740 713.390 1905.800 ;
        RECT 713.530 1860.040 713.850 1860.100 ;
        RECT 713.335 1859.900 713.850 1860.040 ;
        RECT 713.530 1859.840 713.850 1859.900 ;
        RECT 713.530 1832.160 713.850 1832.220 ;
        RECT 713.335 1832.020 713.850 1832.160 ;
        RECT 713.530 1831.960 713.850 1832.020 ;
        RECT 712.165 1769.940 712.455 1769.985 ;
        RECT 713.530 1769.940 713.850 1770.000 ;
        RECT 712.165 1769.800 713.850 1769.940 ;
        RECT 712.165 1769.755 712.455 1769.800 ;
        RECT 713.530 1769.740 713.850 1769.800 ;
        RECT 712.150 1747.500 712.470 1747.560 ;
        RECT 711.955 1747.360 712.470 1747.500 ;
        RECT 712.150 1747.300 712.470 1747.360 ;
        RECT 712.150 1661.480 712.470 1661.540 ;
        RECT 711.955 1661.340 712.470 1661.480 ;
        RECT 712.150 1661.280 712.470 1661.340 ;
        RECT 717.210 1657.740 717.530 1657.800 ;
        RECT 717.015 1657.600 717.530 1657.740 ;
        RECT 717.210 1657.540 717.530 1657.600 ;
        RECT 712.165 1638.020 712.455 1638.065 ;
        RECT 713.990 1638.020 714.310 1638.080 ;
        RECT 712.165 1637.880 714.310 1638.020 ;
        RECT 712.165 1637.835 712.455 1637.880 ;
        RECT 713.990 1637.820 714.310 1637.880 ;
        RECT 713.530 1631.900 713.850 1631.960 ;
        RECT 717.225 1631.900 717.515 1631.945 ;
        RECT 713.530 1631.760 717.515 1631.900 ;
        RECT 713.530 1631.700 713.850 1631.760 ;
        RECT 717.225 1631.715 717.515 1631.760 ;
        RECT 730.565 1332.700 730.855 1332.745 ;
        RECT 1148.245 1332.700 1148.535 1332.745 ;
        RECT 730.565 1332.560 1148.535 1332.700 ;
        RECT 730.565 1332.515 730.855 1332.560 ;
        RECT 1148.245 1332.515 1148.535 1332.560 ;
        RECT 1148.230 1326.580 1148.550 1326.640 ;
        RECT 1148.035 1326.440 1148.550 1326.580 ;
        RECT 1148.230 1326.380 1148.550 1326.440 ;
        RECT 730.550 1326.240 730.870 1326.300 ;
        RECT 730.355 1326.100 730.870 1326.240 ;
        RECT 730.550 1326.040 730.870 1326.100 ;
        RECT 897.990 20.640 898.310 20.700 ;
        RECT 900.750 20.640 901.070 20.700 ;
        RECT 897.990 20.500 901.070 20.640 ;
        RECT 897.990 20.440 898.310 20.500 ;
        RECT 900.750 20.440 901.070 20.500 ;
        RECT 1008.390 20.640 1008.710 20.700 ;
        RECT 1013.450 20.640 1013.770 20.700 ;
        RECT 1008.390 20.500 1013.770 20.640 ;
        RECT 1008.390 20.440 1008.710 20.500 ;
        RECT 1013.450 20.440 1013.770 20.500 ;
      LAYER via ;
        RECT 975.300 2387.860 975.560 2388.120 ;
        RECT 979.900 2387.860 980.160 2388.120 ;
        RECT 713.100 1936.000 713.360 1936.260 ;
        RECT 717.700 1936.000 717.960 1936.260 ;
        RECT 713.100 1912.200 713.360 1912.460 ;
        RECT 713.100 1905.740 713.360 1906.000 ;
        RECT 713.560 1859.840 713.820 1860.100 ;
        RECT 713.560 1831.960 713.820 1832.220 ;
        RECT 713.560 1769.740 713.820 1770.000 ;
        RECT 712.180 1747.300 712.440 1747.560 ;
        RECT 712.180 1661.280 712.440 1661.540 ;
        RECT 717.240 1657.540 717.500 1657.800 ;
        RECT 714.020 1637.820 714.280 1638.080 ;
        RECT 713.560 1631.700 713.820 1631.960 ;
        RECT 1148.260 1326.380 1148.520 1326.640 ;
        RECT 730.580 1326.040 730.840 1326.300 ;
        RECT 898.020 20.440 898.280 20.700 ;
        RECT 900.780 20.440 901.040 20.700 ;
        RECT 1008.420 20.440 1008.680 20.700 ;
        RECT 1013.480 20.440 1013.740 20.700 ;
      LAYER met2 ;
        RECT 759.090 2394.435 759.370 2394.805 ;
        RECT 759.160 2392.085 759.300 2394.435 ;
        RECT 810.610 2393.755 810.890 2394.125 ;
        RECT 855.690 2393.755 855.970 2394.125 ;
        RECT 903.530 2393.755 903.810 2394.125 ;
        RECT 810.680 2392.085 810.820 2393.755 ;
        RECT 855.760 2392.085 855.900 2393.755 ;
        RECT 903.600 2392.085 903.740 2393.755 ;
        RECT 1131.690 2393.075 1131.970 2393.445 ;
        RECT 759.090 2391.715 759.370 2392.085 ;
        RECT 810.610 2391.715 810.890 2392.085 ;
        RECT 855.690 2391.715 855.970 2392.085 ;
        RECT 903.530 2391.715 903.810 2392.085 ;
        RECT 975.290 2391.715 975.570 2392.085 ;
        RECT 975.360 2388.150 975.500 2391.715 ;
        RECT 975.300 2387.830 975.560 2388.150 ;
        RECT 979.900 2387.830 980.160 2388.150 ;
        RECT 979.960 2377.690 980.100 2387.830 ;
        RECT 1131.760 2377.880 1131.900 2393.075 ;
        RECT 981.780 2377.690 982.060 2377.880 ;
        RECT 979.960 2377.550 982.060 2377.690 ;
        RECT 821.190 2374.715 821.470 2375.085 ;
        RECT 823.490 2374.715 823.770 2375.085 ;
        RECT 821.260 2374.290 821.400 2374.715 ;
        RECT 823.560 2374.290 823.700 2374.715 ;
        RECT 821.260 2374.150 823.700 2374.290 ;
        RECT 981.780 2373.880 982.060 2377.550 ;
        RECT 1021.290 2374.970 1021.570 2375.085 ;
        RECT 1022.260 2374.970 1022.540 2377.880 ;
        RECT 1021.290 2374.830 1022.540 2374.970 ;
        RECT 1021.290 2374.715 1021.570 2374.830 ;
        RECT 1022.260 2373.880 1022.540 2374.830 ;
        RECT 1037.850 2374.290 1038.130 2374.405 ;
        RECT 1039.740 2374.290 1040.020 2377.880 ;
        RECT 1037.850 2374.150 1040.020 2374.290 ;
        RECT 1037.850 2374.035 1038.130 2374.150 ;
        RECT 1039.740 2373.880 1040.020 2374.150 ;
        RECT 1131.740 2373.880 1132.020 2377.880 ;
        RECT 1304.190 2374.290 1304.470 2374.405 ;
        RECT 1305.620 2374.290 1305.900 2377.880 ;
        RECT 1304.190 2374.150 1305.900 2374.290 ;
        RECT 1304.190 2374.035 1304.470 2374.150 ;
        RECT 1305.620 2373.880 1305.900 2374.150 ;
        RECT 716.770 2218.315 717.050 2218.685 ;
        RECT 716.840 2201.005 716.980 2218.315 ;
        RECT 716.770 2200.635 717.050 2201.005 ;
        RECT 715.850 2195.195 716.130 2195.565 ;
        RECT 715.920 2187.405 716.060 2195.195 ;
        RECT 716.310 2194.515 716.590 2194.885 ;
        RECT 715.850 2187.035 716.130 2187.405 ;
        RECT 716.380 2184.005 716.520 2194.515 ;
        RECT 717.690 2187.715 717.970 2188.085 ;
        RECT 716.310 2183.635 716.590 2184.005 ;
        RECT 717.760 2180.605 717.900 2187.715 ;
        RECT 717.690 2180.235 717.970 2180.605 ;
        RECT 718.610 2000.715 718.890 2001.085 ;
        RECT 714.010 1997.315 714.290 1997.685 ;
        RECT 714.080 1956.885 714.220 1997.315 ;
        RECT 718.680 1997.005 718.820 2000.715 ;
        RECT 718.610 1996.635 718.890 1997.005 ;
        RECT 714.010 1956.515 714.290 1956.885 ;
        RECT 713.090 1946.315 713.370 1946.685 ;
        RECT 713.160 1936.290 713.300 1946.315 ;
        RECT 713.100 1935.970 713.360 1936.290 ;
        RECT 717.700 1935.970 717.960 1936.290 ;
        RECT 713.550 1924.555 713.830 1924.925 ;
        RECT 713.090 1921.835 713.370 1922.205 ;
        RECT 713.160 1912.490 713.300 1921.835 ;
        RECT 713.100 1912.170 713.360 1912.490 ;
        RECT 713.090 1911.635 713.370 1912.005 ;
        RECT 713.160 1906.565 713.300 1911.635 ;
        RECT 713.090 1906.195 713.370 1906.565 ;
        RECT 713.100 1905.885 713.360 1906.030 ;
        RECT 713.090 1905.515 713.370 1905.885 ;
        RECT 713.620 1860.130 713.760 1924.555 ;
        RECT 717.760 1909.285 717.900 1935.970 ;
        RECT 717.690 1908.915 717.970 1909.285 ;
        RECT 713.560 1859.810 713.820 1860.130 ;
        RECT 713.560 1831.930 713.820 1832.250 ;
        RECT 713.620 1820.885 713.760 1831.930 ;
        RECT 713.550 1820.515 713.830 1820.885 ;
        RECT 713.550 1776.995 713.830 1777.365 ;
        RECT 713.620 1770.030 713.760 1776.995 ;
        RECT 713.560 1769.710 713.820 1770.030 ;
        RECT 712.180 1747.270 712.440 1747.590 ;
        RECT 710.330 1721.235 710.610 1721.605 ;
        RECT 710.400 1718.885 710.540 1721.235 ;
        RECT 710.330 1718.515 710.610 1718.885 ;
        RECT 712.240 1681.485 712.380 1747.270 ;
        RECT 713.090 1738.915 713.370 1739.285 ;
        RECT 712.170 1681.115 712.450 1681.485 ;
        RECT 713.160 1671.285 713.300 1738.915 ;
        RECT 713.090 1670.915 713.370 1671.285 ;
        RECT 717.230 1664.115 717.510 1664.485 ;
        RECT 712.170 1662.075 712.450 1662.445 ;
        RECT 712.240 1661.570 712.380 1662.075 ;
        RECT 712.180 1661.250 712.440 1661.570 ;
        RECT 717.300 1657.830 717.440 1664.115 ;
        RECT 717.240 1657.510 717.500 1657.830 ;
        RECT 713.550 1652.555 713.830 1652.925 ;
        RECT 713.620 1638.645 713.760 1652.555 ;
        RECT 713.550 1638.275 713.830 1638.645 ;
        RECT 714.020 1637.965 714.280 1638.110 ;
        RECT 714.010 1637.595 714.290 1637.965 ;
        RECT 713.560 1631.845 713.820 1631.990 ;
        RECT 713.550 1631.475 713.830 1631.845 ;
        RECT 1148.260 1326.525 1148.520 1326.670 ;
        RECT 730.570 1326.155 730.850 1326.525 ;
        RECT 1008.870 1326.410 1009.150 1326.525 ;
        RECT 1008.480 1326.270 1009.150 1326.410 ;
        RECT 730.580 1326.010 730.840 1326.155 ;
        RECT 898.470 1325.730 898.750 1325.845 ;
        RECT 898.080 1325.590 898.750 1325.730 ;
        RECT 898.080 20.730 898.220 1325.590 ;
        RECT 898.470 1325.475 898.750 1325.590 ;
        RECT 953.670 1158.875 953.950 1159.245 ;
        RECT 953.740 1111.645 953.880 1158.875 ;
        RECT 953.670 1111.275 953.950 1111.645 ;
        RECT 953.670 1062.315 953.950 1062.685 ;
        RECT 953.740 1015.085 953.880 1062.315 ;
        RECT 953.670 1014.715 953.950 1015.085 ;
        RECT 952.750 965.755 953.030 966.125 ;
        RECT 952.820 919.205 952.960 965.755 ;
        RECT 952.750 918.835 953.030 919.205 ;
        RECT 952.750 869.195 953.030 869.565 ;
        RECT 952.820 821.285 952.960 869.195 ;
        RECT 952.750 820.915 953.030 821.285 ;
        RECT 953.670 771.955 953.950 772.325 ;
        RECT 953.740 724.725 953.880 771.955 ;
        RECT 953.670 724.355 953.950 724.725 ;
        RECT 953.670 674.715 953.950 675.085 ;
        RECT 953.740 628.165 953.880 674.715 ;
        RECT 953.670 627.795 953.950 628.165 ;
        RECT 952.750 426.515 953.030 426.885 ;
        RECT 952.820 380.645 952.960 426.515 ;
        RECT 952.750 380.275 953.030 380.645 ;
        RECT 953.670 288.475 953.950 288.845 ;
        RECT 953.740 241.925 953.880 288.475 ;
        RECT 953.670 241.555 953.950 241.925 ;
        RECT 952.750 192.595 953.030 192.965 ;
        RECT 952.820 146.045 952.960 192.595 ;
        RECT 952.750 145.675 953.030 146.045 ;
        RECT 953.670 95.355 953.950 95.725 ;
        RECT 953.740 48.805 953.880 95.355 ;
        RECT 953.670 48.435 953.950 48.805 ;
        RECT 954.130 24.635 954.410 25.005 ;
        RECT 898.020 20.410 898.280 20.730 ;
        RECT 900.780 20.410 901.040 20.730 ;
        RECT 900.840 2.400 900.980 20.410 ;
        RECT 954.200 2.400 954.340 24.635 ;
        RECT 1008.480 20.730 1008.620 1326.270 ;
        RECT 1008.870 1326.155 1009.150 1326.270 ;
        RECT 1148.250 1326.155 1148.530 1326.525 ;
        RECT 1008.420 20.410 1008.680 20.730 ;
        RECT 1013.480 20.410 1013.740 20.730 ;
        RECT 1013.540 2.400 1013.680 20.410 ;
        RECT 1150.550 18.515 1150.830 18.885 ;
        RECT 1037.390 14.435 1037.670 14.805 ;
        RECT 1037.460 2.400 1037.600 14.435 ;
        RECT 1150.620 2.400 1150.760 18.515 ;
        RECT 900.630 -4.800 901.190 2.400 ;
        RECT 953.990 -4.800 954.550 2.400 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
        RECT 1150.410 -4.800 1150.970 2.400 ;
      LAYER via2 ;
        RECT 759.090 2394.480 759.370 2394.760 ;
        RECT 810.610 2393.800 810.890 2394.080 ;
        RECT 855.690 2393.800 855.970 2394.080 ;
        RECT 903.530 2393.800 903.810 2394.080 ;
        RECT 1131.690 2393.120 1131.970 2393.400 ;
        RECT 759.090 2391.760 759.370 2392.040 ;
        RECT 810.610 2391.760 810.890 2392.040 ;
        RECT 855.690 2391.760 855.970 2392.040 ;
        RECT 903.530 2391.760 903.810 2392.040 ;
        RECT 975.290 2391.760 975.570 2392.040 ;
        RECT 821.190 2374.760 821.470 2375.040 ;
        RECT 823.490 2374.760 823.770 2375.040 ;
        RECT 1021.290 2374.760 1021.570 2375.040 ;
        RECT 1037.850 2374.080 1038.130 2374.360 ;
        RECT 1304.190 2374.080 1304.470 2374.360 ;
        RECT 716.770 2218.360 717.050 2218.640 ;
        RECT 716.770 2200.680 717.050 2200.960 ;
        RECT 715.850 2195.240 716.130 2195.520 ;
        RECT 716.310 2194.560 716.590 2194.840 ;
        RECT 715.850 2187.080 716.130 2187.360 ;
        RECT 717.690 2187.760 717.970 2188.040 ;
        RECT 716.310 2183.680 716.590 2183.960 ;
        RECT 717.690 2180.280 717.970 2180.560 ;
        RECT 718.610 2000.760 718.890 2001.040 ;
        RECT 714.010 1997.360 714.290 1997.640 ;
        RECT 718.610 1996.680 718.890 1996.960 ;
        RECT 714.010 1956.560 714.290 1956.840 ;
        RECT 713.090 1946.360 713.370 1946.640 ;
        RECT 713.550 1924.600 713.830 1924.880 ;
        RECT 713.090 1921.880 713.370 1922.160 ;
        RECT 713.090 1911.680 713.370 1911.960 ;
        RECT 713.090 1906.240 713.370 1906.520 ;
        RECT 713.090 1905.560 713.370 1905.840 ;
        RECT 717.690 1908.960 717.970 1909.240 ;
        RECT 713.550 1820.560 713.830 1820.840 ;
        RECT 713.550 1777.040 713.830 1777.320 ;
        RECT 710.330 1721.280 710.610 1721.560 ;
        RECT 710.330 1718.560 710.610 1718.840 ;
        RECT 713.090 1738.960 713.370 1739.240 ;
        RECT 712.170 1681.160 712.450 1681.440 ;
        RECT 713.090 1670.960 713.370 1671.240 ;
        RECT 717.230 1664.160 717.510 1664.440 ;
        RECT 712.170 1662.120 712.450 1662.400 ;
        RECT 713.550 1652.600 713.830 1652.880 ;
        RECT 713.550 1638.320 713.830 1638.600 ;
        RECT 714.010 1637.640 714.290 1637.920 ;
        RECT 713.550 1631.520 713.830 1631.800 ;
        RECT 730.570 1326.200 730.850 1326.480 ;
        RECT 898.470 1325.520 898.750 1325.800 ;
        RECT 953.670 1158.920 953.950 1159.200 ;
        RECT 953.670 1111.320 953.950 1111.600 ;
        RECT 953.670 1062.360 953.950 1062.640 ;
        RECT 953.670 1014.760 953.950 1015.040 ;
        RECT 952.750 965.800 953.030 966.080 ;
        RECT 952.750 918.880 953.030 919.160 ;
        RECT 952.750 869.240 953.030 869.520 ;
        RECT 952.750 820.960 953.030 821.240 ;
        RECT 953.670 772.000 953.950 772.280 ;
        RECT 953.670 724.400 953.950 724.680 ;
        RECT 953.670 674.760 953.950 675.040 ;
        RECT 953.670 627.840 953.950 628.120 ;
        RECT 952.750 426.560 953.030 426.840 ;
        RECT 952.750 380.320 953.030 380.600 ;
        RECT 953.670 288.520 953.950 288.800 ;
        RECT 953.670 241.600 953.950 241.880 ;
        RECT 952.750 192.640 953.030 192.920 ;
        RECT 952.750 145.720 953.030 146.000 ;
        RECT 953.670 95.400 953.950 95.680 ;
        RECT 953.670 48.480 953.950 48.760 ;
        RECT 954.130 24.680 954.410 24.960 ;
        RECT 1008.870 1326.200 1009.150 1326.480 ;
        RECT 1148.250 1326.200 1148.530 1326.480 ;
        RECT 1150.550 18.560 1150.830 18.840 ;
        RECT 1037.390 14.480 1037.670 14.760 ;
      LAYER met3 ;
        RECT 759.065 2394.770 759.395 2394.785 ;
        RECT 759.065 2394.470 788.130 2394.770 ;
        RECT 759.065 2394.455 759.395 2394.470 ;
        RECT 787.830 2394.090 788.130 2394.470 ;
        RECT 810.585 2394.090 810.915 2394.105 ;
        RECT 787.830 2393.790 810.915 2394.090 ;
        RECT 810.585 2393.775 810.915 2393.790 ;
        RECT 855.665 2394.090 855.995 2394.105 ;
        RECT 903.505 2394.090 903.835 2394.105 ;
        RECT 855.665 2393.790 903.835 2394.090 ;
        RECT 855.665 2393.775 855.995 2393.790 ;
        RECT 903.505 2393.775 903.835 2393.790 ;
        RECT 730.750 2393.410 731.130 2393.420 ;
        RECT 1131.665 2393.410 1131.995 2393.425 ;
        RECT 730.750 2393.110 1131.995 2393.410 ;
        RECT 730.750 2393.100 731.130 2393.110 ;
        RECT 1131.665 2393.095 1131.995 2393.110 ;
        RECT 729.830 2392.050 730.210 2392.060 ;
        RECT 759.065 2392.050 759.395 2392.065 ;
        RECT 729.830 2391.750 759.395 2392.050 ;
        RECT 729.830 2391.740 730.210 2391.750 ;
        RECT 759.065 2391.735 759.395 2391.750 ;
        RECT 810.585 2392.050 810.915 2392.065 ;
        RECT 855.665 2392.050 855.995 2392.065 ;
        RECT 810.585 2391.750 855.995 2392.050 ;
        RECT 810.585 2391.735 810.915 2391.750 ;
        RECT 855.665 2391.735 855.995 2391.750 ;
        RECT 903.505 2392.050 903.835 2392.065 ;
        RECT 975.265 2392.050 975.595 2392.065 ;
        RECT 903.505 2391.750 975.595 2392.050 ;
        RECT 903.505 2391.735 903.835 2391.750 ;
        RECT 975.265 2391.735 975.595 2391.750 ;
        RECT 738.110 2375.050 738.490 2375.060 ;
        RECT 821.165 2375.050 821.495 2375.065 ;
        RECT 738.110 2374.750 821.495 2375.050 ;
        RECT 738.110 2374.740 738.490 2374.750 ;
        RECT 821.165 2374.735 821.495 2374.750 ;
        RECT 823.465 2375.050 823.795 2375.065 ;
        RECT 1021.265 2375.050 1021.595 2375.065 ;
        RECT 823.465 2374.750 1021.595 2375.050 ;
        RECT 823.465 2374.735 823.795 2374.750 ;
        RECT 1021.265 2374.735 1021.595 2374.750 ;
        RECT 739.030 2374.370 739.410 2374.380 ;
        RECT 1037.825 2374.370 1038.155 2374.385 ;
        RECT 1304.165 2374.380 1304.495 2374.385 ;
        RECT 1303.910 2374.370 1304.495 2374.380 ;
        RECT 739.030 2374.070 1038.155 2374.370 ;
        RECT 1303.710 2374.070 1304.495 2374.370 ;
        RECT 739.030 2374.060 739.410 2374.070 ;
        RECT 1037.825 2374.055 1038.155 2374.070 ;
        RECT 1303.910 2374.060 1304.495 2374.070 ;
        RECT 1304.165 2374.055 1304.495 2374.060 ;
        RECT 723.390 2370.290 723.770 2370.300 ;
        RECT 1303.910 2370.290 1304.290 2370.300 ;
        RECT 723.390 2369.990 1304.290 2370.290 ;
        RECT 723.390 2369.980 723.770 2369.990 ;
        RECT 1303.910 2369.980 1304.290 2369.990 ;
        RECT 726.150 2366.890 726.530 2366.900 ;
        RECT 739.030 2366.890 739.410 2366.900 ;
        RECT 726.150 2366.590 739.410 2366.890 ;
        RECT 726.150 2366.580 726.530 2366.590 ;
        RECT 739.030 2366.580 739.410 2366.590 ;
        RECT 725.230 2366.210 725.610 2366.220 ;
        RECT 738.110 2366.210 738.490 2366.220 ;
        RECT 725.230 2365.910 738.490 2366.210 ;
        RECT 725.230 2365.900 725.610 2365.910 ;
        RECT 738.110 2365.900 738.490 2365.910 ;
        RECT 716.745 2218.650 717.075 2218.665 ;
        RECT 718.790 2218.650 719.170 2218.660 ;
        RECT 716.745 2218.350 719.170 2218.650 ;
        RECT 716.745 2218.335 717.075 2218.350 ;
        RECT 718.790 2218.340 719.170 2218.350 ;
        RECT 716.745 2200.970 717.075 2200.985 ;
        RECT 717.870 2200.970 718.250 2200.980 ;
        RECT 716.745 2200.670 718.250 2200.970 ;
        RECT 716.745 2200.655 717.075 2200.670 ;
        RECT 717.870 2200.660 718.250 2200.670 ;
        RECT 715.825 2195.530 716.155 2195.545 ;
        RECT 718.790 2195.530 719.170 2195.540 ;
        RECT 715.825 2195.230 719.170 2195.530 ;
        RECT 715.825 2195.215 716.155 2195.230 ;
        RECT 718.790 2195.220 719.170 2195.230 ;
        RECT 716.285 2194.850 716.615 2194.865 ;
        RECT 718.790 2194.850 719.170 2194.860 ;
        RECT 716.285 2194.550 719.170 2194.850 ;
        RECT 716.285 2194.535 716.615 2194.550 ;
        RECT 718.790 2194.540 719.170 2194.550 ;
        RECT 717.665 2188.050 717.995 2188.065 ;
        RECT 718.790 2188.050 719.170 2188.060 ;
        RECT 717.665 2187.750 719.170 2188.050 ;
        RECT 717.665 2187.735 717.995 2187.750 ;
        RECT 718.790 2187.740 719.170 2187.750 ;
        RECT 715.825 2187.370 716.155 2187.385 ;
        RECT 718.790 2187.370 719.170 2187.380 ;
        RECT 715.825 2187.070 719.170 2187.370 ;
        RECT 715.825 2187.055 716.155 2187.070 ;
        RECT 718.790 2187.060 719.170 2187.070 ;
        RECT 716.285 2183.970 716.615 2183.985 ;
        RECT 718.790 2183.970 719.170 2183.980 ;
        RECT 716.285 2183.670 719.170 2183.970 ;
        RECT 716.285 2183.655 716.615 2183.670 ;
        RECT 718.790 2183.660 719.170 2183.670 ;
        RECT 717.665 2180.570 717.995 2180.585 ;
        RECT 718.790 2180.570 719.170 2180.580 ;
        RECT 717.665 2180.270 719.170 2180.570 ;
        RECT 717.665 2180.255 717.995 2180.270 ;
        RECT 718.790 2180.260 719.170 2180.270 ;
        RECT 718.585 2001.060 718.915 2001.065 ;
        RECT 718.585 2001.050 719.170 2001.060 ;
        RECT 718.585 2000.750 719.370 2001.050 ;
        RECT 718.585 2000.740 719.170 2000.750 ;
        RECT 718.585 2000.735 718.915 2000.740 ;
        RECT 713.985 1997.650 714.315 1997.665 ;
        RECT 718.790 1997.650 719.170 1997.660 ;
        RECT 713.985 1997.350 719.170 1997.650 ;
        RECT 713.985 1997.335 714.315 1997.350 ;
        RECT 718.790 1997.340 719.170 1997.350 ;
        RECT 718.585 1996.980 718.915 1996.985 ;
        RECT 718.585 1996.970 719.170 1996.980 ;
        RECT 718.360 1996.670 719.170 1996.970 ;
        RECT 718.585 1996.660 719.170 1996.670 ;
        RECT 718.585 1996.655 718.915 1996.660 ;
        RECT 713.985 1956.850 714.315 1956.865 ;
        RECT 718.790 1956.850 719.170 1956.860 ;
        RECT 713.985 1956.550 719.170 1956.850 ;
        RECT 713.985 1956.535 714.315 1956.550 ;
        RECT 718.790 1956.540 719.170 1956.550 ;
        RECT 713.065 1946.650 713.395 1946.665 ;
        RECT 718.790 1946.650 719.170 1946.660 ;
        RECT 713.065 1946.350 719.170 1946.650 ;
        RECT 713.065 1946.335 713.395 1946.350 ;
        RECT 718.790 1946.340 719.170 1946.350 ;
        RECT 716.030 1926.930 716.410 1926.940 ;
        RECT 718.790 1926.930 719.170 1926.940 ;
        RECT 716.030 1926.630 719.170 1926.930 ;
        RECT 716.030 1926.620 716.410 1926.630 ;
        RECT 718.790 1926.620 719.170 1926.630 ;
        RECT 713.525 1924.890 713.855 1924.905 ;
        RECT 718.790 1924.890 719.170 1924.900 ;
        RECT 713.525 1924.590 719.170 1924.890 ;
        RECT 713.525 1924.575 713.855 1924.590 ;
        RECT 718.790 1924.580 719.170 1924.590 ;
        RECT 713.065 1922.170 713.395 1922.185 ;
        RECT 718.790 1922.170 719.170 1922.180 ;
        RECT 713.065 1921.870 719.170 1922.170 ;
        RECT 713.065 1921.855 713.395 1921.870 ;
        RECT 718.790 1921.860 719.170 1921.870 ;
        RECT 716.950 1912.650 717.330 1912.660 ;
        RECT 718.790 1912.650 719.170 1912.660 ;
        RECT 716.950 1912.350 719.170 1912.650 ;
        RECT 716.950 1912.340 717.330 1912.350 ;
        RECT 718.790 1912.340 719.170 1912.350 ;
        RECT 713.065 1911.970 713.395 1911.985 ;
        RECT 716.030 1911.970 716.410 1911.980 ;
        RECT 713.065 1911.670 716.410 1911.970 ;
        RECT 713.065 1911.655 713.395 1911.670 ;
        RECT 716.030 1911.660 716.410 1911.670 ;
        RECT 717.665 1909.250 717.995 1909.265 ;
        RECT 718.790 1909.250 719.170 1909.260 ;
        RECT 717.665 1908.950 719.170 1909.250 ;
        RECT 717.665 1908.935 717.995 1908.950 ;
        RECT 718.790 1908.940 719.170 1908.950 ;
        RECT 716.950 1907.210 717.330 1907.220 ;
        RECT 712.390 1906.910 717.330 1907.210 ;
        RECT 712.390 1905.850 712.690 1906.910 ;
        RECT 716.950 1906.900 717.330 1906.910 ;
        RECT 713.065 1906.530 713.395 1906.545 ;
        RECT 718.790 1906.530 719.170 1906.540 ;
        RECT 713.065 1906.230 719.170 1906.530 ;
        RECT 713.065 1906.215 713.395 1906.230 ;
        RECT 718.790 1906.220 719.170 1906.230 ;
        RECT 713.065 1905.850 713.395 1905.865 ;
        RECT 712.390 1905.550 713.395 1905.850 ;
        RECT 713.065 1905.535 713.395 1905.550 ;
        RECT 713.525 1820.850 713.855 1820.865 ;
        RECT 718.790 1820.850 719.170 1820.860 ;
        RECT 713.525 1820.550 719.170 1820.850 ;
        RECT 713.525 1820.535 713.855 1820.550 ;
        RECT 718.790 1820.540 719.170 1820.550 ;
        RECT 713.525 1777.330 713.855 1777.345 ;
        RECT 718.790 1777.330 719.170 1777.340 ;
        RECT 713.525 1777.030 719.170 1777.330 ;
        RECT 713.525 1777.015 713.855 1777.030 ;
        RECT 718.790 1777.020 719.170 1777.030 ;
        RECT 714.190 1742.650 714.570 1742.660 ;
        RECT 718.790 1742.650 719.170 1742.660 ;
        RECT 714.190 1742.350 719.170 1742.650 ;
        RECT 714.190 1742.340 714.570 1742.350 ;
        RECT 718.790 1742.340 719.170 1742.350 ;
        RECT 713.065 1739.250 713.395 1739.265 ;
        RECT 718.790 1739.250 719.170 1739.260 ;
        RECT 713.065 1738.950 719.170 1739.250 ;
        RECT 713.065 1738.935 713.395 1738.950 ;
        RECT 718.790 1738.940 719.170 1738.950 ;
        RECT 712.350 1731.770 712.730 1731.780 ;
        RECT 714.190 1731.770 714.570 1731.780 ;
        RECT 712.350 1731.470 714.570 1731.770 ;
        RECT 712.350 1731.460 712.730 1731.470 ;
        RECT 714.190 1731.460 714.570 1731.470 ;
        RECT 710.305 1721.570 710.635 1721.585 ;
        RECT 718.790 1721.570 719.170 1721.580 ;
        RECT 710.305 1721.270 719.170 1721.570 ;
        RECT 710.305 1721.255 710.635 1721.270 ;
        RECT 718.790 1721.260 719.170 1721.270 ;
        RECT 710.305 1718.850 710.635 1718.865 ;
        RECT 718.790 1718.850 719.170 1718.860 ;
        RECT 710.305 1718.550 719.170 1718.850 ;
        RECT 710.305 1718.535 710.635 1718.550 ;
        RECT 718.790 1718.540 719.170 1718.550 ;
        RECT 712.350 1698.450 712.730 1698.460 ;
        RECT 718.790 1698.450 719.170 1698.460 ;
        RECT 712.350 1698.150 719.170 1698.450 ;
        RECT 712.350 1698.140 712.730 1698.150 ;
        RECT 718.790 1698.140 719.170 1698.150 ;
        RECT 712.145 1681.450 712.475 1681.465 ;
        RECT 718.790 1681.450 719.170 1681.460 ;
        RECT 712.145 1681.150 719.170 1681.450 ;
        RECT 712.145 1681.135 712.475 1681.150 ;
        RECT 718.790 1681.140 719.170 1681.150 ;
        RECT 713.065 1671.250 713.395 1671.265 ;
        RECT 718.790 1671.250 719.170 1671.260 ;
        RECT 713.065 1670.950 719.170 1671.250 ;
        RECT 713.065 1670.935 713.395 1670.950 ;
        RECT 718.790 1670.940 719.170 1670.950 ;
        RECT 714.190 1665.130 714.570 1665.140 ;
        RECT 718.790 1665.130 719.170 1665.140 ;
        RECT 714.190 1664.830 719.170 1665.130 ;
        RECT 714.190 1664.820 714.570 1664.830 ;
        RECT 718.790 1664.820 719.170 1664.830 ;
        RECT 717.205 1664.450 717.535 1664.465 ;
        RECT 718.790 1664.450 719.170 1664.460 ;
        RECT 717.205 1664.150 719.170 1664.450 ;
        RECT 717.205 1664.135 717.535 1664.150 ;
        RECT 718.790 1664.140 719.170 1664.150 ;
        RECT 712.145 1662.410 712.475 1662.425 ;
        RECT 718.790 1662.410 719.170 1662.420 ;
        RECT 712.145 1662.110 719.170 1662.410 ;
        RECT 712.145 1662.095 712.475 1662.110 ;
        RECT 718.790 1662.100 719.170 1662.110 ;
        RECT 718.790 1654.930 719.170 1654.940 ;
        RECT 713.540 1654.630 719.170 1654.930 ;
        RECT 713.540 1652.905 713.840 1654.630 ;
        RECT 718.790 1654.620 719.170 1654.630 ;
        RECT 714.190 1654.250 714.570 1654.260 ;
        RECT 718.790 1654.250 719.170 1654.260 ;
        RECT 714.190 1653.950 719.170 1654.250 ;
        RECT 714.190 1653.940 714.570 1653.950 ;
        RECT 718.790 1653.940 719.170 1653.950 ;
        RECT 713.525 1652.575 713.855 1652.905 ;
        RECT 713.525 1638.610 713.855 1638.625 ;
        RECT 718.790 1638.610 719.170 1638.620 ;
        RECT 713.525 1638.310 719.170 1638.610 ;
        RECT 713.525 1638.295 713.855 1638.310 ;
        RECT 718.790 1638.300 719.170 1638.310 ;
        RECT 713.985 1637.930 714.315 1637.945 ;
        RECT 718.790 1637.930 719.170 1637.940 ;
        RECT 713.985 1637.630 719.170 1637.930 ;
        RECT 713.985 1637.615 714.315 1637.630 ;
        RECT 718.790 1637.620 719.170 1637.630 ;
        RECT 713.525 1631.810 713.855 1631.825 ;
        RECT 718.790 1631.810 719.170 1631.820 ;
        RECT 713.525 1631.510 719.170 1631.810 ;
        RECT 713.525 1631.495 713.855 1631.510 ;
        RECT 718.790 1631.500 719.170 1631.510 ;
        RECT 728.910 1326.490 729.290 1326.500 ;
        RECT 730.545 1326.490 730.875 1326.505 ;
        RECT 728.910 1326.190 730.875 1326.490 ;
        RECT 728.910 1326.180 729.290 1326.190 ;
        RECT 730.545 1326.175 730.875 1326.190 ;
        RECT 731.670 1326.490 732.050 1326.500 ;
        RECT 1008.845 1326.490 1009.175 1326.505 ;
        RECT 1148.225 1326.500 1148.555 1326.505 ;
        RECT 1148.225 1326.490 1148.810 1326.500 ;
        RECT 731.670 1326.190 1009.175 1326.490 ;
        RECT 1148.000 1326.190 1148.810 1326.490 ;
        RECT 731.670 1326.180 732.050 1326.190 ;
        RECT 1008.845 1326.175 1009.175 1326.190 ;
        RECT 1148.225 1326.180 1148.810 1326.190 ;
        RECT 1148.225 1326.175 1148.555 1326.180 ;
        RECT 725.230 1325.810 725.610 1325.820 ;
        RECT 729.830 1325.810 730.210 1325.820 ;
        RECT 725.230 1325.510 730.210 1325.810 ;
        RECT 725.230 1325.500 725.610 1325.510 ;
        RECT 729.830 1325.500 730.210 1325.510 ;
        RECT 730.750 1325.810 731.130 1325.820 ;
        RECT 898.445 1325.810 898.775 1325.825 ;
        RECT 730.750 1325.510 898.775 1325.810 ;
        RECT 730.750 1325.500 731.130 1325.510 ;
        RECT 898.445 1325.495 898.775 1325.510 ;
        RECT 730.750 1324.450 731.130 1324.460 ;
        RECT 735.350 1324.450 735.730 1324.460 ;
        RECT 730.750 1324.150 735.730 1324.450 ;
        RECT 730.750 1324.140 731.130 1324.150 ;
        RECT 735.350 1324.140 735.730 1324.150 ;
        RECT 932.230 1297.930 932.610 1297.940 ;
        RECT 953.390 1297.930 953.770 1297.940 ;
        RECT 932.230 1297.630 953.770 1297.930 ;
        RECT 932.230 1297.620 932.610 1297.630 ;
        RECT 953.390 1297.620 953.770 1297.630 ;
        RECT 953.390 1202.050 953.770 1202.060 ;
        RECT 952.510 1201.750 953.770 1202.050 ;
        RECT 952.510 1201.380 952.810 1201.750 ;
        RECT 953.390 1201.740 953.770 1201.750 ;
        RECT 952.470 1201.060 952.850 1201.380 ;
        RECT 952.470 1173.180 952.850 1173.500 ;
        RECT 952.510 1172.130 952.810 1173.180 ;
        RECT 953.390 1172.130 953.770 1172.140 ;
        RECT 952.510 1171.830 953.770 1172.130 ;
        RECT 953.390 1171.820 953.770 1171.830 ;
        RECT 953.645 1159.220 953.975 1159.225 ;
        RECT 953.390 1159.210 953.975 1159.220 ;
        RECT 953.190 1158.910 953.975 1159.210 ;
        RECT 953.390 1158.900 953.975 1158.910 ;
        RECT 953.645 1158.895 953.975 1158.900 ;
        RECT 953.645 1111.610 953.975 1111.625 ;
        RECT 954.310 1111.610 954.690 1111.620 ;
        RECT 953.645 1111.310 954.690 1111.610 ;
        RECT 953.645 1111.295 953.975 1111.310 ;
        RECT 954.310 1111.300 954.690 1111.310 ;
        RECT 954.310 1077.610 954.690 1077.620 ;
        RECT 953.430 1077.310 954.690 1077.610 ;
        RECT 953.430 1076.260 953.730 1077.310 ;
        RECT 954.310 1077.300 954.690 1077.310 ;
        RECT 953.390 1075.940 953.770 1076.260 ;
        RECT 953.645 1062.660 953.975 1062.665 ;
        RECT 953.390 1062.650 953.975 1062.660 ;
        RECT 953.190 1062.350 953.975 1062.650 ;
        RECT 953.390 1062.340 953.975 1062.350 ;
        RECT 953.645 1062.335 953.975 1062.340 ;
        RECT 953.645 1015.050 953.975 1015.065 ;
        RECT 954.310 1015.050 954.690 1015.060 ;
        RECT 953.645 1014.750 954.690 1015.050 ;
        RECT 953.645 1014.735 953.975 1014.750 ;
        RECT 954.310 1014.740 954.690 1014.750 ;
        RECT 954.310 981.050 954.690 981.060 ;
        RECT 953.430 980.750 954.690 981.050 ;
        RECT 953.430 979.020 953.730 980.750 ;
        RECT 954.310 980.740 954.690 980.750 ;
        RECT 953.390 978.700 953.770 979.020 ;
        RECT 952.725 966.090 953.055 966.105 ;
        RECT 953.390 966.090 953.770 966.100 ;
        RECT 952.725 965.790 953.770 966.090 ;
        RECT 952.725 965.775 953.055 965.790 ;
        RECT 953.390 965.780 953.770 965.790 ;
        RECT 952.725 919.170 953.055 919.185 ;
        RECT 952.510 918.855 953.055 919.170 ;
        RECT 952.510 918.500 952.810 918.855 ;
        RECT 952.470 918.180 952.850 918.500 ;
        RECT 952.470 883.500 952.850 883.820 ;
        RECT 952.510 882.450 952.810 883.500 ;
        RECT 953.390 882.450 953.770 882.460 ;
        RECT 952.510 882.150 953.770 882.450 ;
        RECT 953.390 882.140 953.770 882.150 ;
        RECT 952.725 869.530 953.055 869.545 ;
        RECT 953.390 869.530 953.770 869.540 ;
        RECT 952.725 869.230 953.770 869.530 ;
        RECT 952.725 869.215 953.055 869.230 ;
        RECT 953.390 869.220 953.770 869.230 ;
        RECT 952.725 821.260 953.055 821.265 ;
        RECT 952.470 821.250 953.055 821.260 ;
        RECT 952.270 820.950 953.055 821.250 ;
        RECT 952.470 820.940 953.055 820.950 ;
        RECT 952.725 820.935 953.055 820.940 ;
        RECT 952.470 786.940 952.850 787.260 ;
        RECT 952.510 785.890 952.810 786.940 ;
        RECT 953.390 785.890 953.770 785.900 ;
        RECT 952.510 785.590 953.770 785.890 ;
        RECT 953.390 785.580 953.770 785.590 ;
        RECT 953.645 772.300 953.975 772.305 ;
        RECT 953.390 772.290 953.975 772.300 ;
        RECT 953.390 771.990 954.200 772.290 ;
        RECT 953.390 771.980 953.975 771.990 ;
        RECT 953.645 771.975 953.975 771.980 ;
        RECT 952.470 724.690 952.850 724.700 ;
        RECT 953.645 724.690 953.975 724.705 ;
        RECT 952.470 724.390 953.975 724.690 ;
        RECT 952.470 724.380 952.850 724.390 ;
        RECT 953.645 724.375 953.975 724.390 ;
        RECT 952.470 690.380 952.850 690.700 ;
        RECT 952.510 689.330 952.810 690.380 ;
        RECT 953.390 689.330 953.770 689.340 ;
        RECT 952.510 689.030 953.770 689.330 ;
        RECT 953.390 689.020 953.770 689.030 ;
        RECT 953.390 675.420 953.770 675.740 ;
        RECT 953.430 675.065 953.730 675.420 ;
        RECT 953.430 674.750 953.975 675.065 ;
        RECT 953.645 674.735 953.975 674.750 ;
        RECT 953.645 628.130 953.975 628.145 ;
        RECT 954.310 628.130 954.690 628.140 ;
        RECT 953.645 627.830 954.690 628.130 ;
        RECT 953.645 627.815 953.975 627.830 ;
        RECT 954.310 627.820 954.690 627.830 ;
        RECT 954.310 594.130 954.690 594.140 ;
        RECT 953.430 593.830 954.690 594.130 ;
        RECT 953.430 592.780 953.730 593.830 ;
        RECT 954.310 593.820 954.690 593.830 ;
        RECT 953.390 592.460 953.770 592.780 ;
        RECT 953.390 545.540 953.770 545.860 ;
        RECT 953.430 544.490 953.730 545.540 ;
        RECT 954.310 544.490 954.690 544.500 ;
        RECT 953.430 544.190 954.690 544.490 ;
        RECT 954.310 544.180 954.690 544.190 ;
        RECT 954.310 497.570 954.690 497.580 ;
        RECT 953.430 497.270 954.690 497.570 ;
        RECT 953.430 496.220 953.730 497.270 ;
        RECT 954.310 497.260 954.690 497.270 ;
        RECT 953.390 495.900 953.770 496.220 ;
        RECT 953.390 449.290 953.770 449.300 ;
        RECT 952.510 448.990 953.770 449.290 ;
        RECT 952.510 447.940 952.810 448.990 ;
        RECT 953.390 448.980 953.770 448.990 ;
        RECT 952.470 447.620 952.850 447.940 ;
        RECT 952.470 427.220 952.850 427.540 ;
        RECT 952.510 426.865 952.810 427.220 ;
        RECT 952.510 426.550 953.055 426.865 ;
        RECT 952.725 426.535 953.055 426.550 ;
        RECT 952.725 380.610 953.055 380.625 ;
        RECT 953.390 380.610 953.770 380.620 ;
        RECT 952.725 380.310 953.770 380.610 ;
        RECT 952.725 380.295 953.055 380.310 ;
        RECT 953.390 380.300 953.770 380.310 ;
        RECT 952.470 304.140 952.850 304.460 ;
        RECT 952.510 303.090 952.810 304.140 ;
        RECT 953.390 303.090 953.770 303.100 ;
        RECT 952.510 302.790 953.770 303.090 ;
        RECT 953.390 302.780 953.770 302.790 ;
        RECT 953.390 289.180 953.770 289.500 ;
        RECT 953.430 288.825 953.730 289.180 ;
        RECT 953.430 288.510 953.975 288.825 ;
        RECT 953.645 288.495 953.975 288.510 ;
        RECT 953.645 241.890 953.975 241.905 ;
        RECT 954.310 241.890 954.690 241.900 ;
        RECT 953.645 241.590 954.690 241.890 ;
        RECT 953.645 241.575 953.975 241.590 ;
        RECT 954.310 241.580 954.690 241.590 ;
        RECT 954.310 207.890 954.690 207.900 ;
        RECT 953.430 207.590 954.690 207.890 ;
        RECT 953.430 206.540 953.730 207.590 ;
        RECT 954.310 207.580 954.690 207.590 ;
        RECT 953.390 206.220 953.770 206.540 ;
        RECT 952.725 192.930 953.055 192.945 ;
        RECT 953.390 192.930 953.770 192.940 ;
        RECT 952.725 192.630 953.770 192.930 ;
        RECT 952.725 192.615 953.055 192.630 ;
        RECT 953.390 192.620 953.770 192.630 ;
        RECT 952.725 146.010 953.055 146.025 ;
        RECT 952.510 145.695 953.055 146.010 ;
        RECT 952.510 145.340 952.810 145.695 ;
        RECT 952.470 145.020 952.850 145.340 ;
        RECT 953.390 96.060 953.770 96.380 ;
        RECT 953.430 95.705 953.730 96.060 ;
        RECT 953.430 95.390 953.975 95.705 ;
        RECT 953.645 95.375 953.975 95.390 ;
        RECT 953.645 48.770 953.975 48.785 ;
        RECT 954.310 48.770 954.690 48.780 ;
        RECT 953.645 48.470 954.690 48.770 ;
        RECT 953.645 48.455 953.975 48.470 ;
        RECT 954.310 48.460 954.690 48.470 ;
        RECT 954.105 24.980 954.435 24.985 ;
        RECT 954.105 24.970 954.690 24.980 ;
        RECT 953.880 24.670 954.690 24.970 ;
        RECT 954.105 24.660 954.690 24.670 ;
        RECT 954.105 24.655 954.435 24.660 ;
        RECT 1148.430 18.850 1148.810 18.860 ;
        RECT 1150.525 18.850 1150.855 18.865 ;
        RECT 1148.430 18.550 1150.855 18.850 ;
        RECT 1148.430 18.540 1148.810 18.550 ;
        RECT 1150.525 18.535 1150.855 18.550 ;
        RECT 1035.270 14.770 1035.650 14.780 ;
        RECT 1037.365 14.770 1037.695 14.785 ;
        RECT 1035.270 14.470 1037.695 14.770 ;
        RECT 1035.270 14.460 1035.650 14.470 ;
        RECT 1037.365 14.455 1037.695 14.470 ;
      LAYER via3 ;
        RECT 730.780 2393.100 731.100 2393.420 ;
        RECT 729.860 2391.740 730.180 2392.060 ;
        RECT 738.140 2374.740 738.460 2375.060 ;
        RECT 739.060 2374.060 739.380 2374.380 ;
        RECT 1303.940 2374.060 1304.260 2374.380 ;
        RECT 723.420 2369.980 723.740 2370.300 ;
        RECT 1303.940 2369.980 1304.260 2370.300 ;
        RECT 726.180 2366.580 726.500 2366.900 ;
        RECT 739.060 2366.580 739.380 2366.900 ;
        RECT 725.260 2365.900 725.580 2366.220 ;
        RECT 738.140 2365.900 738.460 2366.220 ;
        RECT 718.820 2218.340 719.140 2218.660 ;
        RECT 717.900 2200.660 718.220 2200.980 ;
        RECT 718.820 2195.220 719.140 2195.540 ;
        RECT 718.820 2194.540 719.140 2194.860 ;
        RECT 718.820 2187.740 719.140 2188.060 ;
        RECT 718.820 2187.060 719.140 2187.380 ;
        RECT 718.820 2183.660 719.140 2183.980 ;
        RECT 718.820 2180.260 719.140 2180.580 ;
        RECT 718.820 2000.740 719.140 2001.060 ;
        RECT 718.820 1997.340 719.140 1997.660 ;
        RECT 718.820 1996.660 719.140 1996.980 ;
        RECT 718.820 1956.540 719.140 1956.860 ;
        RECT 718.820 1946.340 719.140 1946.660 ;
        RECT 716.060 1926.620 716.380 1926.940 ;
        RECT 718.820 1926.620 719.140 1926.940 ;
        RECT 718.820 1924.580 719.140 1924.900 ;
        RECT 718.820 1921.860 719.140 1922.180 ;
        RECT 716.980 1912.340 717.300 1912.660 ;
        RECT 718.820 1912.340 719.140 1912.660 ;
        RECT 716.060 1911.660 716.380 1911.980 ;
        RECT 718.820 1908.940 719.140 1909.260 ;
        RECT 716.980 1906.900 717.300 1907.220 ;
        RECT 718.820 1906.220 719.140 1906.540 ;
        RECT 718.820 1820.540 719.140 1820.860 ;
        RECT 718.820 1777.020 719.140 1777.340 ;
        RECT 714.220 1742.340 714.540 1742.660 ;
        RECT 718.820 1742.340 719.140 1742.660 ;
        RECT 718.820 1738.940 719.140 1739.260 ;
        RECT 712.380 1731.460 712.700 1731.780 ;
        RECT 714.220 1731.460 714.540 1731.780 ;
        RECT 718.820 1721.260 719.140 1721.580 ;
        RECT 718.820 1718.540 719.140 1718.860 ;
        RECT 712.380 1698.140 712.700 1698.460 ;
        RECT 718.820 1698.140 719.140 1698.460 ;
        RECT 718.820 1681.140 719.140 1681.460 ;
        RECT 718.820 1670.940 719.140 1671.260 ;
        RECT 714.220 1664.820 714.540 1665.140 ;
        RECT 718.820 1664.820 719.140 1665.140 ;
        RECT 718.820 1664.140 719.140 1664.460 ;
        RECT 718.820 1662.100 719.140 1662.420 ;
        RECT 718.820 1654.620 719.140 1654.940 ;
        RECT 714.220 1653.940 714.540 1654.260 ;
        RECT 718.820 1653.940 719.140 1654.260 ;
        RECT 718.820 1638.300 719.140 1638.620 ;
        RECT 718.820 1637.620 719.140 1637.940 ;
        RECT 718.820 1631.500 719.140 1631.820 ;
        RECT 728.940 1326.180 729.260 1326.500 ;
        RECT 731.700 1326.180 732.020 1326.500 ;
        RECT 1148.460 1326.180 1148.780 1326.500 ;
        RECT 725.260 1325.500 725.580 1325.820 ;
        RECT 729.860 1325.500 730.180 1325.820 ;
        RECT 730.780 1325.500 731.100 1325.820 ;
        RECT 730.780 1324.140 731.100 1324.460 ;
        RECT 735.380 1324.140 735.700 1324.460 ;
        RECT 932.260 1297.620 932.580 1297.940 ;
        RECT 953.420 1297.620 953.740 1297.940 ;
        RECT 953.420 1201.740 953.740 1202.060 ;
        RECT 952.500 1201.060 952.820 1201.380 ;
        RECT 952.500 1173.180 952.820 1173.500 ;
        RECT 953.420 1171.820 953.740 1172.140 ;
        RECT 953.420 1158.900 953.740 1159.220 ;
        RECT 954.340 1111.300 954.660 1111.620 ;
        RECT 954.340 1077.300 954.660 1077.620 ;
        RECT 953.420 1075.940 953.740 1076.260 ;
        RECT 953.420 1062.340 953.740 1062.660 ;
        RECT 954.340 1014.740 954.660 1015.060 ;
        RECT 954.340 980.740 954.660 981.060 ;
        RECT 953.420 978.700 953.740 979.020 ;
        RECT 953.420 965.780 953.740 966.100 ;
        RECT 952.500 918.180 952.820 918.500 ;
        RECT 952.500 883.500 952.820 883.820 ;
        RECT 953.420 882.140 953.740 882.460 ;
        RECT 953.420 869.220 953.740 869.540 ;
        RECT 952.500 820.940 952.820 821.260 ;
        RECT 952.500 786.940 952.820 787.260 ;
        RECT 953.420 785.580 953.740 785.900 ;
        RECT 953.420 771.980 953.740 772.300 ;
        RECT 952.500 724.380 952.820 724.700 ;
        RECT 952.500 690.380 952.820 690.700 ;
        RECT 953.420 689.020 953.740 689.340 ;
        RECT 953.420 675.420 953.740 675.740 ;
        RECT 954.340 627.820 954.660 628.140 ;
        RECT 954.340 593.820 954.660 594.140 ;
        RECT 953.420 592.460 953.740 592.780 ;
        RECT 953.420 545.540 953.740 545.860 ;
        RECT 954.340 544.180 954.660 544.500 ;
        RECT 954.340 497.260 954.660 497.580 ;
        RECT 953.420 495.900 953.740 496.220 ;
        RECT 953.420 448.980 953.740 449.300 ;
        RECT 952.500 447.620 952.820 447.940 ;
        RECT 952.500 427.220 952.820 427.540 ;
        RECT 953.420 380.300 953.740 380.620 ;
        RECT 952.500 304.140 952.820 304.460 ;
        RECT 953.420 302.780 953.740 303.100 ;
        RECT 953.420 289.180 953.740 289.500 ;
        RECT 954.340 241.580 954.660 241.900 ;
        RECT 954.340 207.580 954.660 207.900 ;
        RECT 953.420 206.220 953.740 206.540 ;
        RECT 953.420 192.620 953.740 192.940 ;
        RECT 952.500 145.020 952.820 145.340 ;
        RECT 953.420 96.060 953.740 96.380 ;
        RECT 954.340 48.460 954.660 48.780 ;
        RECT 954.340 24.660 954.660 24.980 ;
        RECT 1148.460 18.540 1148.780 18.860 ;
        RECT 1035.300 14.460 1035.620 14.780 ;
      LAYER met4 ;
        RECT 730.775 2393.095 731.105 2393.425 ;
        RECT 729.855 2391.735 730.185 2392.065 ;
        RECT 723.415 2369.975 723.745 2370.305 ;
        RECT 723.430 2355.090 723.730 2369.975 ;
        RECT 726.175 2366.575 726.505 2366.905 ;
        RECT 725.255 2365.895 725.585 2366.225 ;
        RECT 722.990 2353.910 724.170 2355.090 ;
        RECT 725.270 2320.650 725.570 2365.895 ;
        RECT 724.350 2320.350 725.570 2320.650 ;
        RECT 724.350 2314.530 724.650 2320.350 ;
        RECT 726.190 2317.250 726.490 2366.575 ;
        RECT 727.590 2350.510 728.770 2351.690 ;
        RECT 728.030 2344.450 728.330 2350.510 ;
        RECT 728.030 2344.150 729.250 2344.450 ;
        RECT 726.190 2316.950 727.410 2317.250 ;
        RECT 724.350 2314.230 725.570 2314.530 ;
        RECT 725.270 2266.250 725.570 2314.230 ;
        RECT 724.350 2265.950 725.570 2266.250 ;
        RECT 718.815 2218.650 719.145 2218.665 ;
        RECT 724.350 2218.650 724.650 2265.950 ;
        RECT 727.110 2259.450 727.410 2316.950 ;
        RECT 718.815 2218.350 724.650 2218.650 ;
        RECT 725.270 2259.150 727.410 2259.450 ;
        RECT 718.815 2218.335 719.145 2218.350 ;
        RECT 725.270 2208.450 725.570 2259.150 ;
        RECT 728.950 2249.250 729.250 2344.150 ;
        RECT 718.830 2208.150 725.570 2208.450 ;
        RECT 726.190 2248.950 729.250 2249.250 ;
        RECT 717.895 2200.655 718.225 2200.985 ;
        RECT 717.910 2164.250 718.210 2200.655 ;
        RECT 718.830 2195.545 719.130 2208.150 ;
        RECT 718.815 2195.215 719.145 2195.545 ;
        RECT 718.815 2194.850 719.145 2194.865 ;
        RECT 726.190 2194.850 726.490 2248.950 ;
        RECT 729.870 2243.130 730.170 2391.735 ;
        RECT 730.790 2351.250 731.090 2393.095 ;
        RECT 738.135 2374.735 738.465 2375.065 ;
        RECT 738.150 2366.225 738.450 2374.735 ;
        RECT 739.055 2374.055 739.385 2374.385 ;
        RECT 1303.935 2374.055 1304.265 2374.385 ;
        RECT 739.070 2366.905 739.370 2374.055 ;
        RECT 1303.950 2370.305 1304.250 2374.055 ;
        RECT 1303.935 2369.975 1304.265 2370.305 ;
        RECT 739.055 2366.575 739.385 2366.905 ;
        RECT 738.135 2365.895 738.465 2366.225 ;
        RECT 730.790 2350.950 732.010 2351.250 ;
        RECT 731.710 2262.850 732.010 2350.950 ;
        RECT 718.815 2194.550 726.490 2194.850 ;
        RECT 728.950 2242.830 730.170 2243.130 ;
        RECT 730.790 2262.550 732.010 2262.850 ;
        RECT 718.815 2194.535 719.145 2194.550 ;
        RECT 728.950 2188.730 729.250 2242.830 ;
        RECT 730.790 2225.450 731.090 2262.550 ;
        RECT 718.830 2188.430 729.250 2188.730 ;
        RECT 729.870 2225.150 731.090 2225.450 ;
        RECT 718.830 2188.065 719.130 2188.430 ;
        RECT 718.815 2187.735 719.145 2188.065 ;
        RECT 729.870 2188.050 730.170 2225.150 ;
        RECT 729.870 2187.750 732.010 2188.050 ;
        RECT 718.815 2187.370 719.145 2187.385 ;
        RECT 718.815 2187.070 728.330 2187.370 ;
        RECT 718.815 2187.055 719.145 2187.070 ;
        RECT 718.815 2183.655 719.145 2183.985 ;
        RECT 718.830 2181.930 719.130 2183.655 ;
        RECT 718.830 2181.630 727.410 2181.930 ;
        RECT 718.815 2180.255 719.145 2180.585 ;
        RECT 718.830 2174.450 719.130 2180.255 ;
        RECT 718.830 2174.150 722.810 2174.450 ;
        RECT 717.910 2163.950 719.130 2164.250 ;
        RECT 718.830 2162.210 719.130 2163.950 ;
        RECT 718.830 2161.910 720.970 2162.210 ;
        RECT 720.670 2147.250 720.970 2161.910 ;
        RECT 720.670 2146.950 721.890 2147.250 ;
        RECT 721.590 2143.850 721.890 2146.950 ;
        RECT 719.750 2143.550 721.890 2143.850 ;
        RECT 722.510 2143.850 722.810 2174.150 ;
        RECT 722.510 2143.550 723.730 2143.850 ;
        RECT 719.750 2096.250 720.050 2143.550 ;
        RECT 723.430 2130.250 723.730 2143.550 ;
        RECT 727.110 2133.650 727.410 2181.630 ;
        RECT 721.590 2129.950 723.730 2130.250 ;
        RECT 724.350 2133.350 727.410 2133.650 ;
        RECT 721.590 2099.650 721.890 2129.950 ;
        RECT 724.350 2126.850 724.650 2133.350 ;
        RECT 722.510 2126.550 724.650 2126.850 ;
        RECT 722.510 2116.650 722.810 2126.550 ;
        RECT 722.510 2116.350 723.730 2116.650 ;
        RECT 723.430 2109.850 723.730 2116.350 ;
        RECT 728.030 2109.850 728.330 2187.070 ;
        RECT 731.710 2137.050 732.010 2187.750 ;
        RECT 729.870 2136.750 732.010 2137.050 ;
        RECT 729.870 2130.250 730.170 2136.750 ;
        RECT 729.870 2129.950 732.010 2130.250 ;
        RECT 731.710 2126.850 732.010 2129.950 ;
        RECT 730.790 2126.550 732.010 2126.850 ;
        RECT 723.430 2109.550 725.570 2109.850 ;
        RECT 728.030 2109.550 730.170 2109.850 ;
        RECT 725.270 2106.450 725.570 2109.550 ;
        RECT 725.270 2106.150 728.330 2106.450 ;
        RECT 721.590 2099.350 724.650 2099.650 ;
        RECT 719.750 2095.950 723.730 2096.250 ;
        RECT 723.430 2052.730 723.730 2095.950 ;
        RECT 724.350 2073.810 724.650 2099.350 ;
        RECT 728.030 2073.810 728.330 2106.150 ;
        RECT 724.350 2073.510 725.570 2073.810 ;
        RECT 725.270 2071.770 725.570 2073.510 ;
        RECT 724.350 2071.470 725.570 2071.770 ;
        RECT 727.110 2073.510 728.330 2073.810 ;
        RECT 724.350 2065.650 724.650 2071.470 ;
        RECT 724.350 2065.350 726.490 2065.650 ;
        RECT 726.190 2055.450 726.490 2065.350 ;
        RECT 727.110 2062.250 727.410 2073.510 ;
        RECT 727.110 2061.950 729.250 2062.250 ;
        RECT 726.190 2055.150 728.330 2055.450 ;
        RECT 720.670 2052.430 723.730 2052.730 ;
        RECT 720.670 2048.650 720.970 2052.430 ;
        RECT 728.030 2048.650 728.330 2055.150 ;
        RECT 728.950 2048.650 729.250 2061.950 ;
        RECT 729.870 2052.050 730.170 2109.550 ;
        RECT 730.790 2052.050 731.090 2126.550 ;
        RECT 729.870 2051.750 732.010 2052.050 ;
        RECT 719.750 2048.350 720.970 2048.650 ;
        RECT 722.510 2048.350 729.250 2048.650 ;
        RECT 718.815 2001.050 719.145 2001.065 ;
        RECT 719.750 2001.050 720.050 2048.350 ;
        RECT 722.510 2045.250 722.810 2048.350 ;
        RECT 728.030 2045.250 728.330 2048.350 ;
        RECT 730.790 2045.250 731.090 2051.750 ;
        RECT 720.670 2044.950 731.090 2045.250 ;
        RECT 720.670 2028.250 720.970 2044.950 ;
        RECT 722.510 2038.450 722.810 2044.950 ;
        RECT 721.590 2038.150 722.810 2038.450 ;
        RECT 721.590 2034.370 721.890 2038.150 ;
        RECT 721.590 2034.070 725.570 2034.370 ;
        RECT 725.270 2028.250 725.570 2034.070 ;
        RECT 720.670 2027.950 723.730 2028.250 ;
        RECT 723.430 2001.050 723.730 2027.950 ;
        RECT 724.350 2027.950 725.570 2028.250 ;
        RECT 724.350 2014.650 724.650 2027.950 ;
        RECT 728.030 2014.650 728.330 2044.950 ;
        RECT 724.350 2014.350 729.250 2014.650 ;
        RECT 728.030 2011.250 728.330 2014.350 ;
        RECT 718.815 2000.750 720.050 2001.050 ;
        RECT 720.670 2000.750 723.730 2001.050 ;
        RECT 724.350 2010.950 728.330 2011.250 ;
        RECT 718.815 2000.735 719.145 2000.750 ;
        RECT 718.815 1997.650 719.145 1997.665 ;
        RECT 720.670 1997.650 720.970 2000.750 ;
        RECT 718.815 1997.350 720.970 1997.650 ;
        RECT 718.815 1997.335 719.145 1997.350 ;
        RECT 718.815 1996.655 719.145 1996.985 ;
        RECT 724.350 1996.970 724.650 2010.950 ;
        RECT 728.950 2001.050 729.250 2014.350 ;
        RECT 728.030 2000.750 729.250 2001.050 ;
        RECT 724.350 1996.670 726.490 1996.970 ;
        RECT 718.830 1994.250 719.130 1996.655 ;
        RECT 718.830 1993.950 723.730 1994.250 ;
        RECT 723.430 1967.050 723.730 1993.950 ;
        RECT 726.190 1990.850 726.490 1996.670 ;
        RECT 721.590 1966.750 723.730 1967.050 ;
        RECT 724.350 1990.550 726.490 1990.850 ;
        RECT 721.590 1964.330 721.890 1966.750 ;
        RECT 720.670 1964.030 721.890 1964.330 ;
        RECT 718.815 1956.850 719.145 1956.865 ;
        RECT 718.815 1956.550 720.050 1956.850 ;
        RECT 718.815 1956.535 719.145 1956.550 ;
        RECT 718.815 1946.650 719.145 1946.665 ;
        RECT 719.750 1946.650 720.050 1956.550 ;
        RECT 718.815 1946.350 720.050 1946.650 ;
        RECT 718.815 1946.335 719.145 1946.350 ;
        RECT 720.670 1945.970 720.970 1964.030 ;
        RECT 724.350 1963.650 724.650 1990.550 ;
        RECT 728.030 1973.850 728.330 2000.750 ;
        RECT 731.710 1997.650 732.010 2051.750 ;
        RECT 727.110 1973.550 728.330 1973.850 ;
        RECT 730.790 1997.350 732.010 1997.650 ;
        RECT 724.350 1963.350 725.570 1963.650 ;
        RECT 717.910 1945.670 720.970 1945.970 ;
        RECT 717.910 1943.250 718.210 1945.670 ;
        RECT 716.990 1942.950 718.210 1943.250 ;
        RECT 716.055 1926.615 716.385 1926.945 ;
        RECT 716.070 1911.985 716.370 1926.615 ;
        RECT 716.990 1912.665 717.290 1942.950 ;
        RECT 718.815 1926.930 719.145 1926.945 ;
        RECT 725.270 1926.930 725.570 1963.350 ;
        RECT 718.815 1926.630 725.570 1926.930 ;
        RECT 718.815 1926.615 719.145 1926.630 ;
        RECT 727.110 1926.250 727.410 1973.550 ;
        RECT 718.830 1925.950 727.410 1926.250 ;
        RECT 718.830 1924.905 719.130 1925.950 ;
        RECT 718.815 1924.575 719.145 1924.905 ;
        RECT 718.815 1922.170 719.145 1922.185 ;
        RECT 730.790 1922.170 731.090 1997.350 ;
        RECT 718.815 1921.870 731.090 1922.170 ;
        RECT 718.815 1921.855 719.145 1921.870 ;
        RECT 716.975 1912.335 717.305 1912.665 ;
        RECT 718.815 1912.650 719.145 1912.665 ;
        RECT 718.815 1912.350 732.010 1912.650 ;
        RECT 718.815 1912.335 719.145 1912.350 ;
        RECT 716.055 1911.655 716.385 1911.985 ;
        RECT 718.815 1909.250 719.145 1909.265 ;
        RECT 718.815 1908.950 728.330 1909.250 ;
        RECT 718.815 1908.935 719.145 1908.950 ;
        RECT 716.975 1906.895 717.305 1907.225 ;
        RECT 716.990 1905.850 717.290 1906.895 ;
        RECT 718.815 1906.530 719.145 1906.545 ;
        RECT 718.815 1906.230 726.490 1906.530 ;
        RECT 718.815 1906.215 719.145 1906.230 ;
        RECT 716.990 1905.550 725.570 1905.850 ;
        RECT 725.270 1828.330 725.570 1905.550 ;
        RECT 726.190 1858.250 726.490 1906.230 ;
        RECT 726.190 1857.950 727.410 1858.250 ;
        RECT 727.110 1828.330 727.410 1857.950 ;
        RECT 723.430 1828.030 725.570 1828.330 ;
        RECT 726.190 1828.030 727.410 1828.330 ;
        RECT 718.815 1820.850 719.145 1820.865 ;
        RECT 718.815 1820.550 720.970 1820.850 ;
        RECT 718.815 1820.535 719.145 1820.550 ;
        RECT 720.670 1780.050 720.970 1820.550 ;
        RECT 718.830 1779.750 720.970 1780.050 ;
        RECT 718.830 1777.345 719.130 1779.750 ;
        RECT 718.815 1777.015 719.145 1777.345 ;
        RECT 723.430 1746.050 723.730 1828.030 ;
        RECT 726.190 1827.650 726.490 1828.030 ;
        RECT 725.270 1827.350 726.490 1827.650 ;
        RECT 725.270 1807.950 725.570 1827.350 ;
        RECT 728.030 1824.250 728.330 1908.950 ;
        RECT 731.710 1834.450 732.010 1912.350 ;
        RECT 729.870 1834.150 732.010 1834.450 ;
        RECT 729.870 1828.330 730.170 1834.150 ;
        RECT 727.110 1823.950 728.330 1824.250 ;
        RECT 728.950 1828.030 730.170 1828.330 ;
        RECT 725.270 1807.650 726.490 1807.950 ;
        RECT 726.190 1807.250 726.490 1807.650 ;
        RECT 727.110 1807.250 727.410 1823.950 ;
        RECT 728.950 1821.530 729.250 1828.030 ;
        RECT 728.950 1821.230 732.010 1821.530 ;
        RECT 731.710 1807.250 732.010 1821.230 ;
        RECT 724.350 1806.950 732.010 1807.250 ;
        RECT 724.350 1769.850 724.650 1806.950 ;
        RECT 726.190 1793.650 726.490 1806.950 ;
        RECT 727.110 1793.650 727.410 1806.950 ;
        RECT 726.190 1793.350 731.090 1793.650 ;
        RECT 727.110 1790.250 727.410 1793.350 ;
        RECT 727.110 1789.950 728.330 1790.250 ;
        RECT 724.350 1769.550 727.410 1769.850 ;
        RECT 727.110 1763.050 727.410 1769.550 ;
        RECT 728.030 1766.450 728.330 1789.950 ;
        RECT 730.790 1780.050 731.090 1793.350 ;
        RECT 730.790 1779.750 732.010 1780.050 ;
        RECT 728.030 1766.150 730.170 1766.450 ;
        RECT 727.110 1762.750 728.330 1763.050 ;
        RECT 723.430 1745.750 727.410 1746.050 ;
        RECT 714.215 1742.335 714.545 1742.665 ;
        RECT 718.815 1742.650 719.145 1742.665 ;
        RECT 727.110 1742.650 727.410 1745.750 ;
        RECT 718.815 1742.350 727.410 1742.650 ;
        RECT 718.815 1742.335 719.145 1742.350 ;
        RECT 714.230 1731.785 714.530 1742.335 ;
        RECT 718.815 1739.250 719.145 1739.265 ;
        RECT 728.030 1739.250 728.330 1762.750 ;
        RECT 718.815 1738.950 728.330 1739.250 ;
        RECT 718.815 1738.935 719.145 1738.950 ;
        RECT 729.870 1732.450 730.170 1766.150 ;
        RECT 718.830 1732.150 730.170 1732.450 ;
        RECT 712.375 1731.455 712.705 1731.785 ;
        RECT 714.215 1731.455 714.545 1731.785 ;
        RECT 712.390 1698.465 712.690 1731.455 ;
        RECT 718.830 1721.585 719.130 1732.150 ;
        RECT 718.815 1721.255 719.145 1721.585 ;
        RECT 718.815 1718.850 719.145 1718.865 ;
        RECT 718.815 1718.550 728.330 1718.850 ;
        RECT 718.815 1718.535 719.145 1718.550 ;
        RECT 712.375 1698.135 712.705 1698.465 ;
        RECT 718.815 1698.135 719.145 1698.465 ;
        RECT 718.830 1684.850 719.130 1698.135 ;
        RECT 728.030 1691.650 728.330 1718.550 ;
        RECT 728.030 1691.350 731.090 1691.650 ;
        RECT 718.830 1684.550 728.330 1684.850 ;
        RECT 718.815 1681.450 719.145 1681.465 ;
        RECT 718.815 1681.150 725.570 1681.450 ;
        RECT 718.815 1681.135 719.145 1681.150 ;
        RECT 718.815 1671.250 719.145 1671.265 ;
        RECT 725.270 1671.250 725.570 1681.150 ;
        RECT 718.815 1670.950 722.810 1671.250 ;
        RECT 725.270 1670.950 726.490 1671.250 ;
        RECT 718.815 1670.935 719.145 1670.950 ;
        RECT 714.215 1664.815 714.545 1665.145 ;
        RECT 718.815 1665.130 719.145 1665.145 ;
        RECT 722.510 1665.130 722.810 1670.950 ;
        RECT 718.815 1664.830 722.810 1665.130 ;
        RECT 718.815 1664.815 719.145 1664.830 ;
        RECT 714.230 1654.265 714.530 1664.815 ;
        RECT 718.815 1664.450 719.145 1664.465 ;
        RECT 726.190 1664.450 726.490 1670.950 ;
        RECT 728.030 1667.850 728.330 1684.550 ;
        RECT 718.815 1664.150 726.490 1664.450 ;
        RECT 727.110 1667.550 728.330 1667.850 ;
        RECT 718.815 1664.135 719.145 1664.150 ;
        RECT 718.815 1662.095 719.145 1662.425 ;
        RECT 718.830 1661.050 719.130 1662.095 ;
        RECT 727.110 1661.730 727.410 1667.550 ;
        RECT 730.790 1662.410 731.090 1691.350 ;
        RECT 722.510 1661.430 727.410 1661.730 ;
        RECT 729.870 1662.110 731.090 1662.410 ;
        RECT 722.510 1661.050 722.810 1661.430 ;
        RECT 718.830 1660.750 722.810 1661.050 ;
        RECT 729.870 1657.650 730.170 1662.110 ;
        RECT 731.710 1661.730 732.010 1779.750 ;
        RECT 717.910 1657.350 730.170 1657.650 ;
        RECT 730.790 1661.430 732.010 1661.730 ;
        RECT 714.215 1653.935 714.545 1654.265 ;
        RECT 717.910 1639.970 718.210 1657.350 ;
        RECT 718.815 1654.930 719.145 1654.945 ;
        RECT 730.790 1654.930 731.090 1661.430 ;
        RECT 718.815 1654.630 731.090 1654.930 ;
        RECT 718.815 1654.615 719.145 1654.630 ;
        RECT 718.815 1654.250 719.145 1654.265 ;
        RECT 718.815 1653.950 720.970 1654.250 ;
        RECT 718.815 1653.935 719.145 1653.950 ;
        RECT 720.670 1653.570 720.970 1653.950 ;
        RECT 720.670 1653.270 732.010 1653.570 ;
        RECT 717.910 1639.670 731.090 1639.970 ;
        RECT 718.815 1638.610 719.145 1638.625 ;
        RECT 718.815 1638.310 730.170 1638.610 ;
        RECT 718.815 1638.295 719.145 1638.310 ;
        RECT 718.815 1637.615 719.145 1637.945 ;
        RECT 718.830 1637.250 719.130 1637.615 ;
        RECT 718.830 1636.950 727.410 1637.250 ;
        RECT 718.815 1631.810 719.145 1631.825 ;
        RECT 718.815 1631.510 724.650 1631.810 ;
        RECT 718.815 1631.495 719.145 1631.510 ;
        RECT 724.350 1582.850 724.650 1631.510 ;
        RECT 727.110 1609.370 727.410 1636.950 ;
        RECT 727.110 1609.070 728.330 1609.370 ;
        RECT 728.030 1596.450 728.330 1609.070 ;
        RECT 728.030 1596.150 729.250 1596.450 ;
        RECT 724.350 1582.550 728.330 1582.850 ;
        RECT 728.030 1379.530 728.330 1582.550 ;
        RECT 727.110 1379.230 728.330 1379.530 ;
        RECT 727.110 1355.730 727.410 1379.230 ;
        RECT 727.110 1355.430 728.330 1355.730 ;
        RECT 725.060 1337.310 726.240 1338.490 ;
        RECT 725.270 1325.825 725.570 1337.310 ;
        RECT 725.255 1325.495 725.585 1325.825 ;
        RECT 728.030 1325.130 728.330 1355.430 ;
        RECT 728.950 1326.505 729.250 1596.150 ;
        RECT 728.935 1326.175 729.265 1326.505 ;
        RECT 729.870 1325.825 730.170 1638.310 ;
        RECT 730.790 1325.825 731.090 1639.670 ;
        RECT 731.710 1326.505 732.010 1653.270 ;
        RECT 931.830 1330.510 933.010 1331.690 ;
        RECT 734.950 1327.110 736.130 1328.290 ;
        RECT 731.695 1326.175 732.025 1326.505 ;
        RECT 729.855 1325.495 730.185 1325.825 ;
        RECT 730.775 1325.495 731.105 1325.825 ;
        RECT 728.030 1324.830 731.090 1325.130 ;
        RECT 730.790 1324.465 731.090 1324.830 ;
        RECT 735.390 1324.465 735.690 1327.110 ;
        RECT 730.775 1324.135 731.105 1324.465 ;
        RECT 735.375 1324.135 735.705 1324.465 ;
        RECT 932.270 1297.945 932.570 1330.510 ;
        RECT 1034.870 1327.110 1036.050 1328.290 ;
        RECT 932.255 1297.615 932.585 1297.945 ;
        RECT 953.415 1297.615 953.745 1297.945 ;
        RECT 953.430 1202.065 953.730 1297.615 ;
        RECT 953.415 1201.735 953.745 1202.065 ;
        RECT 952.495 1201.055 952.825 1201.385 ;
        RECT 952.510 1173.505 952.810 1201.055 ;
        RECT 952.495 1173.175 952.825 1173.505 ;
        RECT 953.415 1171.815 953.745 1172.145 ;
        RECT 953.430 1159.225 953.730 1171.815 ;
        RECT 953.415 1158.895 953.745 1159.225 ;
        RECT 954.335 1111.295 954.665 1111.625 ;
        RECT 954.350 1077.625 954.650 1111.295 ;
        RECT 954.335 1077.295 954.665 1077.625 ;
        RECT 953.415 1075.935 953.745 1076.265 ;
        RECT 953.430 1062.665 953.730 1075.935 ;
        RECT 953.415 1062.335 953.745 1062.665 ;
        RECT 954.335 1014.735 954.665 1015.065 ;
        RECT 954.350 981.065 954.650 1014.735 ;
        RECT 954.335 980.735 954.665 981.065 ;
        RECT 953.415 978.695 953.745 979.025 ;
        RECT 953.430 966.105 953.730 978.695 ;
        RECT 953.415 965.775 953.745 966.105 ;
        RECT 952.495 918.175 952.825 918.505 ;
        RECT 952.510 883.825 952.810 918.175 ;
        RECT 952.495 883.495 952.825 883.825 ;
        RECT 953.415 882.135 953.745 882.465 ;
        RECT 953.430 869.545 953.730 882.135 ;
        RECT 953.415 869.215 953.745 869.545 ;
        RECT 952.495 820.935 952.825 821.265 ;
        RECT 952.510 787.265 952.810 820.935 ;
        RECT 952.495 786.935 952.825 787.265 ;
        RECT 953.415 785.575 953.745 785.905 ;
        RECT 953.430 772.305 953.730 785.575 ;
        RECT 953.415 771.975 953.745 772.305 ;
        RECT 952.495 724.375 952.825 724.705 ;
        RECT 952.510 690.705 952.810 724.375 ;
        RECT 952.495 690.375 952.825 690.705 ;
        RECT 953.415 689.015 953.745 689.345 ;
        RECT 953.430 675.745 953.730 689.015 ;
        RECT 953.415 675.415 953.745 675.745 ;
        RECT 954.335 627.815 954.665 628.145 ;
        RECT 954.350 594.145 954.650 627.815 ;
        RECT 954.335 593.815 954.665 594.145 ;
        RECT 953.415 592.455 953.745 592.785 ;
        RECT 953.430 545.865 953.730 592.455 ;
        RECT 953.415 545.535 953.745 545.865 ;
        RECT 954.335 544.175 954.665 544.505 ;
        RECT 954.350 497.585 954.650 544.175 ;
        RECT 954.335 497.255 954.665 497.585 ;
        RECT 953.415 495.895 953.745 496.225 ;
        RECT 953.430 449.305 953.730 495.895 ;
        RECT 953.415 448.975 953.745 449.305 ;
        RECT 952.495 447.615 952.825 447.945 ;
        RECT 952.510 427.545 952.810 447.615 ;
        RECT 952.495 427.215 952.825 427.545 ;
        RECT 953.415 380.295 953.745 380.625 ;
        RECT 953.430 362.250 953.730 380.295 ;
        RECT 952.510 361.950 953.730 362.250 ;
        RECT 952.510 304.465 952.810 361.950 ;
        RECT 952.495 304.135 952.825 304.465 ;
        RECT 953.415 302.775 953.745 303.105 ;
        RECT 953.430 289.505 953.730 302.775 ;
        RECT 953.415 289.175 953.745 289.505 ;
        RECT 954.335 241.575 954.665 241.905 ;
        RECT 954.350 207.905 954.650 241.575 ;
        RECT 954.335 207.575 954.665 207.905 ;
        RECT 953.415 206.215 953.745 206.545 ;
        RECT 953.430 192.945 953.730 206.215 ;
        RECT 953.415 192.615 953.745 192.945 ;
        RECT 952.495 145.015 952.825 145.345 ;
        RECT 952.510 107.250 952.810 145.015 ;
        RECT 952.510 106.950 953.730 107.250 ;
        RECT 953.430 96.385 953.730 106.950 ;
        RECT 953.415 96.055 953.745 96.385 ;
        RECT 954.335 48.455 954.665 48.785 ;
        RECT 954.350 24.985 954.650 48.455 ;
        RECT 954.335 24.655 954.665 24.985 ;
        RECT 1035.310 14.785 1035.610 1327.110 ;
        RECT 1148.455 1326.175 1148.785 1326.505 ;
        RECT 1148.470 18.865 1148.770 1326.175 ;
        RECT 1148.455 18.535 1148.785 18.865 ;
        RECT 1035.295 14.455 1035.625 14.785 ;
      LAYER met5 ;
        RECT 722.780 2353.700 728.060 2355.300 ;
        RECT 726.460 2351.900 728.060 2353.700 ;
        RECT 726.460 2350.300 728.980 2351.900 ;
        RECT 724.850 1337.100 933.220 1338.700 ;
        RECT 931.620 1330.300 933.220 1337.100 ;
        RECT 734.740 1326.900 1036.260 1328.500 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 682.250 2353.040 682.570 2353.100 ;
        RECT 705.250 2353.040 705.570 2353.100 ;
        RECT 682.250 2352.900 705.570 2353.040 ;
        RECT 682.250 2352.840 682.570 2352.900 ;
        RECT 705.250 2352.840 705.570 2352.900 ;
        RECT 682.250 15.880 682.570 15.940 ;
        RECT 918.690 15.880 919.010 15.940 ;
        RECT 682.250 15.740 919.010 15.880 ;
        RECT 682.250 15.680 682.570 15.740 ;
        RECT 918.690 15.680 919.010 15.740 ;
      LAYER via ;
        RECT 682.280 2352.840 682.540 2353.100 ;
        RECT 705.280 2352.840 705.540 2353.100 ;
        RECT 682.280 15.680 682.540 15.940 ;
        RECT 918.720 15.680 918.980 15.940 ;
      LAYER met2 ;
        RECT 682.280 2352.810 682.540 2353.130 ;
        RECT 705.270 2352.955 705.550 2353.325 ;
        RECT 705.280 2352.810 705.540 2352.955 ;
        RECT 682.340 15.970 682.480 2352.810 ;
        RECT 682.280 15.650 682.540 15.970 ;
        RECT 918.720 15.650 918.980 15.970 ;
        RECT 918.780 2.400 918.920 15.650 ;
        RECT 918.570 -4.800 919.130 2.400 ;
      LAYER via2 ;
        RECT 705.270 2353.000 705.550 2353.280 ;
      LAYER met3 ;
        RECT 705.245 2353.290 705.575 2353.305 ;
        RECT 715.810 2353.290 719.810 2353.295 ;
        RECT 705.245 2352.990 719.810 2353.290 ;
        RECT 705.245 2352.975 705.575 2352.990 ;
        RECT 715.810 2352.695 719.810 2352.990 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 792.650 46.140 792.970 46.200 ;
        RECT 936.170 46.140 936.490 46.200 ;
        RECT 792.650 46.000 936.490 46.140 ;
        RECT 792.650 45.940 792.970 46.000 ;
        RECT 936.170 45.940 936.490 46.000 ;
      LAYER via ;
        RECT 792.680 45.940 792.940 46.200 ;
        RECT 936.200 45.940 936.460 46.200 ;
      LAYER met2 ;
        RECT 793.180 1323.690 793.460 1327.135 ;
        RECT 792.740 1323.550 793.460 1323.690 ;
        RECT 792.740 46.230 792.880 1323.550 ;
        RECT 793.180 1323.135 793.460 1323.550 ;
        RECT 792.680 45.910 792.940 46.230 ;
        RECT 936.200 45.910 936.460 46.230 ;
        RECT 936.260 2.400 936.400 45.910 ;
        RECT 936.050 -4.800 936.610 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1650.165 641.325 1650.335 717.655 ;
        RECT 1649.245 386.325 1649.415 434.775 ;
        RECT 1650.165 144.925 1650.335 193.035 ;
      LAYER mcon ;
        RECT 1650.165 717.485 1650.335 717.655 ;
        RECT 1649.245 434.605 1649.415 434.775 ;
        RECT 1650.165 192.865 1650.335 193.035 ;
      LAYER met1 ;
        RECT 1649.630 1304.480 1649.950 1304.540 ;
        RECT 1655.150 1304.480 1655.470 1304.540 ;
        RECT 1649.630 1304.340 1655.470 1304.480 ;
        RECT 1649.630 1304.280 1649.950 1304.340 ;
        RECT 1655.150 1304.280 1655.470 1304.340 ;
        RECT 1650.090 1207.240 1650.410 1207.300 ;
        RECT 1650.550 1207.240 1650.870 1207.300 ;
        RECT 1650.090 1207.100 1650.870 1207.240 ;
        RECT 1650.090 1207.040 1650.410 1207.100 ;
        RECT 1650.550 1207.040 1650.870 1207.100 ;
        RECT 1650.090 1110.680 1650.410 1110.740 ;
        RECT 1650.550 1110.680 1650.870 1110.740 ;
        RECT 1650.090 1110.540 1650.870 1110.680 ;
        RECT 1650.090 1110.480 1650.410 1110.540 ;
        RECT 1650.550 1110.480 1650.870 1110.540 ;
        RECT 1650.090 1014.120 1650.410 1014.180 ;
        RECT 1650.550 1014.120 1650.870 1014.180 ;
        RECT 1650.090 1013.980 1650.870 1014.120 ;
        RECT 1650.090 1013.920 1650.410 1013.980 ;
        RECT 1650.550 1013.920 1650.870 1013.980 ;
        RECT 1650.090 917.560 1650.410 917.620 ;
        RECT 1650.550 917.560 1650.870 917.620 ;
        RECT 1650.090 917.420 1650.870 917.560 ;
        RECT 1650.090 917.360 1650.410 917.420 ;
        RECT 1650.550 917.360 1650.870 917.420 ;
        RECT 1650.090 821.000 1650.410 821.060 ;
        RECT 1650.550 821.000 1650.870 821.060 ;
        RECT 1650.090 820.860 1650.870 821.000 ;
        RECT 1650.090 820.800 1650.410 820.860 ;
        RECT 1650.550 820.800 1650.870 820.860 ;
        RECT 1650.090 717.640 1650.410 717.700 ;
        RECT 1649.895 717.500 1650.410 717.640 ;
        RECT 1650.090 717.440 1650.410 717.500 ;
        RECT 1650.090 641.480 1650.410 641.540 ;
        RECT 1649.895 641.340 1650.410 641.480 ;
        RECT 1650.090 641.280 1650.410 641.340 ;
        RECT 1650.090 593.340 1650.410 593.600 ;
        RECT 1650.180 593.200 1650.320 593.340 ;
        RECT 1650.550 593.200 1650.870 593.260 ;
        RECT 1650.180 593.060 1650.870 593.200 ;
        RECT 1650.550 593.000 1650.870 593.060 ;
        RECT 1650.090 496.780 1650.410 497.040 ;
        RECT 1650.180 496.640 1650.320 496.780 ;
        RECT 1650.550 496.640 1650.870 496.700 ;
        RECT 1650.180 496.500 1650.870 496.640 ;
        RECT 1650.550 496.440 1650.870 496.500 ;
        RECT 1649.185 434.760 1649.475 434.805 ;
        RECT 1649.630 434.760 1649.950 434.820 ;
        RECT 1649.185 434.620 1649.950 434.760 ;
        RECT 1649.185 434.575 1649.475 434.620 ;
        RECT 1649.630 434.560 1649.950 434.620 ;
        RECT 1649.170 386.480 1649.490 386.540 ;
        RECT 1648.975 386.340 1649.490 386.480 ;
        RECT 1649.170 386.280 1649.490 386.340 ;
        RECT 1649.630 303.520 1649.950 303.580 ;
        RECT 1650.550 303.520 1650.870 303.580 ;
        RECT 1649.630 303.380 1650.870 303.520 ;
        RECT 1649.630 303.320 1649.950 303.380 ;
        RECT 1650.550 303.320 1650.870 303.380 ;
        RECT 1650.550 255.580 1650.870 255.640 ;
        RECT 1650.180 255.440 1650.870 255.580 ;
        RECT 1650.180 255.300 1650.320 255.440 ;
        RECT 1650.550 255.380 1650.870 255.440 ;
        RECT 1650.090 255.040 1650.410 255.300 ;
        RECT 1649.630 206.960 1649.950 207.020 ;
        RECT 1650.550 206.960 1650.870 207.020 ;
        RECT 1649.630 206.820 1650.870 206.960 ;
        RECT 1649.630 206.760 1649.950 206.820 ;
        RECT 1650.550 206.760 1650.870 206.820 ;
        RECT 1650.105 193.020 1650.395 193.065 ;
        RECT 1650.550 193.020 1650.870 193.080 ;
        RECT 1650.105 192.880 1650.870 193.020 ;
        RECT 1650.105 192.835 1650.395 192.880 ;
        RECT 1650.550 192.820 1650.870 192.880 ;
        RECT 1650.090 145.080 1650.410 145.140 ;
        RECT 1649.895 144.940 1650.410 145.080 ;
        RECT 1650.090 144.880 1650.410 144.940 ;
        RECT 972.050 26.420 972.370 26.480 ;
        RECT 1650.090 26.420 1650.410 26.480 ;
        RECT 972.050 26.280 1650.410 26.420 ;
        RECT 972.050 26.220 972.370 26.280 ;
        RECT 1650.090 26.220 1650.410 26.280 ;
      LAYER via ;
        RECT 1649.660 1304.280 1649.920 1304.540 ;
        RECT 1655.180 1304.280 1655.440 1304.540 ;
        RECT 1650.120 1207.040 1650.380 1207.300 ;
        RECT 1650.580 1207.040 1650.840 1207.300 ;
        RECT 1650.120 1110.480 1650.380 1110.740 ;
        RECT 1650.580 1110.480 1650.840 1110.740 ;
        RECT 1650.120 1013.920 1650.380 1014.180 ;
        RECT 1650.580 1013.920 1650.840 1014.180 ;
        RECT 1650.120 917.360 1650.380 917.620 ;
        RECT 1650.580 917.360 1650.840 917.620 ;
        RECT 1650.120 820.800 1650.380 821.060 ;
        RECT 1650.580 820.800 1650.840 821.060 ;
        RECT 1650.120 717.440 1650.380 717.700 ;
        RECT 1650.120 641.280 1650.380 641.540 ;
        RECT 1650.120 593.340 1650.380 593.600 ;
        RECT 1650.580 593.000 1650.840 593.260 ;
        RECT 1650.120 496.780 1650.380 497.040 ;
        RECT 1650.580 496.440 1650.840 496.700 ;
        RECT 1649.660 434.560 1649.920 434.820 ;
        RECT 1649.200 386.280 1649.460 386.540 ;
        RECT 1649.660 303.320 1649.920 303.580 ;
        RECT 1650.580 303.320 1650.840 303.580 ;
        RECT 1650.580 255.380 1650.840 255.640 ;
        RECT 1650.120 255.040 1650.380 255.300 ;
        RECT 1649.660 206.760 1649.920 207.020 ;
        RECT 1650.580 206.760 1650.840 207.020 ;
        RECT 1650.580 192.820 1650.840 193.080 ;
        RECT 1650.120 144.880 1650.380 145.140 ;
        RECT 972.080 26.220 972.340 26.480 ;
        RECT 1650.120 26.220 1650.380 26.480 ;
      LAYER met2 ;
        RECT 1655.220 1323.135 1655.500 1327.135 ;
        RECT 1655.240 1304.570 1655.380 1323.135 ;
        RECT 1649.660 1304.250 1649.920 1304.570 ;
        RECT 1655.180 1304.250 1655.440 1304.570 ;
        RECT 1649.720 1303.970 1649.860 1304.250 ;
        RECT 1649.720 1303.830 1650.780 1303.970 ;
        RECT 1650.640 1221.010 1650.780 1303.830 ;
        RECT 1650.180 1220.870 1650.780 1221.010 ;
        RECT 1650.180 1207.330 1650.320 1220.870 ;
        RECT 1650.120 1207.010 1650.380 1207.330 ;
        RECT 1650.580 1207.010 1650.840 1207.330 ;
        RECT 1650.640 1124.450 1650.780 1207.010 ;
        RECT 1650.180 1124.310 1650.780 1124.450 ;
        RECT 1650.180 1110.770 1650.320 1124.310 ;
        RECT 1650.120 1110.450 1650.380 1110.770 ;
        RECT 1650.580 1110.450 1650.840 1110.770 ;
        RECT 1650.640 1027.890 1650.780 1110.450 ;
        RECT 1650.180 1027.750 1650.780 1027.890 ;
        RECT 1650.180 1014.210 1650.320 1027.750 ;
        RECT 1650.120 1013.890 1650.380 1014.210 ;
        RECT 1650.580 1013.890 1650.840 1014.210 ;
        RECT 1650.640 931.330 1650.780 1013.890 ;
        RECT 1650.180 931.190 1650.780 931.330 ;
        RECT 1650.180 917.650 1650.320 931.190 ;
        RECT 1650.120 917.330 1650.380 917.650 ;
        RECT 1650.580 917.330 1650.840 917.650 ;
        RECT 1650.640 834.770 1650.780 917.330 ;
        RECT 1650.180 834.630 1650.780 834.770 ;
        RECT 1650.180 821.090 1650.320 834.630 ;
        RECT 1650.120 820.770 1650.380 821.090 ;
        RECT 1650.580 820.770 1650.840 821.090 ;
        RECT 1650.640 738.210 1650.780 820.770 ;
        RECT 1650.180 738.070 1650.780 738.210 ;
        RECT 1650.180 717.730 1650.320 738.070 ;
        RECT 1650.120 717.410 1650.380 717.730 ;
        RECT 1650.120 641.250 1650.380 641.570 ;
        RECT 1650.180 593.630 1650.320 641.250 ;
        RECT 1650.120 593.310 1650.380 593.630 ;
        RECT 1650.580 592.970 1650.840 593.290 ;
        RECT 1650.640 545.090 1650.780 592.970 ;
        RECT 1650.180 544.950 1650.780 545.090 ;
        RECT 1650.180 497.070 1650.320 544.950 ;
        RECT 1650.120 496.750 1650.380 497.070 ;
        RECT 1650.580 496.410 1650.840 496.730 ;
        RECT 1650.640 448.530 1650.780 496.410 ;
        RECT 1649.720 448.390 1650.780 448.530 ;
        RECT 1649.720 434.850 1649.860 448.390 ;
        RECT 1649.660 434.530 1649.920 434.850 ;
        RECT 1649.200 386.250 1649.460 386.570 ;
        RECT 1649.260 351.290 1649.400 386.250 ;
        RECT 1649.260 351.150 1649.860 351.290 ;
        RECT 1649.720 303.610 1649.860 351.150 ;
        RECT 1649.660 303.290 1649.920 303.610 ;
        RECT 1650.580 303.290 1650.840 303.610 ;
        RECT 1650.640 255.670 1650.780 303.290 ;
        RECT 1650.580 255.350 1650.840 255.670 ;
        RECT 1650.120 255.010 1650.380 255.330 ;
        RECT 1650.180 207.130 1650.320 255.010 ;
        RECT 1649.720 207.050 1650.320 207.130 ;
        RECT 1649.660 206.990 1650.320 207.050 ;
        RECT 1649.660 206.730 1649.920 206.990 ;
        RECT 1650.580 206.730 1650.840 207.050 ;
        RECT 1650.640 193.110 1650.780 206.730 ;
        RECT 1650.580 192.790 1650.840 193.110 ;
        RECT 1650.120 144.850 1650.380 145.170 ;
        RECT 1650.180 110.570 1650.320 144.850 ;
        RECT 1649.720 110.430 1650.320 110.570 ;
        RECT 1649.720 109.890 1649.860 110.430 ;
        RECT 1649.720 109.750 1650.320 109.890 ;
        RECT 1650.180 26.510 1650.320 109.750 ;
        RECT 972.080 26.190 972.340 26.510 ;
        RECT 1650.120 26.190 1650.380 26.510 ;
        RECT 972.140 2.400 972.280 26.190 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1559.930 2376.500 1560.250 2376.560 ;
        RECT 1564.070 2376.500 1564.390 2376.560 ;
        RECT 1559.930 2376.360 1564.390 2376.500 ;
        RECT 1559.930 2376.300 1560.250 2376.360 ;
        RECT 1564.070 2376.300 1564.390 2376.360 ;
        RECT 650.970 17.240 651.290 17.300 ;
        RECT 655.110 17.240 655.430 17.300 ;
        RECT 650.970 17.100 655.430 17.240 ;
        RECT 650.970 17.040 651.290 17.100 ;
        RECT 655.110 17.040 655.430 17.100 ;
      LAYER via ;
        RECT 1559.960 2376.300 1560.220 2376.560 ;
        RECT 1564.100 2376.300 1564.360 2376.560 ;
        RECT 651.000 17.040 651.260 17.300 ;
        RECT 655.140 17.040 655.400 17.300 ;
      LAYER met2 ;
        RECT 1558.640 2378.230 1560.160 2378.370 ;
        RECT 1558.640 2377.805 1558.780 2378.230 ;
        RECT 655.130 2377.435 655.410 2377.805 ;
        RECT 1558.570 2377.435 1558.850 2377.805 ;
        RECT 655.200 17.330 655.340 2377.435 ;
        RECT 1560.020 2376.590 1560.160 2378.230 ;
        RECT 1559.960 2376.270 1560.220 2376.590 ;
        RECT 1564.100 2376.330 1564.360 2376.590 ;
        RECT 1565.980 2376.330 1566.260 2377.880 ;
        RECT 1564.100 2376.270 1566.260 2376.330 ;
        RECT 1564.160 2376.190 1566.260 2376.270 ;
        RECT 1565.980 2373.880 1566.260 2376.190 ;
        RECT 651.000 17.010 651.260 17.330 ;
        RECT 655.140 17.010 655.400 17.330 ;
        RECT 651.060 2.400 651.200 17.010 ;
        RECT 650.850 -4.800 651.410 2.400 ;
      LAYER via2 ;
        RECT 655.130 2377.480 655.410 2377.760 ;
        RECT 1558.570 2377.480 1558.850 2377.760 ;
      LAYER met3 ;
        RECT 655.105 2377.770 655.435 2377.785 ;
        RECT 1558.545 2377.770 1558.875 2377.785 ;
        RECT 655.105 2377.470 1558.875 2377.770 ;
        RECT 655.105 2377.455 655.435 2377.470 ;
        RECT 1558.545 2377.455 1558.875 2377.470 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1756.425 1476.365 1756.595 1498.975 ;
      LAYER mcon ;
        RECT 1756.425 1498.805 1756.595 1498.975 ;
      LAYER met1 ;
        RECT 1754.970 1525.140 1755.290 1525.200 ;
        RECT 1758.190 1525.140 1758.510 1525.200 ;
        RECT 1754.970 1525.000 1758.510 1525.140 ;
        RECT 1754.970 1524.940 1755.290 1525.000 ;
        RECT 1758.190 1524.940 1758.510 1525.000 ;
        RECT 1754.970 1498.960 1755.290 1499.020 ;
        RECT 1756.365 1498.960 1756.655 1499.005 ;
        RECT 1754.970 1498.820 1756.655 1498.960 ;
        RECT 1754.970 1498.760 1755.290 1498.820 ;
        RECT 1756.365 1498.775 1756.655 1498.820 ;
        RECT 1754.970 1476.520 1755.290 1476.580 ;
        RECT 1756.365 1476.520 1756.655 1476.565 ;
        RECT 1754.970 1476.380 1756.655 1476.520 ;
        RECT 1754.970 1476.320 1755.290 1476.380 ;
        RECT 1756.365 1476.335 1756.655 1476.380 ;
        RECT 989.990 25.400 990.310 25.460 ;
        RECT 1754.970 25.400 1755.290 25.460 ;
        RECT 989.990 25.260 1755.290 25.400 ;
        RECT 989.990 25.200 990.310 25.260 ;
        RECT 1754.970 25.200 1755.290 25.260 ;
      LAYER via ;
        RECT 1755.000 1524.940 1755.260 1525.200 ;
        RECT 1758.220 1524.940 1758.480 1525.200 ;
        RECT 1755.000 1498.760 1755.260 1499.020 ;
        RECT 1755.000 1476.320 1755.260 1476.580 ;
        RECT 990.020 25.200 990.280 25.460 ;
        RECT 1755.000 25.200 1755.260 25.460 ;
      LAYER met2 ;
        RECT 1758.210 1525.395 1758.490 1525.765 ;
        RECT 1758.280 1525.230 1758.420 1525.395 ;
        RECT 1755.000 1524.910 1755.260 1525.230 ;
        RECT 1758.220 1524.910 1758.480 1525.230 ;
        RECT 1755.060 1499.050 1755.200 1524.910 ;
        RECT 1755.000 1498.730 1755.260 1499.050 ;
        RECT 1755.000 1476.290 1755.260 1476.610 ;
        RECT 1755.060 25.490 1755.200 1476.290 ;
        RECT 990.020 25.170 990.280 25.490 ;
        RECT 1755.000 25.170 1755.260 25.490 ;
        RECT 990.080 2.400 990.220 25.170 ;
        RECT 989.870 -4.800 990.430 2.400 ;
      LAYER via2 ;
        RECT 1758.210 1525.440 1758.490 1525.720 ;
      LAYER met3 ;
        RECT 1755.835 1527.175 1759.835 1527.775 ;
        RECT 1758.430 1525.745 1758.730 1527.175 ;
        RECT 1758.185 1525.430 1758.730 1525.745 ;
        RECT 1758.185 1525.415 1758.515 1525.430 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1007.470 27.440 1007.790 27.500 ;
        RECT 1386.970 27.440 1387.290 27.500 ;
        RECT 1007.470 27.300 1387.290 27.440 ;
        RECT 1007.470 27.240 1007.790 27.300 ;
        RECT 1386.970 27.240 1387.290 27.300 ;
      LAYER via ;
        RECT 1007.500 27.240 1007.760 27.500 ;
        RECT 1387.000 27.240 1387.260 27.500 ;
      LAYER met2 ;
        RECT 1389.340 1323.690 1389.620 1327.135 ;
        RECT 1387.060 1323.550 1389.620 1323.690 ;
        RECT 1387.060 27.530 1387.200 1323.550 ;
        RECT 1389.340 1323.135 1389.620 1323.550 ;
        RECT 1007.500 27.210 1007.760 27.530 ;
        RECT 1387.000 27.210 1387.260 27.530 ;
        RECT 1007.560 2.400 1007.700 27.210 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 806.450 24.720 806.770 24.780 ;
        RECT 1025.410 24.720 1025.730 24.780 ;
        RECT 806.450 24.580 1025.730 24.720 ;
        RECT 806.450 24.520 806.770 24.580 ;
        RECT 1025.410 24.520 1025.730 24.580 ;
      LAYER via ;
        RECT 806.480 24.520 806.740 24.780 ;
        RECT 1025.440 24.520 1025.700 24.780 ;
      LAYER met2 ;
        RECT 805.140 1323.690 805.420 1327.135 ;
        RECT 805.140 1323.550 806.680 1323.690 ;
        RECT 805.140 1323.135 805.420 1323.550 ;
        RECT 806.540 24.810 806.680 1323.550 ;
        RECT 806.480 24.490 806.740 24.810 ;
        RECT 1025.440 24.490 1025.700 24.810 ;
        RECT 1025.500 2.400 1025.640 24.490 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1757.805 1897.625 1757.975 1945.735 ;
      LAYER mcon ;
        RECT 1757.805 1945.565 1757.975 1945.735 ;
      LAYER met1 ;
        RECT 1757.730 1945.720 1758.050 1945.780 ;
        RECT 1757.535 1945.580 1758.050 1945.720 ;
        RECT 1757.730 1945.520 1758.050 1945.580 ;
        RECT 1757.745 1897.780 1758.035 1897.825 ;
        RECT 1758.190 1897.780 1758.510 1897.840 ;
        RECT 1757.745 1897.640 1758.510 1897.780 ;
        RECT 1757.745 1897.595 1758.035 1897.640 ;
        RECT 1758.190 1897.580 1758.510 1897.640 ;
        RECT 1043.350 20.640 1043.670 20.700 ;
        RECT 1047.490 20.640 1047.810 20.700 ;
        RECT 1043.350 20.500 1047.810 20.640 ;
        RECT 1043.350 20.440 1043.670 20.500 ;
        RECT 1047.490 20.440 1047.810 20.500 ;
      LAYER via ;
        RECT 1757.760 1945.520 1758.020 1945.780 ;
        RECT 1758.220 1897.580 1758.480 1897.840 ;
        RECT 1043.380 20.440 1043.640 20.700 ;
        RECT 1047.520 20.440 1047.780 20.700 ;
      LAYER met2 ;
        RECT 1757.750 1957.195 1758.030 1957.565 ;
        RECT 1757.820 1945.810 1757.960 1957.195 ;
        RECT 1757.760 1945.490 1758.020 1945.810 ;
        RECT 1758.220 1897.550 1758.480 1897.870 ;
        RECT 1758.280 1877.325 1758.420 1897.550 ;
        RECT 1758.210 1876.955 1758.490 1877.325 ;
        RECT 1047.510 86.515 1047.790 86.885 ;
        RECT 1047.580 20.730 1047.720 86.515 ;
        RECT 1043.380 20.410 1043.640 20.730 ;
        RECT 1047.520 20.410 1047.780 20.730 ;
        RECT 1043.440 2.400 1043.580 20.410 ;
        RECT 1043.230 -4.800 1043.790 2.400 ;
      LAYER via2 ;
        RECT 1757.750 1957.240 1758.030 1957.520 ;
        RECT 1758.210 1877.000 1758.490 1877.280 ;
        RECT 1047.510 86.560 1047.790 86.840 ;
      LAYER met3 ;
        RECT 1755.835 2305.095 1759.835 2305.695 ;
        RECT 1756.590 2302.980 1756.890 2305.095 ;
        RECT 1756.550 2302.660 1756.930 2302.980 ;
        RECT 1756.550 1957.530 1756.930 1957.540 ;
        RECT 1757.725 1957.530 1758.055 1957.545 ;
        RECT 1756.550 1957.230 1758.055 1957.530 ;
        RECT 1756.550 1957.220 1756.930 1957.230 ;
        RECT 1757.725 1957.215 1758.055 1957.230 ;
        RECT 1756.550 1877.290 1756.930 1877.300 ;
        RECT 1758.185 1877.290 1758.515 1877.305 ;
        RECT 1756.550 1876.990 1758.515 1877.290 ;
        RECT 1756.550 1876.980 1756.930 1876.990 ;
        RECT 1758.185 1876.975 1758.515 1876.990 ;
        RECT 1753.790 1326.490 1754.170 1326.500 ;
        RECT 1752.910 1326.190 1754.170 1326.490 ;
        RECT 1752.910 1325.140 1753.210 1326.190 ;
        RECT 1753.790 1326.180 1754.170 1326.190 ;
        RECT 1752.870 1324.820 1753.250 1325.140 ;
        RECT 1752.870 1294.530 1753.250 1294.540 ;
        RECT 1755.630 1294.530 1756.010 1294.540 ;
        RECT 1752.870 1294.230 1756.010 1294.530 ;
        RECT 1752.870 1294.220 1753.250 1294.230 ;
        RECT 1755.630 1294.220 1756.010 1294.230 ;
        RECT 1752.870 1245.570 1753.250 1245.580 ;
        RECT 1755.630 1245.570 1756.010 1245.580 ;
        RECT 1752.870 1245.270 1756.010 1245.570 ;
        RECT 1752.870 1245.260 1753.250 1245.270 ;
        RECT 1755.630 1245.260 1756.010 1245.270 ;
        RECT 1752.870 911.690 1753.250 911.700 ;
        RECT 1756.550 911.690 1756.930 911.700 ;
        RECT 1752.870 911.390 1756.930 911.690 ;
        RECT 1752.870 911.380 1753.250 911.390 ;
        RECT 1756.550 911.380 1756.930 911.390 ;
        RECT 1752.870 859.330 1753.250 859.340 ;
        RECT 1756.550 859.330 1756.930 859.340 ;
        RECT 1752.870 859.030 1756.930 859.330 ;
        RECT 1752.870 859.020 1753.250 859.030 ;
        RECT 1756.550 859.020 1756.930 859.030 ;
        RECT 1752.870 133.770 1753.250 133.780 ;
        RECT 1756.550 133.770 1756.930 133.780 ;
        RECT 1752.870 133.470 1756.930 133.770 ;
        RECT 1752.870 133.460 1753.250 133.470 ;
        RECT 1756.550 133.460 1756.930 133.470 ;
        RECT 1047.485 86.850 1047.815 86.865 ;
        RECT 1756.550 86.850 1756.930 86.860 ;
        RECT 1047.485 86.550 1756.930 86.850 ;
        RECT 1047.485 86.535 1047.815 86.550 ;
        RECT 1756.550 86.540 1756.930 86.550 ;
      LAYER via3 ;
        RECT 1756.580 2302.660 1756.900 2302.980 ;
        RECT 1756.580 1957.220 1756.900 1957.540 ;
        RECT 1756.580 1876.980 1756.900 1877.300 ;
        RECT 1753.820 1326.180 1754.140 1326.500 ;
        RECT 1752.900 1324.820 1753.220 1325.140 ;
        RECT 1752.900 1294.220 1753.220 1294.540 ;
        RECT 1755.660 1294.220 1755.980 1294.540 ;
        RECT 1752.900 1245.260 1753.220 1245.580 ;
        RECT 1755.660 1245.260 1755.980 1245.580 ;
        RECT 1752.900 911.380 1753.220 911.700 ;
        RECT 1756.580 911.380 1756.900 911.700 ;
        RECT 1752.900 859.020 1753.220 859.340 ;
        RECT 1756.580 859.020 1756.900 859.340 ;
        RECT 1752.900 133.460 1753.220 133.780 ;
        RECT 1756.580 133.460 1756.900 133.780 ;
        RECT 1756.580 86.540 1756.900 86.860 ;
      LAYER met4 ;
        RECT 1756.575 2302.970 1756.905 2302.985 ;
        RECT 1753.830 2302.670 1756.905 2302.970 ;
        RECT 1753.830 2262.850 1754.130 2302.670 ;
        RECT 1756.575 2302.655 1756.905 2302.670 ;
        RECT 1752.910 2262.550 1754.130 2262.850 ;
        RECT 1752.910 2256.050 1753.210 2262.550 ;
        RECT 1751.070 2255.750 1753.210 2256.050 ;
        RECT 1751.070 2208.450 1751.370 2255.750 ;
        RECT 1751.070 2208.150 1754.130 2208.450 ;
        RECT 1753.830 2174.450 1754.130 2208.150 ;
        RECT 1752.910 2174.150 1754.130 2174.450 ;
        RECT 1752.910 2167.650 1753.210 2174.150 ;
        RECT 1752.910 2167.350 1754.130 2167.650 ;
        RECT 1753.830 2076.530 1754.130 2167.350 ;
        RECT 1751.990 2076.230 1754.130 2076.530 ;
        RECT 1751.990 2018.050 1752.290 2076.230 ;
        RECT 1751.990 2017.750 1754.130 2018.050 ;
        RECT 1753.830 2014.650 1754.130 2017.750 ;
        RECT 1753.830 2014.350 1757.810 2014.650 ;
        RECT 1757.510 2007.850 1757.810 2014.350 ;
        RECT 1756.590 2007.550 1757.810 2007.850 ;
        RECT 1756.590 1997.650 1756.890 2007.550 ;
        RECT 1754.750 1997.350 1756.890 1997.650 ;
        RECT 1754.750 1960.250 1755.050 1997.350 ;
        RECT 1754.750 1959.950 1756.890 1960.250 ;
        RECT 1756.590 1957.545 1756.890 1959.950 ;
        RECT 1756.575 1957.215 1756.905 1957.545 ;
        RECT 1756.575 1877.290 1756.905 1877.305 ;
        RECT 1754.750 1876.990 1756.905 1877.290 ;
        RECT 1754.750 1859.610 1755.050 1876.990 ;
        RECT 1756.575 1876.975 1756.905 1876.990 ;
        RECT 1751.990 1859.310 1755.050 1859.610 ;
        RECT 1751.990 1803.850 1752.290 1859.310 ;
        RECT 1750.150 1803.550 1752.290 1803.850 ;
        RECT 1750.150 1769.850 1750.450 1803.550 ;
        RECT 1750.150 1769.550 1751.370 1769.850 ;
        RECT 1751.070 1678.050 1751.370 1769.550 ;
        RECT 1751.070 1677.750 1753.210 1678.050 ;
        RECT 1752.910 1582.850 1753.210 1677.750 ;
        RECT 1751.990 1582.550 1753.210 1582.850 ;
        RECT 1751.990 1528.450 1752.290 1582.550 ;
        RECT 1751.990 1528.150 1753.210 1528.450 ;
        RECT 1752.910 1404.010 1753.210 1528.150 ;
        RECT 1752.910 1403.710 1754.130 1404.010 ;
        RECT 1753.830 1396.530 1754.130 1403.710 ;
        RECT 1752.910 1396.230 1754.130 1396.530 ;
        RECT 1752.910 1367.290 1753.210 1396.230 ;
        RECT 1752.910 1366.990 1754.130 1367.290 ;
        RECT 1753.830 1326.505 1754.130 1366.990 ;
        RECT 1753.815 1326.175 1754.145 1326.505 ;
        RECT 1752.895 1324.815 1753.225 1325.145 ;
        RECT 1752.910 1294.545 1753.210 1324.815 ;
        RECT 1752.895 1294.215 1753.225 1294.545 ;
        RECT 1755.655 1294.215 1755.985 1294.545 ;
        RECT 1755.670 1245.585 1755.970 1294.215 ;
        RECT 1752.895 1245.255 1753.225 1245.585 ;
        RECT 1755.655 1245.255 1755.985 1245.585 ;
        RECT 1752.910 911.705 1753.210 1245.255 ;
        RECT 1752.895 911.375 1753.225 911.705 ;
        RECT 1756.575 911.375 1756.905 911.705 ;
        RECT 1756.590 859.345 1756.890 911.375 ;
        RECT 1752.895 859.015 1753.225 859.345 ;
        RECT 1756.575 859.015 1756.905 859.345 ;
        RECT 1752.910 133.785 1753.210 859.015 ;
        RECT 1752.895 133.455 1753.225 133.785 ;
        RECT 1756.575 133.455 1756.905 133.785 ;
        RECT 1756.590 86.865 1756.890 133.455 ;
        RECT 1756.575 86.535 1756.905 86.865 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1754.585 1745.305 1754.755 1808.375 ;
        RECT 1754.585 1704.165 1754.755 1738.675 ;
        RECT 1755.045 1635.485 1755.215 1649.255 ;
      LAYER mcon ;
        RECT 1754.585 1808.205 1754.755 1808.375 ;
        RECT 1754.585 1738.505 1754.755 1738.675 ;
        RECT 1755.045 1649.085 1755.215 1649.255 ;
      LAYER met1 ;
        RECT 1754.510 1850.860 1754.830 1850.920 ;
        RECT 1757.270 1850.860 1757.590 1850.920 ;
        RECT 1754.510 1850.720 1757.590 1850.860 ;
        RECT 1754.510 1850.660 1754.830 1850.720 ;
        RECT 1757.270 1850.660 1757.590 1850.720 ;
        RECT 1754.510 1808.360 1754.830 1808.420 ;
        RECT 1754.315 1808.220 1754.830 1808.360 ;
        RECT 1754.510 1808.160 1754.830 1808.220 ;
        RECT 1754.510 1745.460 1754.830 1745.520 ;
        RECT 1754.315 1745.320 1754.830 1745.460 ;
        RECT 1754.510 1745.260 1754.830 1745.320 ;
        RECT 1754.510 1738.660 1754.830 1738.720 ;
        RECT 1754.315 1738.520 1754.830 1738.660 ;
        RECT 1754.510 1738.460 1754.830 1738.520 ;
        RECT 1754.510 1704.320 1754.830 1704.380 ;
        RECT 1754.315 1704.180 1754.830 1704.320 ;
        RECT 1754.510 1704.120 1754.830 1704.180 ;
        RECT 1754.510 1649.240 1754.830 1649.300 ;
        RECT 1754.985 1649.240 1755.275 1649.285 ;
        RECT 1754.510 1649.100 1755.275 1649.240 ;
        RECT 1754.510 1649.040 1754.830 1649.100 ;
        RECT 1754.985 1649.055 1755.275 1649.100 ;
        RECT 1754.970 1635.640 1755.290 1635.700 ;
        RECT 1754.775 1635.500 1755.290 1635.640 ;
        RECT 1754.970 1635.440 1755.290 1635.500 ;
        RECT 1752.670 1332.700 1752.990 1332.760 ;
        RECT 1753.590 1332.700 1753.910 1332.760 ;
        RECT 1752.670 1332.560 1753.910 1332.700 ;
        RECT 1752.670 1332.500 1752.990 1332.560 ;
        RECT 1753.590 1332.500 1753.910 1332.560 ;
        RECT 1752.670 907.360 1752.990 907.420 ;
        RECT 1753.590 907.360 1753.910 907.420 ;
        RECT 1752.670 907.220 1753.910 907.360 ;
        RECT 1752.670 907.160 1752.990 907.220 ;
        RECT 1753.590 907.160 1753.910 907.220 ;
        RECT 1753.590 158.820 1753.910 159.080 ;
        RECT 1753.680 158.400 1753.820 158.820 ;
        RECT 1753.590 158.140 1753.910 158.400 ;
        RECT 1753.590 135.360 1753.910 135.620 ;
        RECT 1753.680 134.540 1753.820 135.360 ;
        RECT 1754.050 134.540 1754.370 134.600 ;
        RECT 1753.680 134.400 1754.370 134.540 ;
        RECT 1754.050 134.340 1754.370 134.400 ;
        RECT 1062.210 86.940 1062.530 87.000 ;
        RECT 1754.050 86.940 1754.370 87.000 ;
        RECT 1062.210 86.800 1754.370 86.940 ;
        RECT 1062.210 86.740 1062.530 86.800 ;
        RECT 1754.050 86.740 1754.370 86.800 ;
        RECT 1061.290 2.960 1061.610 3.020 ;
        RECT 1062.210 2.960 1062.530 3.020 ;
        RECT 1061.290 2.820 1062.530 2.960 ;
        RECT 1061.290 2.760 1061.610 2.820 ;
        RECT 1062.210 2.760 1062.530 2.820 ;
      LAYER via ;
        RECT 1754.540 1850.660 1754.800 1850.920 ;
        RECT 1757.300 1850.660 1757.560 1850.920 ;
        RECT 1754.540 1808.160 1754.800 1808.420 ;
        RECT 1754.540 1745.260 1754.800 1745.520 ;
        RECT 1754.540 1738.460 1754.800 1738.720 ;
        RECT 1754.540 1704.120 1754.800 1704.380 ;
        RECT 1754.540 1649.040 1754.800 1649.300 ;
        RECT 1755.000 1635.440 1755.260 1635.700 ;
        RECT 1752.700 1332.500 1752.960 1332.760 ;
        RECT 1753.620 1332.500 1753.880 1332.760 ;
        RECT 1752.700 907.160 1752.960 907.420 ;
        RECT 1753.620 907.160 1753.880 907.420 ;
        RECT 1753.620 158.820 1753.880 159.080 ;
        RECT 1753.620 158.140 1753.880 158.400 ;
        RECT 1753.620 135.360 1753.880 135.620 ;
        RECT 1754.080 134.340 1754.340 134.600 ;
        RECT 1062.240 86.740 1062.500 87.000 ;
        RECT 1754.080 86.740 1754.340 87.000 ;
        RECT 1061.320 2.760 1061.580 3.020 ;
        RECT 1062.240 2.760 1062.500 3.020 ;
      LAYER met2 ;
        RECT 1757.290 1851.115 1757.570 1851.485 ;
        RECT 1757.360 1850.950 1757.500 1851.115 ;
        RECT 1754.540 1850.630 1754.800 1850.950 ;
        RECT 1757.300 1850.630 1757.560 1850.950 ;
        RECT 1754.600 1808.450 1754.740 1850.630 ;
        RECT 1754.540 1808.130 1754.800 1808.450 ;
        RECT 1754.540 1745.230 1754.800 1745.550 ;
        RECT 1754.600 1738.750 1754.740 1745.230 ;
        RECT 1754.540 1738.430 1754.800 1738.750 ;
        RECT 1754.540 1704.090 1754.800 1704.410 ;
        RECT 1754.600 1690.890 1754.740 1704.090 ;
        RECT 1753.680 1690.750 1754.740 1690.890 ;
        RECT 1753.680 1690.210 1753.820 1690.750 ;
        RECT 1753.680 1690.070 1754.280 1690.210 ;
        RECT 1754.140 1649.240 1754.280 1690.070 ;
        RECT 1754.540 1649.240 1754.800 1649.330 ;
        RECT 1754.140 1649.100 1754.800 1649.240 ;
        RECT 1754.540 1649.010 1754.800 1649.100 ;
        RECT 1755.000 1635.410 1755.260 1635.730 ;
        RECT 1755.060 1606.570 1755.200 1635.410 ;
        RECT 1752.760 1606.430 1755.200 1606.570 ;
        RECT 1752.760 1498.450 1752.900 1606.430 ;
        RECT 1752.760 1498.310 1753.360 1498.450 ;
        RECT 1753.220 1497.770 1753.360 1498.310 ;
        RECT 1753.220 1497.630 1755.200 1497.770 ;
        RECT 1755.060 1483.490 1755.200 1497.630 ;
        RECT 1753.680 1483.350 1755.200 1483.490 ;
        RECT 1753.680 1332.790 1753.820 1483.350 ;
        RECT 1752.700 1332.470 1752.960 1332.790 ;
        RECT 1753.620 1332.470 1753.880 1332.790 ;
        RECT 1752.760 1246.170 1752.900 1332.470 ;
        RECT 1752.760 1246.030 1753.360 1246.170 ;
        RECT 1753.220 1244.810 1753.360 1246.030 ;
        RECT 1753.220 1244.670 1753.820 1244.810 ;
        RECT 1753.680 907.450 1753.820 1244.670 ;
        RECT 1752.700 907.130 1752.960 907.450 ;
        RECT 1753.620 907.130 1753.880 907.450 ;
        RECT 1752.760 859.930 1752.900 907.130 ;
        RECT 1752.760 859.790 1753.360 859.930 ;
        RECT 1753.220 858.570 1753.360 859.790 ;
        RECT 1753.220 858.430 1753.820 858.570 ;
        RECT 1753.680 159.110 1753.820 858.430 ;
        RECT 1753.620 158.790 1753.880 159.110 ;
        RECT 1753.620 158.110 1753.880 158.430 ;
        RECT 1753.680 135.650 1753.820 158.110 ;
        RECT 1753.620 135.330 1753.880 135.650 ;
        RECT 1754.080 134.310 1754.340 134.630 ;
        RECT 1754.140 87.030 1754.280 134.310 ;
        RECT 1062.240 86.710 1062.500 87.030 ;
        RECT 1754.080 86.710 1754.340 87.030 ;
        RECT 1062.300 3.050 1062.440 86.710 ;
        RECT 1061.320 2.730 1061.580 3.050 ;
        RECT 1062.240 2.730 1062.500 3.050 ;
        RECT 1061.380 2.400 1061.520 2.730 ;
        RECT 1061.170 -4.800 1061.730 2.400 ;
      LAYER via2 ;
        RECT 1757.290 1851.160 1757.570 1851.440 ;
      LAYER met3 ;
        RECT 1755.835 1852.215 1759.835 1852.815 ;
        RECT 1757.510 1851.465 1757.810 1852.215 ;
        RECT 1757.265 1851.150 1757.810 1851.465 ;
        RECT 1757.265 1851.135 1757.595 1851.150 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1082.985 1297.185 1083.155 1322.515 ;
        RECT 1082.065 1110.865 1082.235 1124.975 ;
        RECT 1082.065 1014.305 1082.235 1028.415 ;
        RECT 1082.525 786.505 1082.695 821.015 ;
        RECT 1082.525 689.605 1082.695 724.455 ;
        RECT 1082.525 579.785 1082.695 593.895 ;
        RECT 1082.525 496.485 1082.695 531.335 ;
        RECT 1082.525 386.325 1082.695 434.775 ;
        RECT 1082.525 241.485 1082.695 289.595 ;
      LAYER mcon ;
        RECT 1082.985 1322.345 1083.155 1322.515 ;
        RECT 1082.065 1124.805 1082.235 1124.975 ;
        RECT 1082.065 1028.245 1082.235 1028.415 ;
        RECT 1082.525 820.845 1082.695 821.015 ;
        RECT 1082.525 724.285 1082.695 724.455 ;
        RECT 1082.525 593.725 1082.695 593.895 ;
        RECT 1082.525 531.165 1082.695 531.335 ;
        RECT 1082.525 434.605 1082.695 434.775 ;
        RECT 1082.525 289.425 1082.695 289.595 ;
      LAYER met1 ;
        RECT 1771.990 2021.880 1772.310 2021.940 ;
        RECT 1786.710 2021.880 1787.030 2021.940 ;
        RECT 1771.990 2021.740 1787.030 2021.880 ;
        RECT 1771.990 2021.680 1772.310 2021.740 ;
        RECT 1786.710 2021.680 1787.030 2021.740 ;
        RECT 1082.925 1322.500 1083.215 1322.545 ;
        RECT 1786.710 1322.500 1787.030 1322.560 ;
        RECT 1082.925 1322.360 1787.030 1322.500 ;
        RECT 1082.925 1322.315 1083.215 1322.360 ;
        RECT 1786.710 1322.300 1787.030 1322.360 ;
        RECT 1082.910 1297.340 1083.230 1297.400 ;
        RECT 1082.715 1297.200 1083.230 1297.340 ;
        RECT 1082.910 1297.140 1083.230 1297.200 ;
        RECT 1082.910 1173.580 1083.230 1173.640 ;
        RECT 1082.540 1173.440 1083.230 1173.580 ;
        RECT 1082.540 1172.960 1082.680 1173.440 ;
        RECT 1082.910 1173.380 1083.230 1173.440 ;
        RECT 1082.450 1172.700 1082.770 1172.960 ;
        RECT 1081.990 1124.960 1082.310 1125.020 ;
        RECT 1081.795 1124.820 1082.310 1124.960 ;
        RECT 1081.990 1124.760 1082.310 1124.820 ;
        RECT 1081.990 1111.020 1082.310 1111.080 ;
        RECT 1081.795 1110.880 1082.310 1111.020 ;
        RECT 1081.990 1110.820 1082.310 1110.880 ;
        RECT 1081.990 1076.480 1082.310 1076.740 ;
        RECT 1082.080 1076.000 1082.220 1076.480 ;
        RECT 1082.450 1076.000 1082.770 1076.060 ;
        RECT 1082.080 1075.860 1082.770 1076.000 ;
        RECT 1082.450 1075.800 1082.770 1075.860 ;
        RECT 1081.990 1028.400 1082.310 1028.460 ;
        RECT 1081.795 1028.260 1082.310 1028.400 ;
        RECT 1081.990 1028.200 1082.310 1028.260 ;
        RECT 1081.990 1014.460 1082.310 1014.520 ;
        RECT 1081.795 1014.320 1082.310 1014.460 ;
        RECT 1081.990 1014.260 1082.310 1014.320 ;
        RECT 1081.990 980.260 1082.310 980.520 ;
        RECT 1082.080 979.840 1082.220 980.260 ;
        RECT 1081.990 979.580 1082.310 979.840 ;
        RECT 1081.530 869.620 1081.850 869.680 ;
        RECT 1082.910 869.620 1083.230 869.680 ;
        RECT 1081.530 869.480 1083.230 869.620 ;
        RECT 1081.530 869.420 1081.850 869.480 ;
        RECT 1082.910 869.420 1083.230 869.480 ;
        RECT 1081.990 835.280 1082.310 835.340 ;
        RECT 1082.910 835.280 1083.230 835.340 ;
        RECT 1081.990 835.140 1083.230 835.280 ;
        RECT 1081.990 835.080 1082.310 835.140 ;
        RECT 1082.910 835.080 1083.230 835.140 ;
        RECT 1082.450 821.000 1082.770 821.060 ;
        RECT 1082.255 820.860 1082.770 821.000 ;
        RECT 1082.450 820.800 1082.770 820.860 ;
        RECT 1082.450 786.660 1082.770 786.720 ;
        RECT 1082.255 786.520 1082.770 786.660 ;
        RECT 1082.450 786.460 1082.770 786.520 ;
        RECT 1081.990 738.380 1082.310 738.440 ;
        RECT 1082.910 738.380 1083.230 738.440 ;
        RECT 1081.990 738.240 1083.230 738.380 ;
        RECT 1081.990 738.180 1082.310 738.240 ;
        RECT 1082.910 738.180 1083.230 738.240 ;
        RECT 1082.450 724.440 1082.770 724.500 ;
        RECT 1082.255 724.300 1082.770 724.440 ;
        RECT 1082.450 724.240 1082.770 724.300 ;
        RECT 1082.450 689.760 1082.770 689.820 ;
        RECT 1082.255 689.620 1082.770 689.760 ;
        RECT 1082.450 689.560 1082.770 689.620 ;
        RECT 1081.990 641.820 1082.310 641.880 ;
        RECT 1082.910 641.820 1083.230 641.880 ;
        RECT 1081.990 641.680 1083.230 641.820 ;
        RECT 1081.990 641.620 1082.310 641.680 ;
        RECT 1082.910 641.620 1083.230 641.680 ;
        RECT 1082.465 593.880 1082.755 593.925 ;
        RECT 1082.910 593.880 1083.230 593.940 ;
        RECT 1082.465 593.740 1083.230 593.880 ;
        RECT 1082.465 593.695 1082.755 593.740 ;
        RECT 1082.910 593.680 1083.230 593.740 ;
        RECT 1082.450 579.940 1082.770 580.000 ;
        RECT 1082.255 579.800 1082.770 579.940 ;
        RECT 1082.450 579.740 1082.770 579.800 ;
        RECT 1082.450 531.320 1082.770 531.380 ;
        RECT 1082.255 531.180 1082.770 531.320 ;
        RECT 1082.450 531.120 1082.770 531.180 ;
        RECT 1082.450 496.640 1082.770 496.700 ;
        RECT 1082.255 496.500 1082.770 496.640 ;
        RECT 1082.450 496.440 1082.770 496.500 ;
        RECT 1081.990 448.700 1082.310 448.760 ;
        RECT 1082.910 448.700 1083.230 448.760 ;
        RECT 1081.990 448.560 1083.230 448.700 ;
        RECT 1081.990 448.500 1082.310 448.560 ;
        RECT 1082.910 448.500 1083.230 448.560 ;
        RECT 1082.450 434.760 1082.770 434.820 ;
        RECT 1082.255 434.620 1082.770 434.760 ;
        RECT 1082.450 434.560 1082.770 434.620 ;
        RECT 1082.465 386.480 1082.755 386.525 ;
        RECT 1082.910 386.480 1083.230 386.540 ;
        RECT 1082.465 386.340 1083.230 386.480 ;
        RECT 1082.465 386.295 1082.755 386.340 ;
        RECT 1082.910 386.280 1083.230 386.340 ;
        RECT 1082.465 289.580 1082.755 289.625 ;
        RECT 1082.910 289.580 1083.230 289.640 ;
        RECT 1082.465 289.440 1083.230 289.580 ;
        RECT 1082.465 289.395 1082.755 289.440 ;
        RECT 1082.910 289.380 1083.230 289.440 ;
        RECT 1082.450 241.640 1082.770 241.700 ;
        RECT 1082.255 241.500 1082.770 241.640 ;
        RECT 1082.450 241.440 1082.770 241.500 ;
        RECT 1079.230 15.200 1079.550 15.260 ;
        RECT 1081.990 15.200 1082.310 15.260 ;
        RECT 1079.230 15.060 1082.310 15.200 ;
        RECT 1079.230 15.000 1079.550 15.060 ;
        RECT 1081.990 15.000 1082.310 15.060 ;
      LAYER via ;
        RECT 1772.020 2021.680 1772.280 2021.940 ;
        RECT 1786.740 2021.680 1787.000 2021.940 ;
        RECT 1786.740 1322.300 1787.000 1322.560 ;
        RECT 1082.940 1297.140 1083.200 1297.400 ;
        RECT 1082.940 1173.380 1083.200 1173.640 ;
        RECT 1082.480 1172.700 1082.740 1172.960 ;
        RECT 1082.020 1124.760 1082.280 1125.020 ;
        RECT 1082.020 1110.820 1082.280 1111.080 ;
        RECT 1082.020 1076.480 1082.280 1076.740 ;
        RECT 1082.480 1075.800 1082.740 1076.060 ;
        RECT 1082.020 1028.200 1082.280 1028.460 ;
        RECT 1082.020 1014.260 1082.280 1014.520 ;
        RECT 1082.020 980.260 1082.280 980.520 ;
        RECT 1082.020 979.580 1082.280 979.840 ;
        RECT 1081.560 869.420 1081.820 869.680 ;
        RECT 1082.940 869.420 1083.200 869.680 ;
        RECT 1082.020 835.080 1082.280 835.340 ;
        RECT 1082.940 835.080 1083.200 835.340 ;
        RECT 1082.480 820.800 1082.740 821.060 ;
        RECT 1082.480 786.460 1082.740 786.720 ;
        RECT 1082.020 738.180 1082.280 738.440 ;
        RECT 1082.940 738.180 1083.200 738.440 ;
        RECT 1082.480 724.240 1082.740 724.500 ;
        RECT 1082.480 689.560 1082.740 689.820 ;
        RECT 1082.020 641.620 1082.280 641.880 ;
        RECT 1082.940 641.620 1083.200 641.880 ;
        RECT 1082.940 593.680 1083.200 593.940 ;
        RECT 1082.480 579.740 1082.740 580.000 ;
        RECT 1082.480 531.120 1082.740 531.380 ;
        RECT 1082.480 496.440 1082.740 496.700 ;
        RECT 1082.020 448.500 1082.280 448.760 ;
        RECT 1082.940 448.500 1083.200 448.760 ;
        RECT 1082.480 434.560 1082.740 434.820 ;
        RECT 1082.940 386.280 1083.200 386.540 ;
        RECT 1082.940 289.380 1083.200 289.640 ;
        RECT 1082.480 241.440 1082.740 241.700 ;
        RECT 1079.260 15.000 1079.520 15.260 ;
        RECT 1082.020 15.000 1082.280 15.260 ;
      LAYER met2 ;
        RECT 1772.010 2023.835 1772.290 2024.205 ;
        RECT 1772.080 2021.970 1772.220 2023.835 ;
        RECT 1772.020 2021.650 1772.280 2021.970 ;
        RECT 1786.740 2021.650 1787.000 2021.970 ;
        RECT 1786.800 1322.590 1786.940 2021.650 ;
        RECT 1786.740 1322.270 1787.000 1322.590 ;
        RECT 1082.940 1297.110 1083.200 1297.430 ;
        RECT 1083.000 1173.670 1083.140 1297.110 ;
        RECT 1082.940 1173.350 1083.200 1173.670 ;
        RECT 1082.480 1172.670 1082.740 1172.990 ;
        RECT 1082.540 1159.130 1082.680 1172.670 ;
        RECT 1082.080 1158.990 1082.680 1159.130 ;
        RECT 1082.080 1125.050 1082.220 1158.990 ;
        RECT 1082.020 1124.730 1082.280 1125.050 ;
        RECT 1082.020 1110.790 1082.280 1111.110 ;
        RECT 1082.080 1076.770 1082.220 1110.790 ;
        RECT 1082.020 1076.450 1082.280 1076.770 ;
        RECT 1082.480 1075.770 1082.740 1076.090 ;
        RECT 1082.540 1062.570 1082.680 1075.770 ;
        RECT 1082.080 1062.430 1082.680 1062.570 ;
        RECT 1082.080 1028.490 1082.220 1062.430 ;
        RECT 1082.020 1028.170 1082.280 1028.490 ;
        RECT 1082.020 1014.230 1082.280 1014.550 ;
        RECT 1082.080 980.550 1082.220 1014.230 ;
        RECT 1082.020 980.230 1082.280 980.550 ;
        RECT 1082.020 979.550 1082.280 979.870 ;
        RECT 1082.080 978.930 1082.220 979.550 ;
        RECT 1082.080 978.790 1082.680 978.930 ;
        RECT 1082.540 932.010 1082.680 978.790 ;
        RECT 1082.080 931.870 1082.680 932.010 ;
        RECT 1082.080 931.330 1082.220 931.870 ;
        RECT 1082.080 931.190 1082.680 931.330 ;
        RECT 1082.540 917.845 1082.680 931.190 ;
        RECT 1081.550 917.475 1081.830 917.845 ;
        RECT 1082.470 917.475 1082.750 917.845 ;
        RECT 1081.620 869.710 1081.760 917.475 ;
        RECT 1081.560 869.390 1081.820 869.710 ;
        RECT 1082.940 869.390 1083.200 869.710 ;
        RECT 1083.000 835.370 1083.140 869.390 ;
        RECT 1082.020 835.050 1082.280 835.370 ;
        RECT 1082.940 835.050 1083.200 835.370 ;
        RECT 1082.080 834.770 1082.220 835.050 ;
        RECT 1082.080 834.630 1082.680 834.770 ;
        RECT 1082.540 821.090 1082.680 834.630 ;
        RECT 1082.480 820.770 1082.740 821.090 ;
        RECT 1082.480 786.430 1082.740 786.750 ;
        RECT 1082.540 772.890 1082.680 786.430 ;
        RECT 1082.540 772.750 1083.140 772.890 ;
        RECT 1083.000 738.470 1083.140 772.750 ;
        RECT 1082.020 738.210 1082.280 738.470 ;
        RECT 1082.020 738.150 1082.680 738.210 ;
        RECT 1082.940 738.150 1083.200 738.470 ;
        RECT 1082.080 738.070 1082.680 738.150 ;
        RECT 1082.540 724.530 1082.680 738.070 ;
        RECT 1082.480 724.210 1082.740 724.530 ;
        RECT 1082.480 689.530 1082.740 689.850 ;
        RECT 1082.540 676.330 1082.680 689.530 ;
        RECT 1082.540 676.190 1083.140 676.330 ;
        RECT 1083.000 641.910 1083.140 676.190 ;
        RECT 1082.020 641.650 1082.280 641.910 ;
        RECT 1082.940 641.650 1083.200 641.910 ;
        RECT 1082.020 641.590 1083.200 641.650 ;
        RECT 1082.080 641.510 1083.140 641.590 ;
        RECT 1083.000 593.970 1083.140 641.510 ;
        RECT 1082.940 593.650 1083.200 593.970 ;
        RECT 1082.480 579.710 1082.740 580.030 ;
        RECT 1082.540 545.770 1082.680 579.710 ;
        RECT 1082.080 545.630 1082.680 545.770 ;
        RECT 1082.080 545.090 1082.220 545.630 ;
        RECT 1082.080 544.950 1082.680 545.090 ;
        RECT 1082.540 531.410 1082.680 544.950 ;
        RECT 1082.480 531.090 1082.740 531.410 ;
        RECT 1082.480 496.410 1082.740 496.730 ;
        RECT 1082.540 483.210 1082.680 496.410 ;
        RECT 1082.540 483.070 1083.140 483.210 ;
        RECT 1083.000 448.790 1083.140 483.070 ;
        RECT 1082.020 448.530 1082.280 448.790 ;
        RECT 1082.020 448.470 1082.680 448.530 ;
        RECT 1082.940 448.470 1083.200 448.790 ;
        RECT 1082.080 448.390 1082.680 448.470 ;
        RECT 1082.540 434.850 1082.680 448.390 ;
        RECT 1082.480 434.530 1082.740 434.850 ;
        RECT 1082.940 386.250 1083.200 386.570 ;
        RECT 1083.000 351.290 1083.140 386.250 ;
        RECT 1082.540 351.150 1083.140 351.290 ;
        RECT 1082.540 303.690 1082.680 351.150 ;
        RECT 1082.540 303.550 1083.140 303.690 ;
        RECT 1083.000 289.670 1083.140 303.550 ;
        RECT 1082.940 289.350 1083.200 289.670 ;
        RECT 1082.480 241.410 1082.740 241.730 ;
        RECT 1082.540 207.130 1082.680 241.410 ;
        RECT 1082.540 206.990 1083.140 207.130 ;
        RECT 1083.000 158.850 1083.140 206.990 ;
        RECT 1082.080 158.710 1083.140 158.850 ;
        RECT 1082.080 158.170 1082.220 158.710 ;
        RECT 1082.080 158.030 1082.680 158.170 ;
        RECT 1082.540 62.290 1082.680 158.030 ;
        RECT 1082.080 62.150 1082.680 62.290 ;
        RECT 1082.080 15.290 1082.220 62.150 ;
        RECT 1079.260 14.970 1079.520 15.290 ;
        RECT 1082.020 14.970 1082.280 15.290 ;
        RECT 1079.320 2.400 1079.460 14.970 ;
        RECT 1079.110 -4.800 1079.670 2.400 ;
      LAYER via2 ;
        RECT 1772.010 2023.880 1772.290 2024.160 ;
        RECT 1081.550 917.520 1081.830 917.800 ;
        RECT 1082.470 917.520 1082.750 917.800 ;
      LAYER met3 ;
        RECT 1755.835 2024.170 1759.835 2024.175 ;
        RECT 1771.985 2024.170 1772.315 2024.185 ;
        RECT 1755.835 2023.870 1772.315 2024.170 ;
        RECT 1755.835 2023.575 1759.835 2023.870 ;
        RECT 1771.985 2023.855 1772.315 2023.870 ;
        RECT 1081.525 917.810 1081.855 917.825 ;
        RECT 1082.445 917.810 1082.775 917.825 ;
        RECT 1081.525 917.510 1082.775 917.810 ;
        RECT 1081.525 917.495 1081.855 917.510 ;
        RECT 1082.445 917.495 1082.775 917.510 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 702.030 2386.360 702.350 2386.420 ;
        RECT 1080.150 2386.360 1080.470 2386.420 ;
        RECT 702.030 2386.220 1080.470 2386.360 ;
        RECT 702.030 2386.160 702.350 2386.220 ;
        RECT 1080.150 2386.160 1080.470 2386.220 ;
        RECT 702.030 31.180 702.350 31.240 ;
        RECT 1096.250 31.180 1096.570 31.240 ;
        RECT 702.030 31.040 1096.570 31.180 ;
        RECT 702.030 30.980 702.350 31.040 ;
        RECT 1096.250 30.980 1096.570 31.040 ;
      LAYER via ;
        RECT 702.060 2386.160 702.320 2386.420 ;
        RECT 1080.180 2386.160 1080.440 2386.420 ;
        RECT 702.060 30.980 702.320 31.240 ;
        RECT 1096.280 30.980 1096.540 31.240 ;
      LAYER met2 ;
        RECT 702.060 2386.130 702.320 2386.450 ;
        RECT 1080.180 2386.130 1080.440 2386.450 ;
        RECT 702.120 1393.845 702.260 2386.130 ;
        RECT 1080.240 2377.880 1080.380 2386.130 ;
        RECT 1080.220 2373.880 1080.500 2377.880 ;
        RECT 702.050 1393.475 702.330 1393.845 ;
        RECT 702.050 1392.115 702.330 1392.485 ;
        RECT 702.120 31.270 702.260 1392.115 ;
        RECT 702.060 30.950 702.320 31.270 ;
        RECT 1096.280 30.950 1096.540 31.270 ;
        RECT 1096.340 20.130 1096.480 30.950 ;
        RECT 1096.340 19.990 1096.940 20.130 ;
        RECT 1096.800 2.400 1096.940 19.990 ;
        RECT 1096.590 -4.800 1097.150 2.400 ;
      LAYER via2 ;
        RECT 702.050 1393.520 702.330 1393.800 ;
        RECT 702.050 1392.160 702.330 1392.440 ;
      LAYER met3 ;
        RECT 702.025 1393.810 702.355 1393.825 ;
        RECT 702.025 1393.495 702.570 1393.810 ;
        RECT 702.270 1392.465 702.570 1393.495 ;
        RECT 702.025 1392.150 702.570 1392.465 ;
        RECT 702.025 1392.135 702.355 1392.150 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 692.830 61.440 693.150 61.500 ;
        RECT 693.750 61.440 694.070 61.500 ;
        RECT 692.830 61.300 694.070 61.440 ;
        RECT 692.830 61.240 693.150 61.300 ;
        RECT 693.750 61.240 694.070 61.300 ;
        RECT 693.750 16.220 694.070 16.280 ;
        RECT 1114.650 16.220 1114.970 16.280 ;
        RECT 693.750 16.080 1114.970 16.220 ;
        RECT 693.750 16.020 694.070 16.080 ;
        RECT 1114.650 16.020 1114.970 16.080 ;
      LAYER via ;
        RECT 692.860 61.240 693.120 61.500 ;
        RECT 693.780 61.240 694.040 61.500 ;
        RECT 693.780 16.020 694.040 16.280 ;
        RECT 1114.680 16.020 1114.940 16.280 ;
      LAYER met2 ;
        RECT 692.850 1968.075 693.130 1968.445 ;
        RECT 692.920 1393.845 693.060 1968.075 ;
        RECT 692.850 1393.475 693.130 1393.845 ;
        RECT 692.850 1392.115 693.130 1392.485 ;
        RECT 692.920 61.530 693.060 1392.115 ;
        RECT 692.860 61.210 693.120 61.530 ;
        RECT 693.780 61.210 694.040 61.530 ;
        RECT 693.840 16.310 693.980 61.210 ;
        RECT 693.780 15.990 694.040 16.310 ;
        RECT 1114.680 15.990 1114.940 16.310 ;
        RECT 1114.740 2.400 1114.880 15.990 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
      LAYER via2 ;
        RECT 692.850 1968.120 693.130 1968.400 ;
        RECT 692.850 1393.520 693.130 1393.800 ;
        RECT 692.850 1392.160 693.130 1392.440 ;
      LAYER met3 ;
        RECT 692.825 1968.410 693.155 1968.425 ;
        RECT 715.810 1968.410 719.810 1968.415 ;
        RECT 692.825 1968.110 719.810 1968.410 ;
        RECT 692.825 1968.095 693.155 1968.110 ;
        RECT 715.810 1967.815 719.810 1968.110 ;
        RECT 692.825 1393.810 693.155 1393.825 ;
        RECT 692.825 1393.495 693.370 1393.810 ;
        RECT 693.070 1392.465 693.370 1393.495 ;
        RECT 692.825 1392.150 693.370 1392.465 ;
        RECT 692.825 1392.135 693.155 1392.150 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1755.505 1331.525 1756.135 1331.695 ;
        RECT 1755.505 1310.105 1755.675 1331.525 ;
      LAYER mcon ;
        RECT 1755.965 1331.525 1756.135 1331.695 ;
      LAYER met1 ;
        RECT 1754.510 1487.060 1754.830 1487.120 ;
        RECT 1759.110 1487.060 1759.430 1487.120 ;
        RECT 1754.510 1486.920 1759.430 1487.060 ;
        RECT 1754.510 1486.860 1754.830 1486.920 ;
        RECT 1759.110 1486.860 1759.430 1486.920 ;
        RECT 1752.670 1333.380 1752.990 1333.440 ;
        RECT 1755.890 1333.380 1756.210 1333.440 ;
        RECT 1752.670 1333.240 1756.210 1333.380 ;
        RECT 1752.670 1333.180 1752.990 1333.240 ;
        RECT 1755.890 1333.180 1756.210 1333.240 ;
        RECT 1755.890 1331.680 1756.210 1331.740 ;
        RECT 1755.890 1331.540 1756.405 1331.680 ;
        RECT 1755.890 1331.480 1756.210 1331.540 ;
        RECT 1138.110 1310.260 1138.430 1310.320 ;
        RECT 1755.445 1310.260 1755.735 1310.305 ;
        RECT 1138.110 1310.120 1755.735 1310.260 ;
        RECT 1138.110 1310.060 1138.430 1310.120 ;
        RECT 1755.445 1310.075 1755.735 1310.120 ;
        RECT 1132.590 20.640 1132.910 20.700 ;
        RECT 1138.110 20.640 1138.430 20.700 ;
        RECT 1132.590 20.500 1138.430 20.640 ;
        RECT 1132.590 20.440 1132.910 20.500 ;
        RECT 1138.110 20.440 1138.430 20.500 ;
      LAYER via ;
        RECT 1754.540 1486.860 1754.800 1487.120 ;
        RECT 1759.140 1486.860 1759.400 1487.120 ;
        RECT 1752.700 1333.180 1752.960 1333.440 ;
        RECT 1755.920 1333.180 1756.180 1333.440 ;
        RECT 1755.920 1331.480 1756.180 1331.740 ;
        RECT 1138.140 1310.060 1138.400 1310.320 ;
        RECT 1132.620 20.440 1132.880 20.700 ;
        RECT 1138.140 20.440 1138.400 20.700 ;
      LAYER met2 ;
        RECT 1759.130 1516.555 1759.410 1516.925 ;
        RECT 1759.200 1487.150 1759.340 1516.555 ;
        RECT 1754.540 1486.830 1754.800 1487.150 ;
        RECT 1759.140 1486.830 1759.400 1487.150 ;
        RECT 1754.600 1484.850 1754.740 1486.830 ;
        RECT 1752.760 1484.710 1754.740 1484.850 ;
        RECT 1752.760 1333.470 1752.900 1484.710 ;
        RECT 1752.700 1333.150 1752.960 1333.470 ;
        RECT 1755.920 1333.150 1756.180 1333.470 ;
        RECT 1755.980 1331.770 1756.120 1333.150 ;
        RECT 1755.920 1331.450 1756.180 1331.770 ;
        RECT 1138.140 1310.030 1138.400 1310.350 ;
        RECT 1138.200 20.730 1138.340 1310.030 ;
        RECT 1132.620 20.410 1132.880 20.730 ;
        RECT 1138.140 20.410 1138.400 20.730 ;
        RECT 1132.680 2.400 1132.820 20.410 ;
        RECT 1132.470 -4.800 1133.030 2.400 ;
      LAYER via2 ;
        RECT 1759.130 1516.600 1759.410 1516.880 ;
      LAYER met3 ;
        RECT 1755.835 1519.015 1759.835 1519.615 ;
        RECT 1759.350 1516.905 1759.650 1519.015 ;
        RECT 1759.105 1516.890 1759.650 1516.905 ;
        RECT 1758.700 1516.590 1759.650 1516.890 ;
        RECT 1759.105 1516.575 1759.435 1516.590 ;
    END
  END la_data_in[28]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 668.910 2049.420 669.230 2049.480 ;
        RECT 706.170 2049.420 706.490 2049.480 ;
        RECT 668.910 2049.280 706.490 2049.420 ;
        RECT 668.910 2049.220 669.230 2049.280 ;
        RECT 706.170 2049.220 706.490 2049.280 ;
      LAYER via ;
        RECT 668.940 2049.220 669.200 2049.480 ;
        RECT 706.200 2049.220 706.460 2049.480 ;
      LAYER met2 ;
        RECT 706.190 2053.755 706.470 2054.125 ;
        RECT 706.260 2049.510 706.400 2053.755 ;
        RECT 668.940 2049.190 669.200 2049.510 ;
        RECT 706.200 2049.190 706.460 2049.510 ;
        RECT 669.000 2.400 669.140 2049.190 ;
        RECT 668.790 -4.800 669.350 2.400 ;
      LAYER via2 ;
        RECT 706.190 2053.800 706.470 2054.080 ;
      LAYER met3 ;
        RECT 706.165 2054.090 706.495 2054.105 ;
        RECT 715.810 2054.090 719.810 2054.095 ;
        RECT 706.165 2053.790 719.810 2054.090 ;
        RECT 706.165 2053.775 706.495 2053.790 ;
        RECT 715.810 2053.495 719.810 2053.790 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1030.470 1311.280 1030.790 1311.340 ;
        RECT 1034.610 1311.280 1034.930 1311.340 ;
        RECT 1030.470 1311.140 1034.930 1311.280 ;
        RECT 1030.470 1311.080 1030.790 1311.140 ;
        RECT 1034.610 1311.080 1034.930 1311.140 ;
        RECT 1034.610 23.700 1034.930 23.760 ;
        RECT 1168.470 23.700 1168.790 23.760 ;
        RECT 1034.610 23.560 1168.790 23.700 ;
        RECT 1034.610 23.500 1034.930 23.560 ;
        RECT 1168.470 23.500 1168.790 23.560 ;
      LAYER via ;
        RECT 1030.500 1311.080 1030.760 1311.340 ;
        RECT 1034.640 1311.080 1034.900 1311.340 ;
        RECT 1034.640 23.500 1034.900 23.760 ;
        RECT 1168.500 23.500 1168.760 23.760 ;
      LAYER met2 ;
        RECT 1030.540 1323.135 1030.820 1327.135 ;
        RECT 1030.560 1311.370 1030.700 1323.135 ;
        RECT 1030.500 1311.050 1030.760 1311.370 ;
        RECT 1034.640 1311.050 1034.900 1311.370 ;
        RECT 1034.700 23.790 1034.840 1311.050 ;
        RECT 1034.640 23.470 1034.900 23.790 ;
        RECT 1168.500 23.470 1168.760 23.790 ;
        RECT 1168.560 2.400 1168.700 23.470 ;
        RECT 1168.350 -4.800 1168.910 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1761.870 1341.540 1762.190 1341.600 ;
        RECT 1764.170 1341.540 1764.490 1341.600 ;
        RECT 1761.870 1341.400 1764.490 1341.540 ;
        RECT 1761.870 1341.340 1762.190 1341.400 ;
        RECT 1764.170 1341.340 1764.490 1341.400 ;
        RECT 1185.950 1310.600 1186.270 1310.660 ;
        RECT 1764.170 1310.600 1764.490 1310.660 ;
        RECT 1185.950 1310.460 1764.490 1310.600 ;
        RECT 1185.950 1310.400 1186.270 1310.460 ;
        RECT 1764.170 1310.400 1764.490 1310.460 ;
      LAYER via ;
        RECT 1761.900 1341.340 1762.160 1341.600 ;
        RECT 1764.200 1341.340 1764.460 1341.600 ;
        RECT 1185.980 1310.400 1186.240 1310.660 ;
        RECT 1764.200 1310.400 1764.460 1310.660 ;
      LAYER met2 ;
        RECT 1761.890 2331.195 1762.170 2331.565 ;
        RECT 1761.960 1341.630 1762.100 2331.195 ;
        RECT 1761.900 1341.310 1762.160 1341.630 ;
        RECT 1764.200 1341.310 1764.460 1341.630 ;
        RECT 1764.260 1310.690 1764.400 1341.310 ;
        RECT 1185.980 1310.370 1186.240 1310.690 ;
        RECT 1764.200 1310.370 1764.460 1310.690 ;
        RECT 1186.040 2.400 1186.180 1310.370 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
      LAYER via2 ;
        RECT 1761.890 2331.240 1762.170 2331.520 ;
      LAYER met3 ;
        RECT 1755.835 2331.530 1759.835 2331.535 ;
        RECT 1761.865 2331.530 1762.195 2331.545 ;
        RECT 1755.835 2331.230 1762.195 2331.530 ;
        RECT 1755.835 2330.935 1759.835 2331.230 ;
        RECT 1761.865 2331.215 1762.195 2331.230 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1768.770 1745.800 1769.090 1745.860 ;
        RECT 1783.490 1745.800 1783.810 1745.860 ;
        RECT 1768.770 1745.660 1783.810 1745.800 ;
        RECT 1768.770 1745.600 1769.090 1745.660 ;
        RECT 1783.490 1745.600 1783.810 1745.660 ;
        RECT 1207.110 1323.180 1207.430 1323.240 ;
        RECT 1783.490 1323.180 1783.810 1323.240 ;
        RECT 1207.110 1323.040 1783.810 1323.180 ;
        RECT 1207.110 1322.980 1207.430 1323.040 ;
        RECT 1783.490 1322.980 1783.810 1323.040 ;
        RECT 1203.890 16.560 1204.210 16.620 ;
        RECT 1207.110 16.560 1207.430 16.620 ;
        RECT 1203.890 16.420 1207.430 16.560 ;
        RECT 1203.890 16.360 1204.210 16.420 ;
        RECT 1207.110 16.360 1207.430 16.420 ;
      LAYER via ;
        RECT 1768.800 1745.600 1769.060 1745.860 ;
        RECT 1783.520 1745.600 1783.780 1745.860 ;
        RECT 1207.140 1322.980 1207.400 1323.240 ;
        RECT 1783.520 1322.980 1783.780 1323.240 ;
        RECT 1203.920 16.360 1204.180 16.620 ;
        RECT 1207.140 16.360 1207.400 16.620 ;
      LAYER met2 ;
        RECT 1768.790 1749.115 1769.070 1749.485 ;
        RECT 1768.860 1745.890 1769.000 1749.115 ;
        RECT 1768.800 1745.570 1769.060 1745.890 ;
        RECT 1783.520 1745.570 1783.780 1745.890 ;
        RECT 1783.580 1323.270 1783.720 1745.570 ;
        RECT 1207.140 1322.950 1207.400 1323.270 ;
        RECT 1783.520 1322.950 1783.780 1323.270 ;
        RECT 1207.200 16.650 1207.340 1322.950 ;
        RECT 1203.920 16.330 1204.180 16.650 ;
        RECT 1207.140 16.330 1207.400 16.650 ;
        RECT 1203.980 2.400 1204.120 16.330 ;
        RECT 1203.770 -4.800 1204.330 2.400 ;
      LAYER via2 ;
        RECT 1768.790 1749.160 1769.070 1749.440 ;
      LAYER met3 ;
        RECT 1755.835 1749.450 1759.835 1749.455 ;
        RECT 1768.765 1749.450 1769.095 1749.465 ;
        RECT 1755.835 1749.150 1769.095 1749.450 ;
        RECT 1755.835 1748.855 1759.835 1749.150 ;
        RECT 1768.765 1749.135 1769.095 1749.150 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 699.805 1368.925 699.975 1393.575 ;
      LAYER mcon ;
        RECT 699.805 1393.405 699.975 1393.575 ;
      LAYER met1 ;
        RECT 699.730 1393.560 700.050 1393.620 ;
        RECT 699.730 1393.420 700.245 1393.560 ;
        RECT 699.730 1393.360 700.050 1393.420 ;
        RECT 699.730 1369.080 700.050 1369.140 ;
        RECT 699.535 1368.940 700.050 1369.080 ;
        RECT 699.730 1368.880 700.050 1368.940 ;
        RECT 699.730 16.560 700.050 16.620 ;
        RECT 699.730 16.420 1197.680 16.560 ;
        RECT 699.730 16.360 700.050 16.420 ;
        RECT 1197.540 16.220 1197.680 16.420 ;
        RECT 1221.830 16.220 1222.150 16.280 ;
        RECT 1197.540 16.080 1222.150 16.220 ;
        RECT 1221.830 16.020 1222.150 16.080 ;
      LAYER via ;
        RECT 699.760 1393.360 700.020 1393.620 ;
        RECT 699.760 1368.880 700.020 1369.140 ;
        RECT 699.760 16.360 700.020 16.620 ;
        RECT 1221.860 16.020 1222.120 16.280 ;
      LAYER met2 ;
        RECT 699.750 1421.355 700.030 1421.725 ;
        RECT 699.820 1393.650 699.960 1421.355 ;
        RECT 699.760 1393.330 700.020 1393.650 ;
        RECT 699.760 1368.850 700.020 1369.170 ;
        RECT 699.820 16.650 699.960 1368.850 ;
        RECT 699.760 16.330 700.020 16.650 ;
        RECT 1221.860 15.990 1222.120 16.310 ;
        RECT 1221.920 2.400 1222.060 15.990 ;
        RECT 1221.710 -4.800 1222.270 2.400 ;
      LAYER via2 ;
        RECT 699.750 1421.400 700.030 1421.680 ;
      LAYER met3 ;
        RECT 699.725 1421.690 700.055 1421.705 ;
        RECT 715.810 1421.690 719.810 1421.695 ;
        RECT 699.725 1421.390 719.810 1421.690 ;
        RECT 699.725 1421.375 700.055 1421.390 ;
        RECT 715.810 1421.095 719.810 1421.390 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1751.365 724.625 1751.535 814.215 ;
        RECT 1242.145 14.705 1242.315 15.555 ;
        RECT 1269.745 14.705 1269.915 16.915 ;
        RECT 1417.865 15.385 1418.035 16.915 ;
        RECT 1704.905 16.575 1705.075 20.655 ;
        RECT 1441.785 15.385 1441.955 16.235 ;
        RECT 1497.445 15.385 1497.615 16.235 ;
        RECT 1538.845 15.385 1539.015 16.235 ;
        RECT 1655.685 15.385 1655.855 16.575 ;
        RECT 1704.445 16.405 1705.075 16.575 ;
      LAYER mcon ;
        RECT 1751.365 814.045 1751.535 814.215 ;
        RECT 1704.905 20.485 1705.075 20.655 ;
        RECT 1269.745 16.745 1269.915 16.915 ;
        RECT 1242.145 15.385 1242.315 15.555 ;
        RECT 1417.865 16.745 1418.035 16.915 ;
        RECT 1655.685 16.405 1655.855 16.575 ;
        RECT 1441.785 16.065 1441.955 16.235 ;
        RECT 1497.445 16.065 1497.615 16.235 ;
        RECT 1538.845 16.065 1539.015 16.235 ;
      LAYER met1 ;
        RECT 1751.290 1325.560 1751.610 1325.620 ;
        RECT 1770.610 1325.560 1770.930 1325.620 ;
        RECT 1751.290 1325.420 1770.930 1325.560 ;
        RECT 1751.290 1325.360 1751.610 1325.420 ;
        RECT 1770.610 1325.360 1770.930 1325.420 ;
        RECT 1751.290 814.200 1751.610 814.260 ;
        RECT 1751.095 814.060 1751.610 814.200 ;
        RECT 1751.290 814.000 1751.610 814.060 ;
        RECT 1751.290 724.780 1751.610 724.840 ;
        RECT 1751.095 724.640 1751.610 724.780 ;
        RECT 1751.290 724.580 1751.610 724.640 ;
        RECT 1704.845 20.640 1705.135 20.685 ;
        RECT 1749.910 20.640 1750.230 20.700 ;
        RECT 1704.845 20.500 1750.230 20.640 ;
        RECT 1704.845 20.455 1705.135 20.500 ;
        RECT 1749.910 20.440 1750.230 20.500 ;
        RECT 1269.685 16.900 1269.975 16.945 ;
        RECT 1417.805 16.900 1418.095 16.945 ;
        RECT 1269.685 16.760 1365.580 16.900 ;
        RECT 1269.685 16.715 1269.975 16.760 ;
        RECT 1365.440 16.560 1365.580 16.760 ;
        RECT 1366.360 16.760 1418.095 16.900 ;
        RECT 1366.360 16.560 1366.500 16.760 ;
        RECT 1417.805 16.715 1418.095 16.760 ;
        RECT 1655.625 16.560 1655.915 16.605 ;
        RECT 1704.385 16.560 1704.675 16.605 ;
        RECT 1365.440 16.420 1366.500 16.560 ;
        RECT 1586.700 16.420 1618.120 16.560 ;
        RECT 1441.725 16.220 1442.015 16.265 ;
        RECT 1497.385 16.220 1497.675 16.265 ;
        RECT 1441.725 16.080 1497.675 16.220 ;
        RECT 1441.725 16.035 1442.015 16.080 ;
        RECT 1497.385 16.035 1497.675 16.080 ;
        RECT 1538.785 16.220 1539.075 16.265 ;
        RECT 1586.700 16.220 1586.840 16.420 ;
        RECT 1538.785 16.080 1586.840 16.220 ;
        RECT 1538.785 16.035 1539.075 16.080 ;
        RECT 1239.770 15.540 1240.090 15.600 ;
        RECT 1242.085 15.540 1242.375 15.585 ;
        RECT 1239.770 15.400 1242.375 15.540 ;
        RECT 1239.770 15.340 1240.090 15.400 ;
        RECT 1242.085 15.355 1242.375 15.400 ;
        RECT 1417.805 15.540 1418.095 15.585 ;
        RECT 1441.725 15.540 1442.015 15.585 ;
        RECT 1417.805 15.400 1442.015 15.540 ;
        RECT 1417.805 15.355 1418.095 15.400 ;
        RECT 1441.725 15.355 1442.015 15.400 ;
        RECT 1497.385 15.540 1497.675 15.585 ;
        RECT 1538.785 15.540 1539.075 15.585 ;
        RECT 1497.385 15.400 1539.075 15.540 ;
        RECT 1617.980 15.540 1618.120 16.420 ;
        RECT 1655.625 16.420 1704.675 16.560 ;
        RECT 1655.625 16.375 1655.915 16.420 ;
        RECT 1704.385 16.375 1704.675 16.420 ;
        RECT 1655.625 15.540 1655.915 15.585 ;
        RECT 1617.980 15.400 1655.915 15.540 ;
        RECT 1497.385 15.355 1497.675 15.400 ;
        RECT 1538.785 15.355 1539.075 15.400 ;
        RECT 1655.625 15.355 1655.915 15.400 ;
        RECT 1242.085 14.860 1242.375 14.905 ;
        RECT 1269.685 14.860 1269.975 14.905 ;
        RECT 1242.085 14.720 1269.975 14.860 ;
        RECT 1242.085 14.675 1242.375 14.720 ;
        RECT 1269.685 14.675 1269.975 14.720 ;
      LAYER via ;
        RECT 1751.320 1325.360 1751.580 1325.620 ;
        RECT 1770.640 1325.360 1770.900 1325.620 ;
        RECT 1751.320 814.000 1751.580 814.260 ;
        RECT 1751.320 724.580 1751.580 724.840 ;
        RECT 1749.940 20.440 1750.200 20.700 ;
        RECT 1239.800 15.340 1240.060 15.600 ;
      LAYER met2 ;
        RECT 1770.630 2125.835 1770.910 2126.205 ;
        RECT 1770.700 1325.650 1770.840 2125.835 ;
        RECT 1751.320 1325.330 1751.580 1325.650 ;
        RECT 1770.640 1325.330 1770.900 1325.650 ;
        RECT 1751.380 814.290 1751.520 1325.330 ;
        RECT 1751.320 813.970 1751.580 814.290 ;
        RECT 1751.320 724.550 1751.580 724.870 ;
        RECT 1751.380 71.810 1751.520 724.550 ;
        RECT 1750.000 71.670 1751.520 71.810 ;
        RECT 1750.000 20.730 1750.140 71.670 ;
        RECT 1749.940 20.410 1750.200 20.730 ;
        RECT 1239.800 15.310 1240.060 15.630 ;
        RECT 1239.860 2.400 1240.000 15.310 ;
        RECT 1239.650 -4.800 1240.210 2.400 ;
      LAYER via2 ;
        RECT 1770.630 2125.880 1770.910 2126.160 ;
      LAYER met3 ;
        RECT 1755.835 2126.170 1759.835 2126.175 ;
        RECT 1770.605 2126.170 1770.935 2126.185 ;
        RECT 1755.835 2125.870 1770.935 2126.170 ;
        RECT 1755.835 2125.575 1759.835 2125.870 ;
        RECT 1770.605 2125.855 1770.935 2125.870 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1261.925 1322.685 1262.095 1329.995 ;
        RECT 1751.825 1329.825 1751.995 1333.395 ;
      LAYER mcon ;
        RECT 1751.825 1333.225 1751.995 1333.395 ;
        RECT 1261.925 1329.825 1262.095 1329.995 ;
      LAYER met1 ;
        RECT 1751.750 1333.380 1752.070 1333.440 ;
        RECT 1751.555 1333.240 1752.070 1333.380 ;
        RECT 1751.750 1333.180 1752.070 1333.240 ;
        RECT 1261.865 1329.980 1262.155 1330.025 ;
        RECT 1751.765 1329.980 1752.055 1330.025 ;
        RECT 1261.865 1329.840 1752.055 1329.980 ;
        RECT 1261.865 1329.795 1262.155 1329.840 ;
        RECT 1751.765 1329.795 1752.055 1329.840 ;
        RECT 1261.850 1322.840 1262.170 1322.900 ;
        RECT 1261.655 1322.700 1262.170 1322.840 ;
        RECT 1261.850 1322.640 1262.170 1322.700 ;
        RECT 1257.250 17.920 1257.570 17.980 ;
        RECT 1261.850 17.920 1262.170 17.980 ;
        RECT 1257.250 17.780 1262.170 17.920 ;
        RECT 1257.250 17.720 1257.570 17.780 ;
        RECT 1261.850 17.720 1262.170 17.780 ;
      LAYER via ;
        RECT 1751.780 1333.180 1752.040 1333.440 ;
        RECT 1261.880 1322.640 1262.140 1322.900 ;
        RECT 1257.280 17.720 1257.540 17.980 ;
        RECT 1261.880 17.720 1262.140 17.980 ;
      LAYER met2 ;
        RECT 1438.970 2379.475 1439.250 2379.845 ;
        RECT 1439.040 2377.880 1439.180 2379.475 ;
        RECT 1439.020 2373.880 1439.300 2377.880 ;
        RECT 1751.770 2371.315 1752.050 2371.685 ;
        RECT 1751.840 1333.470 1751.980 2371.315 ;
        RECT 1751.780 1333.150 1752.040 1333.470 ;
        RECT 1261.880 1322.610 1262.140 1322.930 ;
        RECT 1261.940 18.010 1262.080 1322.610 ;
        RECT 1257.280 17.690 1257.540 18.010 ;
        RECT 1261.880 17.690 1262.140 18.010 ;
        RECT 1257.340 2.400 1257.480 17.690 ;
        RECT 1257.130 -4.800 1257.690 2.400 ;
      LAYER via2 ;
        RECT 1438.970 2379.520 1439.250 2379.800 ;
        RECT 1751.770 2371.360 1752.050 2371.640 ;
      LAYER met3 ;
        RECT 1438.945 2379.820 1439.275 2379.825 ;
        RECT 1438.945 2379.810 1439.530 2379.820 ;
        RECT 1438.945 2379.510 1439.730 2379.810 ;
        RECT 1438.945 2379.500 1439.530 2379.510 ;
        RECT 1438.945 2379.495 1439.275 2379.500 ;
        RECT 1439.150 2371.650 1439.530 2371.660 ;
        RECT 1751.745 2371.650 1752.075 2371.665 ;
        RECT 1439.150 2371.350 1752.075 2371.650 ;
        RECT 1439.150 2371.340 1439.530 2371.350 ;
        RECT 1751.745 2371.335 1752.075 2371.350 ;
      LAYER via3 ;
        RECT 1439.180 2379.500 1439.500 2379.820 ;
        RECT 1439.180 2371.340 1439.500 2371.660 ;
      LAYER met4 ;
        RECT 1439.175 2379.495 1439.505 2379.825 ;
        RECT 1439.190 2371.665 1439.490 2379.495 ;
        RECT 1439.175 2371.335 1439.505 2371.665 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 734.765 19.125 734.935 20.995 ;
        RECT 786.745 18.105 786.915 20.655 ;
        RECT 793.185 18.445 794.275 18.615 ;
        RECT 793.185 18.105 793.355 18.445 ;
        RECT 794.105 14.705 794.275 18.445 ;
        RECT 855.285 14.365 855.455 20.655 ;
        RECT 883.345 14.705 883.515 20.655 ;
        RECT 959.245 14.705 959.415 15.895 ;
        RECT 983.165 14.705 983.335 15.555 ;
        RECT 1014.445 14.365 1014.615 15.555 ;
        RECT 1062.285 14.365 1062.455 15.895 ;
        RECT 1100.465 15.725 1100.635 20.655 ;
        RECT 1152.445 15.725 1152.615 20.315 ;
        RECT 1193.385 15.725 1193.555 20.655 ;
      LAYER mcon ;
        RECT 734.765 20.825 734.935 20.995 ;
        RECT 786.745 20.485 786.915 20.655 ;
        RECT 855.285 20.485 855.455 20.655 ;
        RECT 883.345 20.485 883.515 20.655 ;
        RECT 1100.465 20.485 1100.635 20.655 ;
        RECT 1193.385 20.485 1193.555 20.655 ;
        RECT 959.245 15.725 959.415 15.895 ;
        RECT 1062.285 15.725 1062.455 15.895 ;
        RECT 1152.445 20.145 1152.615 20.315 ;
        RECT 983.165 15.385 983.335 15.555 ;
        RECT 1014.445 15.385 1014.615 15.555 ;
      LAYER met1 ;
        RECT 694.670 2189.500 694.990 2189.560 ;
        RECT 707.550 2189.500 707.870 2189.560 ;
        RECT 694.670 2189.360 707.870 2189.500 ;
        RECT 694.670 2189.300 694.990 2189.360 ;
        RECT 707.550 2189.300 707.870 2189.360 ;
        RECT 734.705 20.980 734.995 21.025 ;
        RECT 734.705 20.840 770.340 20.980 ;
        RECT 734.705 20.795 734.995 20.840 ;
        RECT 770.200 20.300 770.340 20.840 ;
        RECT 786.300 20.840 786.900 20.980 ;
        RECT 786.300 20.300 786.440 20.840 ;
        RECT 786.760 20.685 786.900 20.840 ;
        RECT 786.685 20.455 786.975 20.685 ;
        RECT 855.225 20.640 855.515 20.685 ;
        RECT 883.285 20.640 883.575 20.685 ;
        RECT 855.225 20.500 883.575 20.640 ;
        RECT 855.225 20.455 855.515 20.500 ;
        RECT 883.285 20.455 883.575 20.500 ;
        RECT 1100.405 20.640 1100.695 20.685 ;
        RECT 1193.325 20.640 1193.615 20.685 ;
        RECT 1275.190 20.640 1275.510 20.700 ;
        RECT 1100.405 20.500 1132.360 20.640 ;
        RECT 1100.405 20.455 1100.695 20.500 ;
        RECT 770.200 20.160 786.440 20.300 ;
        RECT 1132.220 20.300 1132.360 20.500 ;
        RECT 1193.325 20.500 1275.510 20.640 ;
        RECT 1193.325 20.455 1193.615 20.500 ;
        RECT 1275.190 20.440 1275.510 20.500 ;
        RECT 1152.385 20.300 1152.675 20.345 ;
        RECT 1132.220 20.160 1152.675 20.300 ;
        RECT 1152.385 20.115 1152.675 20.160 ;
        RECT 694.670 19.280 694.990 19.340 ;
        RECT 734.705 19.280 734.995 19.325 ;
        RECT 694.670 19.140 734.995 19.280 ;
        RECT 694.670 19.080 694.990 19.140 ;
        RECT 734.705 19.095 734.995 19.140 ;
        RECT 786.685 18.260 786.975 18.305 ;
        RECT 793.125 18.260 793.415 18.305 ;
        RECT 786.685 18.120 793.415 18.260 ;
        RECT 786.685 18.075 786.975 18.120 ;
        RECT 793.125 18.075 793.415 18.120 ;
        RECT 959.185 15.880 959.475 15.925 ;
        RECT 926.600 15.740 959.475 15.880 ;
        RECT 794.045 14.860 794.335 14.905 ;
        RECT 883.285 14.860 883.575 14.905 ;
        RECT 926.600 14.860 926.740 15.740 ;
        RECT 959.185 15.695 959.475 15.740 ;
        RECT 1062.225 15.880 1062.515 15.925 ;
        RECT 1100.405 15.880 1100.695 15.925 ;
        RECT 1062.225 15.740 1100.695 15.880 ;
        RECT 1062.225 15.695 1062.515 15.740 ;
        RECT 1100.405 15.695 1100.695 15.740 ;
        RECT 1152.385 15.880 1152.675 15.925 ;
        RECT 1193.325 15.880 1193.615 15.925 ;
        RECT 1152.385 15.740 1193.615 15.880 ;
        RECT 1152.385 15.695 1152.675 15.740 ;
        RECT 1193.325 15.695 1193.615 15.740 ;
        RECT 983.105 15.540 983.395 15.585 ;
        RECT 1014.385 15.540 1014.675 15.585 ;
        RECT 983.105 15.400 1014.675 15.540 ;
        RECT 983.105 15.355 983.395 15.400 ;
        RECT 1014.385 15.355 1014.675 15.400 ;
        RECT 794.045 14.720 800.240 14.860 ;
        RECT 794.045 14.675 794.335 14.720 ;
        RECT 800.100 14.520 800.240 14.720 ;
        RECT 883.285 14.720 926.740 14.860 ;
        RECT 959.185 14.860 959.475 14.905 ;
        RECT 983.105 14.860 983.395 14.905 ;
        RECT 959.185 14.720 983.395 14.860 ;
        RECT 883.285 14.675 883.575 14.720 ;
        RECT 959.185 14.675 959.475 14.720 ;
        RECT 983.105 14.675 983.395 14.720 ;
        RECT 855.225 14.520 855.515 14.565 ;
        RECT 800.100 14.380 855.515 14.520 ;
        RECT 855.225 14.335 855.515 14.380 ;
        RECT 1014.385 14.520 1014.675 14.565 ;
        RECT 1062.225 14.520 1062.515 14.565 ;
        RECT 1014.385 14.380 1062.515 14.520 ;
        RECT 1014.385 14.335 1014.675 14.380 ;
        RECT 1062.225 14.335 1062.515 14.380 ;
      LAYER via ;
        RECT 694.700 2189.300 694.960 2189.560 ;
        RECT 707.580 2189.300 707.840 2189.560 ;
        RECT 1275.220 20.440 1275.480 20.700 ;
        RECT 694.700 19.080 694.960 19.340 ;
      LAYER met2 ;
        RECT 707.570 2191.115 707.850 2191.485 ;
        RECT 707.640 2189.590 707.780 2191.115 ;
        RECT 694.700 2189.270 694.960 2189.590 ;
        RECT 707.580 2189.270 707.840 2189.590 ;
        RECT 694.760 1393.845 694.900 2189.270 ;
        RECT 694.690 1393.475 694.970 1393.845 ;
        RECT 694.690 1392.115 694.970 1392.485 ;
        RECT 694.760 19.370 694.900 1392.115 ;
        RECT 1275.220 20.410 1275.480 20.730 ;
        RECT 694.700 19.050 694.960 19.370 ;
        RECT 1275.280 2.400 1275.420 20.410 ;
        RECT 1275.070 -4.800 1275.630 2.400 ;
      LAYER via2 ;
        RECT 707.570 2191.160 707.850 2191.440 ;
        RECT 694.690 1393.520 694.970 1393.800 ;
        RECT 694.690 1392.160 694.970 1392.440 ;
      LAYER met3 ;
        RECT 707.545 2191.450 707.875 2191.465 ;
        RECT 715.810 2191.450 719.810 2191.455 ;
        RECT 707.545 2191.150 719.810 2191.450 ;
        RECT 707.545 2191.135 707.875 2191.150 ;
        RECT 715.810 2190.855 719.810 2191.150 ;
        RECT 694.665 1393.810 694.995 1393.825 ;
        RECT 694.665 1393.495 695.210 1393.810 ;
        RECT 694.910 1392.465 695.210 1393.495 ;
        RECT 694.665 1392.150 695.210 1392.465 ;
        RECT 694.665 1392.135 694.995 1392.150 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 689.150 2332.300 689.470 2332.360 ;
        RECT 709.390 2332.300 709.710 2332.360 ;
        RECT 689.150 2332.160 709.710 2332.300 ;
        RECT 689.150 2332.100 689.470 2332.160 ;
        RECT 709.390 2332.100 709.710 2332.160 ;
        RECT 689.150 19.620 689.470 19.680 ;
        RECT 1293.130 19.620 1293.450 19.680 ;
        RECT 689.150 19.480 1293.450 19.620 ;
        RECT 689.150 19.420 689.470 19.480 ;
        RECT 1293.130 19.420 1293.450 19.480 ;
      LAYER via ;
        RECT 689.180 2332.100 689.440 2332.360 ;
        RECT 709.420 2332.100 709.680 2332.360 ;
        RECT 689.180 19.420 689.440 19.680 ;
        RECT 1293.160 19.420 1293.420 19.680 ;
      LAYER met2 ;
        RECT 709.410 2335.275 709.690 2335.645 ;
        RECT 709.480 2332.390 709.620 2335.275 ;
        RECT 689.180 2332.070 689.440 2332.390 ;
        RECT 709.420 2332.070 709.680 2332.390 ;
        RECT 689.240 1393.845 689.380 2332.070 ;
        RECT 689.170 1393.475 689.450 1393.845 ;
        RECT 689.170 1392.115 689.450 1392.485 ;
        RECT 689.240 19.710 689.380 1392.115 ;
        RECT 689.180 19.390 689.440 19.710 ;
        RECT 1293.160 19.390 1293.420 19.710 ;
        RECT 1293.220 2.400 1293.360 19.390 ;
        RECT 1293.010 -4.800 1293.570 2.400 ;
      LAYER via2 ;
        RECT 709.410 2335.320 709.690 2335.600 ;
        RECT 689.170 1393.520 689.450 1393.800 ;
        RECT 689.170 1392.160 689.450 1392.440 ;
      LAYER met3 ;
        RECT 709.385 2335.610 709.715 2335.625 ;
        RECT 715.810 2335.610 719.810 2335.615 ;
        RECT 709.385 2335.310 719.810 2335.610 ;
        RECT 709.385 2335.295 709.715 2335.310 ;
        RECT 715.810 2335.015 719.810 2335.310 ;
        RECT 689.145 1393.810 689.475 1393.825 ;
        RECT 689.145 1393.495 689.690 1393.810 ;
        RECT 689.390 1392.465 689.690 1393.495 ;
        RECT 689.145 1392.150 689.690 1392.465 ;
        RECT 689.145 1392.135 689.475 1392.150 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1725.605 16.405 1725.775 19.295 ;
      LAYER mcon ;
        RECT 1725.605 19.125 1725.775 19.295 ;
      LAYER met1 ;
        RECT 1751.750 1325.220 1752.070 1325.280 ;
        RECT 1769.690 1325.220 1770.010 1325.280 ;
        RECT 1751.750 1325.080 1770.010 1325.220 ;
        RECT 1751.750 1325.020 1752.070 1325.080 ;
        RECT 1769.690 1325.020 1770.010 1325.080 ;
        RECT 1751.750 717.440 1752.070 717.700 ;
        RECT 1751.840 717.020 1751.980 717.440 ;
        RECT 1751.750 716.760 1752.070 717.020 ;
        RECT 1311.070 19.280 1311.390 19.340 ;
        RECT 1725.545 19.280 1725.835 19.325 ;
        RECT 1311.070 19.140 1725.835 19.280 ;
        RECT 1311.070 19.080 1311.390 19.140 ;
        RECT 1725.545 19.095 1725.835 19.140 ;
        RECT 1725.545 16.560 1725.835 16.605 ;
        RECT 1751.750 16.560 1752.070 16.620 ;
        RECT 1725.545 16.420 1752.070 16.560 ;
        RECT 1725.545 16.375 1725.835 16.420 ;
        RECT 1751.750 16.360 1752.070 16.420 ;
      LAYER via ;
        RECT 1751.780 1325.020 1752.040 1325.280 ;
        RECT 1769.720 1325.020 1769.980 1325.280 ;
        RECT 1751.780 717.440 1752.040 717.700 ;
        RECT 1751.780 716.760 1752.040 717.020 ;
        RECT 1311.100 19.080 1311.360 19.340 ;
        RECT 1751.780 16.360 1752.040 16.620 ;
      LAYER met2 ;
        RECT 1769.710 2203.355 1769.990 2203.725 ;
        RECT 1769.780 1325.310 1769.920 2203.355 ;
        RECT 1751.780 1324.990 1752.040 1325.310 ;
        RECT 1769.720 1324.990 1769.980 1325.310 ;
        RECT 1751.840 717.730 1751.980 1324.990 ;
        RECT 1751.780 717.410 1752.040 717.730 ;
        RECT 1751.780 716.730 1752.040 717.050 ;
        RECT 1311.100 19.050 1311.360 19.370 ;
        RECT 1311.160 2.400 1311.300 19.050 ;
        RECT 1751.840 16.650 1751.980 716.730 ;
        RECT 1751.780 16.330 1752.040 16.650 ;
        RECT 1310.950 -4.800 1311.510 2.400 ;
      LAYER via2 ;
        RECT 1769.710 2203.400 1769.990 2203.680 ;
      LAYER met3 ;
        RECT 1755.835 2203.690 1759.835 2203.695 ;
        RECT 1769.685 2203.690 1770.015 2203.705 ;
        RECT 1755.835 2203.390 1770.015 2203.690 ;
        RECT 1755.835 2203.095 1759.835 2203.390 ;
        RECT 1769.685 2203.375 1770.015 2203.390 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1771.145 1352.265 1771.315 1357.535 ;
      LAYER mcon ;
        RECT 1771.145 1357.365 1771.315 1357.535 ;
      LAYER met1 ;
        RECT 1771.070 1357.520 1771.390 1357.580 ;
        RECT 1770.875 1357.380 1771.390 1357.520 ;
        RECT 1771.070 1357.320 1771.390 1357.380 ;
        RECT 1769.230 1352.420 1769.550 1352.480 ;
        RECT 1771.085 1352.420 1771.375 1352.465 ;
        RECT 1769.230 1352.280 1771.375 1352.420 ;
        RECT 1769.230 1352.220 1769.550 1352.280 ;
        RECT 1771.085 1352.235 1771.375 1352.280 ;
        RECT 1749.450 1319.440 1749.770 1319.500 ;
        RECT 1769.230 1319.440 1769.550 1319.500 ;
        RECT 1749.450 1319.300 1769.550 1319.440 ;
        RECT 1749.450 1319.240 1749.770 1319.300 ;
        RECT 1769.230 1319.240 1769.550 1319.300 ;
        RECT 1329.010 19.620 1329.330 19.680 ;
        RECT 1329.010 19.480 1726.220 19.620 ;
        RECT 1329.010 19.420 1329.330 19.480 ;
        RECT 1726.080 19.280 1726.220 19.480 ;
        RECT 1749.450 19.280 1749.770 19.340 ;
        RECT 1726.080 19.140 1749.770 19.280 ;
        RECT 1749.450 19.080 1749.770 19.140 ;
      LAYER via ;
        RECT 1771.100 1357.320 1771.360 1357.580 ;
        RECT 1769.260 1352.220 1769.520 1352.480 ;
        RECT 1749.480 1319.240 1749.740 1319.500 ;
        RECT 1769.260 1319.240 1769.520 1319.500 ;
        RECT 1329.040 19.420 1329.300 19.680 ;
        RECT 1749.480 19.080 1749.740 19.340 ;
      LAYER met2 ;
        RECT 1771.090 2074.155 1771.370 2074.525 ;
        RECT 1771.160 1357.610 1771.300 2074.155 ;
        RECT 1771.100 1357.290 1771.360 1357.610 ;
        RECT 1769.260 1352.190 1769.520 1352.510 ;
        RECT 1769.320 1319.530 1769.460 1352.190 ;
        RECT 1749.480 1319.210 1749.740 1319.530 ;
        RECT 1769.260 1319.210 1769.520 1319.530 ;
        RECT 1329.040 19.390 1329.300 19.710 ;
        RECT 1329.100 2.400 1329.240 19.390 ;
        RECT 1749.540 19.370 1749.680 1319.210 ;
        RECT 1749.480 19.050 1749.740 19.370 ;
        RECT 1328.890 -4.800 1329.450 2.400 ;
      LAYER via2 ;
        RECT 1771.090 2074.200 1771.370 2074.480 ;
      LAYER met3 ;
        RECT 1755.835 2074.490 1759.835 2074.495 ;
        RECT 1771.065 2074.490 1771.395 2074.505 ;
        RECT 1755.835 2074.190 1771.395 2074.490 ;
        RECT 1755.835 2073.895 1759.835 2074.190 ;
        RECT 1771.065 2074.175 1771.395 2074.190 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 686.850 24.720 687.170 24.780 ;
        RECT 793.570 24.720 793.890 24.780 ;
        RECT 686.850 24.580 793.890 24.720 ;
        RECT 686.850 24.520 687.170 24.580 ;
        RECT 793.570 24.520 793.890 24.580 ;
      LAYER via ;
        RECT 686.880 24.520 687.140 24.780 ;
        RECT 793.600 24.520 793.860 24.780 ;
      LAYER met2 ;
        RECT 799.620 1323.690 799.900 1327.135 ;
        RECT 793.660 1323.550 799.900 1323.690 ;
        RECT 793.660 24.810 793.800 1323.550 ;
        RECT 799.620 1323.135 799.900 1323.550 ;
        RECT 686.880 24.490 687.140 24.810 ;
        RECT 793.600 24.490 793.860 24.810 ;
        RECT 686.940 12.650 687.080 24.490 ;
        RECT 686.480 12.510 687.080 12.650 ;
        RECT 686.480 2.400 686.620 12.510 ;
        RECT 686.270 -4.800 686.830 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 709.850 26.760 710.170 26.820 ;
        RECT 1346.490 26.760 1346.810 26.820 ;
        RECT 709.850 26.620 1346.810 26.760 ;
        RECT 709.850 26.560 710.170 26.620 ;
        RECT 1346.490 26.560 1346.810 26.620 ;
      LAYER via ;
        RECT 709.880 26.560 710.140 26.820 ;
        RECT 1346.520 26.560 1346.780 26.820 ;
      LAYER met2 ;
        RECT 709.870 2215.595 710.150 2215.965 ;
        RECT 709.940 26.850 710.080 2215.595 ;
        RECT 709.880 26.530 710.140 26.850 ;
        RECT 1346.520 26.530 1346.780 26.850 ;
        RECT 1346.580 2.400 1346.720 26.530 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
      LAYER via2 ;
        RECT 709.870 2215.640 710.150 2215.920 ;
      LAYER met3 ;
        RECT 709.845 2215.930 710.175 2215.945 ;
        RECT 715.810 2215.930 719.810 2215.935 ;
        RECT 709.845 2215.630 719.810 2215.930 ;
        RECT 709.845 2215.615 710.175 2215.630 ;
        RECT 715.810 2215.335 719.810 2215.630 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1698.925 2388.245 1699.095 2392.495 ;
      LAYER mcon ;
        RECT 1698.925 2392.325 1699.095 2392.495 ;
      LAYER met1 ;
        RECT 1357.990 2392.480 1358.310 2392.540 ;
        RECT 1698.865 2392.480 1699.155 2392.525 ;
        RECT 1357.990 2392.340 1699.155 2392.480 ;
        RECT 1357.990 2392.280 1358.310 2392.340 ;
        RECT 1698.865 2392.295 1699.155 2392.340 ;
        RECT 1698.865 2388.400 1699.155 2388.445 ;
        RECT 1711.270 2388.400 1711.590 2388.460 ;
        RECT 1698.865 2388.260 1711.590 2388.400 ;
        RECT 1698.865 2388.215 1699.155 2388.260 ;
        RECT 1711.270 2388.200 1711.590 2388.260 ;
        RECT 1711.270 2379.560 1711.590 2379.620 ;
        RECT 1775.670 2379.560 1775.990 2379.620 ;
        RECT 1711.270 2379.420 1775.990 2379.560 ;
        RECT 1711.270 2379.360 1711.590 2379.420 ;
        RECT 1775.670 2379.360 1775.990 2379.420 ;
        RECT 1364.430 32.540 1364.750 32.600 ;
        RECT 1775.670 32.540 1775.990 32.600 ;
        RECT 1364.430 32.400 1775.990 32.540 ;
        RECT 1364.430 32.340 1364.750 32.400 ;
        RECT 1775.670 32.340 1775.990 32.400 ;
      LAYER via ;
        RECT 1358.020 2392.280 1358.280 2392.540 ;
        RECT 1711.300 2388.200 1711.560 2388.460 ;
        RECT 1711.300 2379.360 1711.560 2379.620 ;
        RECT 1775.700 2379.360 1775.960 2379.620 ;
        RECT 1364.460 32.340 1364.720 32.600 ;
        RECT 1775.700 32.340 1775.960 32.600 ;
      LAYER met2 ;
        RECT 1358.020 2392.250 1358.280 2392.570 ;
        RECT 1358.080 2377.880 1358.220 2392.250 ;
        RECT 1711.300 2388.170 1711.560 2388.490 ;
        RECT 1711.360 2379.650 1711.500 2388.170 ;
        RECT 1711.300 2379.330 1711.560 2379.650 ;
        RECT 1775.700 2379.330 1775.960 2379.650 ;
        RECT 1358.060 2373.880 1358.340 2377.880 ;
        RECT 1775.760 32.630 1775.900 2379.330 ;
        RECT 1364.460 32.310 1364.720 32.630 ;
        RECT 1775.700 32.310 1775.960 32.630 ;
        RECT 1364.520 2.400 1364.660 32.310 ;
        RECT 1364.310 -4.800 1364.870 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 706.705 1337.985 706.875 1356.175 ;
        RECT 743.045 1309.085 743.215 1322.855 ;
        RECT 1380.145 338.385 1380.315 386.155 ;
        RECT 1380.145 241.825 1380.315 289.595 ;
        RECT 1380.145 145.265 1380.315 193.035 ;
        RECT 1380.145 48.705 1380.315 96.475 ;
        RECT 1382.445 2.805 1382.615 48.195 ;
      LAYER mcon ;
        RECT 706.705 1356.005 706.875 1356.175 ;
        RECT 743.045 1322.685 743.215 1322.855 ;
        RECT 1380.145 385.985 1380.315 386.155 ;
        RECT 1380.145 289.425 1380.315 289.595 ;
        RECT 1380.145 192.865 1380.315 193.035 ;
        RECT 1380.145 96.305 1380.315 96.475 ;
        RECT 1382.445 48.025 1382.615 48.195 ;
      LAYER met1 ;
        RECT 706.630 1356.160 706.950 1356.220 ;
        RECT 706.435 1356.020 706.950 1356.160 ;
        RECT 706.630 1355.960 706.950 1356.020 ;
        RECT 706.630 1338.140 706.950 1338.200 ;
        RECT 706.435 1338.000 706.950 1338.140 ;
        RECT 706.630 1337.940 706.950 1338.000 ;
        RECT 706.630 1322.840 706.950 1322.900 ;
        RECT 742.985 1322.840 743.275 1322.885 ;
        RECT 706.630 1322.700 743.275 1322.840 ;
        RECT 706.630 1322.640 706.950 1322.700 ;
        RECT 742.985 1322.655 743.275 1322.700 ;
        RECT 742.985 1309.240 743.275 1309.285 ;
        RECT 1380.070 1309.240 1380.390 1309.300 ;
        RECT 742.985 1309.100 1380.390 1309.240 ;
        RECT 742.985 1309.055 743.275 1309.100 ;
        RECT 1380.070 1309.040 1380.390 1309.100 ;
        RECT 1380.070 1256.680 1380.390 1256.940 ;
        RECT 1380.160 1256.260 1380.300 1256.680 ;
        RECT 1380.070 1256.000 1380.390 1256.260 ;
        RECT 1380.070 1207.580 1380.390 1207.640 ;
        RECT 1380.990 1207.580 1381.310 1207.640 ;
        RECT 1380.070 1207.440 1381.310 1207.580 ;
        RECT 1380.070 1207.380 1380.390 1207.440 ;
        RECT 1380.990 1207.380 1381.310 1207.440 ;
        RECT 1380.070 1111.020 1380.390 1111.080 ;
        RECT 1380.990 1111.020 1381.310 1111.080 ;
        RECT 1380.070 1110.880 1381.310 1111.020 ;
        RECT 1380.070 1110.820 1380.390 1110.880 ;
        RECT 1380.990 1110.820 1381.310 1110.880 ;
        RECT 1380.070 1014.460 1380.390 1014.520 ;
        RECT 1380.990 1014.460 1381.310 1014.520 ;
        RECT 1380.070 1014.320 1381.310 1014.460 ;
        RECT 1380.070 1014.260 1380.390 1014.320 ;
        RECT 1380.990 1014.260 1381.310 1014.320 ;
        RECT 1380.070 917.900 1380.390 917.960 ;
        RECT 1380.990 917.900 1381.310 917.960 ;
        RECT 1380.070 917.760 1381.310 917.900 ;
        RECT 1380.070 917.700 1380.390 917.760 ;
        RECT 1380.990 917.700 1381.310 917.760 ;
        RECT 1380.070 869.620 1380.390 869.680 ;
        RECT 1380.990 869.620 1381.310 869.680 ;
        RECT 1380.070 869.480 1381.310 869.620 ;
        RECT 1380.070 869.420 1380.390 869.480 ;
        RECT 1380.990 869.420 1381.310 869.480 ;
        RECT 1380.070 772.720 1380.390 772.780 ;
        RECT 1380.990 772.720 1381.310 772.780 ;
        RECT 1380.070 772.580 1381.310 772.720 ;
        RECT 1380.070 772.520 1380.390 772.580 ;
        RECT 1380.990 772.520 1381.310 772.580 ;
        RECT 1380.070 676.160 1380.390 676.220 ;
        RECT 1380.990 676.160 1381.310 676.220 ;
        RECT 1380.070 676.020 1381.310 676.160 ;
        RECT 1380.070 675.960 1380.390 676.020 ;
        RECT 1380.990 675.960 1381.310 676.020 ;
        RECT 1380.070 579.600 1380.390 579.660 ;
        RECT 1380.990 579.600 1381.310 579.660 ;
        RECT 1380.070 579.460 1381.310 579.600 ;
        RECT 1380.070 579.400 1380.390 579.460 ;
        RECT 1380.990 579.400 1381.310 579.460 ;
        RECT 1380.070 483.040 1380.390 483.100 ;
        RECT 1380.990 483.040 1381.310 483.100 ;
        RECT 1380.070 482.900 1381.310 483.040 ;
        RECT 1380.070 482.840 1380.390 482.900 ;
        RECT 1380.990 482.840 1381.310 482.900 ;
        RECT 1380.070 386.140 1380.390 386.200 ;
        RECT 1379.875 386.000 1380.390 386.140 ;
        RECT 1380.070 385.940 1380.390 386.000 ;
        RECT 1380.070 338.540 1380.390 338.600 ;
        RECT 1379.875 338.400 1380.390 338.540 ;
        RECT 1380.070 338.340 1380.390 338.400 ;
        RECT 1380.070 337.860 1380.390 337.920 ;
        RECT 1380.530 337.860 1380.850 337.920 ;
        RECT 1380.070 337.720 1380.850 337.860 ;
        RECT 1380.070 337.660 1380.390 337.720 ;
        RECT 1380.530 337.660 1380.850 337.720 ;
        RECT 1380.070 289.580 1380.390 289.640 ;
        RECT 1379.875 289.440 1380.390 289.580 ;
        RECT 1380.070 289.380 1380.390 289.440 ;
        RECT 1380.070 241.980 1380.390 242.040 ;
        RECT 1379.875 241.840 1380.390 241.980 ;
        RECT 1380.070 241.780 1380.390 241.840 ;
        RECT 1380.070 241.300 1380.390 241.360 ;
        RECT 1380.530 241.300 1380.850 241.360 ;
        RECT 1380.070 241.160 1380.850 241.300 ;
        RECT 1380.070 241.100 1380.390 241.160 ;
        RECT 1380.530 241.100 1380.850 241.160 ;
        RECT 1380.070 193.020 1380.390 193.080 ;
        RECT 1379.875 192.880 1380.390 193.020 ;
        RECT 1380.070 192.820 1380.390 192.880 ;
        RECT 1380.070 145.420 1380.390 145.480 ;
        RECT 1379.875 145.280 1380.390 145.420 ;
        RECT 1380.070 145.220 1380.390 145.280 ;
        RECT 1380.070 144.740 1380.390 144.800 ;
        RECT 1380.530 144.740 1380.850 144.800 ;
        RECT 1380.070 144.600 1380.850 144.740 ;
        RECT 1380.070 144.540 1380.390 144.600 ;
        RECT 1380.530 144.540 1380.850 144.600 ;
        RECT 1380.070 96.460 1380.390 96.520 ;
        RECT 1379.875 96.320 1380.390 96.460 ;
        RECT 1380.070 96.260 1380.390 96.320 ;
        RECT 1380.070 48.860 1380.390 48.920 ;
        RECT 1379.875 48.720 1380.390 48.860 ;
        RECT 1380.070 48.660 1380.390 48.720 ;
        RECT 1380.070 48.180 1380.390 48.240 ;
        RECT 1382.385 48.180 1382.675 48.225 ;
        RECT 1380.070 48.040 1382.675 48.180 ;
        RECT 1380.070 47.980 1380.390 48.040 ;
        RECT 1382.385 47.995 1382.675 48.040 ;
        RECT 1382.370 2.960 1382.690 3.020 ;
        RECT 1382.175 2.820 1382.690 2.960 ;
        RECT 1382.370 2.760 1382.690 2.820 ;
      LAYER via ;
        RECT 706.660 1355.960 706.920 1356.220 ;
        RECT 706.660 1337.940 706.920 1338.200 ;
        RECT 706.660 1322.640 706.920 1322.900 ;
        RECT 1380.100 1309.040 1380.360 1309.300 ;
        RECT 1380.100 1256.680 1380.360 1256.940 ;
        RECT 1380.100 1256.000 1380.360 1256.260 ;
        RECT 1380.100 1207.380 1380.360 1207.640 ;
        RECT 1381.020 1207.380 1381.280 1207.640 ;
        RECT 1380.100 1110.820 1380.360 1111.080 ;
        RECT 1381.020 1110.820 1381.280 1111.080 ;
        RECT 1380.100 1014.260 1380.360 1014.520 ;
        RECT 1381.020 1014.260 1381.280 1014.520 ;
        RECT 1380.100 917.700 1380.360 917.960 ;
        RECT 1381.020 917.700 1381.280 917.960 ;
        RECT 1380.100 869.420 1380.360 869.680 ;
        RECT 1381.020 869.420 1381.280 869.680 ;
        RECT 1380.100 772.520 1380.360 772.780 ;
        RECT 1381.020 772.520 1381.280 772.780 ;
        RECT 1380.100 675.960 1380.360 676.220 ;
        RECT 1381.020 675.960 1381.280 676.220 ;
        RECT 1380.100 579.400 1380.360 579.660 ;
        RECT 1381.020 579.400 1381.280 579.660 ;
        RECT 1380.100 482.840 1380.360 483.100 ;
        RECT 1381.020 482.840 1381.280 483.100 ;
        RECT 1380.100 385.940 1380.360 386.200 ;
        RECT 1380.100 338.340 1380.360 338.600 ;
        RECT 1380.100 337.660 1380.360 337.920 ;
        RECT 1380.560 337.660 1380.820 337.920 ;
        RECT 1380.100 289.380 1380.360 289.640 ;
        RECT 1380.100 241.780 1380.360 242.040 ;
        RECT 1380.100 241.100 1380.360 241.360 ;
        RECT 1380.560 241.100 1380.820 241.360 ;
        RECT 1380.100 192.820 1380.360 193.080 ;
        RECT 1380.100 145.220 1380.360 145.480 ;
        RECT 1380.100 144.540 1380.360 144.800 ;
        RECT 1380.560 144.540 1380.820 144.800 ;
        RECT 1380.100 96.260 1380.360 96.520 ;
        RECT 1380.100 48.660 1380.360 48.920 ;
        RECT 1380.100 47.980 1380.360 48.240 ;
        RECT 1382.400 2.760 1382.660 3.020 ;
      LAYER met2 ;
        RECT 706.650 1377.835 706.930 1378.205 ;
        RECT 706.720 1356.250 706.860 1377.835 ;
        RECT 706.660 1355.930 706.920 1356.250 ;
        RECT 706.660 1337.910 706.920 1338.230 ;
        RECT 706.720 1322.930 706.860 1337.910 ;
        RECT 706.660 1322.610 706.920 1322.930 ;
        RECT 1380.100 1309.010 1380.360 1309.330 ;
        RECT 1380.160 1256.970 1380.300 1309.010 ;
        RECT 1380.100 1256.650 1380.360 1256.970 ;
        RECT 1380.100 1255.970 1380.360 1256.290 ;
        RECT 1380.160 1255.805 1380.300 1255.970 ;
        RECT 1380.090 1255.435 1380.370 1255.805 ;
        RECT 1381.010 1255.435 1381.290 1255.805 ;
        RECT 1381.080 1207.670 1381.220 1255.435 ;
        RECT 1380.100 1207.350 1380.360 1207.670 ;
        RECT 1381.020 1207.350 1381.280 1207.670 ;
        RECT 1380.160 1159.245 1380.300 1207.350 ;
        RECT 1380.090 1158.875 1380.370 1159.245 ;
        RECT 1381.010 1158.875 1381.290 1159.245 ;
        RECT 1381.080 1111.110 1381.220 1158.875 ;
        RECT 1380.100 1110.790 1380.360 1111.110 ;
        RECT 1381.020 1110.790 1381.280 1111.110 ;
        RECT 1380.160 1062.685 1380.300 1110.790 ;
        RECT 1380.090 1062.315 1380.370 1062.685 ;
        RECT 1381.010 1062.315 1381.290 1062.685 ;
        RECT 1381.080 1014.550 1381.220 1062.315 ;
        RECT 1380.100 1014.230 1380.360 1014.550 ;
        RECT 1381.020 1014.230 1381.280 1014.550 ;
        RECT 1380.160 966.125 1380.300 1014.230 ;
        RECT 1380.090 965.755 1380.370 966.125 ;
        RECT 1381.010 965.755 1381.290 966.125 ;
        RECT 1381.080 917.990 1381.220 965.755 ;
        RECT 1380.100 917.845 1380.360 917.990 ;
        RECT 1381.020 917.845 1381.280 917.990 ;
        RECT 1380.090 917.475 1380.370 917.845 ;
        RECT 1381.010 917.475 1381.290 917.845 ;
        RECT 1381.080 869.710 1381.220 917.475 ;
        RECT 1380.100 869.565 1380.360 869.710 ;
        RECT 1381.020 869.565 1381.280 869.710 ;
        RECT 1380.090 869.195 1380.370 869.565 ;
        RECT 1381.010 869.195 1381.290 869.565 ;
        RECT 1381.080 821.285 1381.220 869.195 ;
        RECT 1380.090 820.915 1380.370 821.285 ;
        RECT 1381.010 820.915 1381.290 821.285 ;
        RECT 1380.160 772.810 1380.300 820.915 ;
        RECT 1380.100 772.490 1380.360 772.810 ;
        RECT 1381.020 772.490 1381.280 772.810 ;
        RECT 1381.080 724.725 1381.220 772.490 ;
        RECT 1380.090 724.355 1380.370 724.725 ;
        RECT 1381.010 724.355 1381.290 724.725 ;
        RECT 1380.160 676.250 1380.300 724.355 ;
        RECT 1380.100 675.930 1380.360 676.250 ;
        RECT 1381.020 675.930 1381.280 676.250 ;
        RECT 1381.080 628.165 1381.220 675.930 ;
        RECT 1380.090 627.795 1380.370 628.165 ;
        RECT 1381.010 627.795 1381.290 628.165 ;
        RECT 1380.160 580.565 1380.300 627.795 ;
        RECT 1380.090 580.195 1380.370 580.565 ;
        RECT 1380.090 579.515 1380.370 579.885 ;
        RECT 1380.100 579.370 1380.360 579.515 ;
        RECT 1381.020 579.370 1381.280 579.690 ;
        RECT 1381.080 531.605 1381.220 579.370 ;
        RECT 1380.090 531.235 1380.370 531.605 ;
        RECT 1381.010 531.235 1381.290 531.605 ;
        RECT 1380.160 484.005 1380.300 531.235 ;
        RECT 1380.090 483.635 1380.370 484.005 ;
        RECT 1380.090 482.955 1380.370 483.325 ;
        RECT 1380.100 482.810 1380.360 482.955 ;
        RECT 1381.020 482.810 1381.280 483.130 ;
        RECT 1381.080 435.045 1381.220 482.810 ;
        RECT 1380.090 434.675 1380.370 435.045 ;
        RECT 1381.010 434.675 1381.290 435.045 ;
        RECT 1380.160 386.230 1380.300 434.675 ;
        RECT 1380.100 385.910 1380.360 386.230 ;
        RECT 1380.100 338.310 1380.360 338.630 ;
        RECT 1380.160 337.950 1380.300 338.310 ;
        RECT 1380.100 337.630 1380.360 337.950 ;
        RECT 1380.560 337.630 1380.820 337.950 ;
        RECT 1380.620 290.090 1380.760 337.630 ;
        RECT 1380.160 289.950 1380.760 290.090 ;
        RECT 1380.160 289.670 1380.300 289.950 ;
        RECT 1380.100 289.350 1380.360 289.670 ;
        RECT 1380.100 241.750 1380.360 242.070 ;
        RECT 1380.160 241.390 1380.300 241.750 ;
        RECT 1380.100 241.070 1380.360 241.390 ;
        RECT 1380.560 241.070 1380.820 241.390 ;
        RECT 1380.620 193.530 1380.760 241.070 ;
        RECT 1380.160 193.390 1380.760 193.530 ;
        RECT 1380.160 193.110 1380.300 193.390 ;
        RECT 1380.100 192.790 1380.360 193.110 ;
        RECT 1380.100 145.190 1380.360 145.510 ;
        RECT 1380.160 144.830 1380.300 145.190 ;
        RECT 1380.100 144.510 1380.360 144.830 ;
        RECT 1380.560 144.510 1380.820 144.830 ;
        RECT 1380.620 96.970 1380.760 144.510 ;
        RECT 1380.160 96.830 1380.760 96.970 ;
        RECT 1380.160 96.550 1380.300 96.830 ;
        RECT 1380.100 96.230 1380.360 96.550 ;
        RECT 1380.100 48.630 1380.360 48.950 ;
        RECT 1380.160 48.270 1380.300 48.630 ;
        RECT 1380.100 47.950 1380.360 48.270 ;
        RECT 1382.400 2.730 1382.660 3.050 ;
        RECT 1382.460 2.400 1382.600 2.730 ;
        RECT 1382.250 -4.800 1382.810 2.400 ;
      LAYER via2 ;
        RECT 706.650 1377.880 706.930 1378.160 ;
        RECT 1380.090 1255.480 1380.370 1255.760 ;
        RECT 1381.010 1255.480 1381.290 1255.760 ;
        RECT 1380.090 1158.920 1380.370 1159.200 ;
        RECT 1381.010 1158.920 1381.290 1159.200 ;
        RECT 1380.090 1062.360 1380.370 1062.640 ;
        RECT 1381.010 1062.360 1381.290 1062.640 ;
        RECT 1380.090 965.800 1380.370 966.080 ;
        RECT 1381.010 965.800 1381.290 966.080 ;
        RECT 1380.090 917.520 1380.370 917.800 ;
        RECT 1381.010 917.520 1381.290 917.800 ;
        RECT 1380.090 869.240 1380.370 869.520 ;
        RECT 1381.010 869.240 1381.290 869.520 ;
        RECT 1380.090 820.960 1380.370 821.240 ;
        RECT 1381.010 820.960 1381.290 821.240 ;
        RECT 1380.090 724.400 1380.370 724.680 ;
        RECT 1381.010 724.400 1381.290 724.680 ;
        RECT 1380.090 627.840 1380.370 628.120 ;
        RECT 1381.010 627.840 1381.290 628.120 ;
        RECT 1380.090 580.240 1380.370 580.520 ;
        RECT 1380.090 579.560 1380.370 579.840 ;
        RECT 1380.090 531.280 1380.370 531.560 ;
        RECT 1381.010 531.280 1381.290 531.560 ;
        RECT 1380.090 483.680 1380.370 483.960 ;
        RECT 1380.090 483.000 1380.370 483.280 ;
        RECT 1380.090 434.720 1380.370 435.000 ;
        RECT 1381.010 434.720 1381.290 435.000 ;
      LAYER met3 ;
        RECT 706.625 1378.170 706.955 1378.185 ;
        RECT 715.810 1378.170 719.810 1378.175 ;
        RECT 706.625 1377.870 719.810 1378.170 ;
        RECT 706.625 1377.855 706.955 1377.870 ;
        RECT 715.810 1377.575 719.810 1377.870 ;
        RECT 1380.065 1255.770 1380.395 1255.785 ;
        RECT 1380.985 1255.770 1381.315 1255.785 ;
        RECT 1380.065 1255.470 1381.315 1255.770 ;
        RECT 1380.065 1255.455 1380.395 1255.470 ;
        RECT 1380.985 1255.455 1381.315 1255.470 ;
        RECT 1380.065 1159.210 1380.395 1159.225 ;
        RECT 1380.985 1159.210 1381.315 1159.225 ;
        RECT 1380.065 1158.910 1381.315 1159.210 ;
        RECT 1380.065 1158.895 1380.395 1158.910 ;
        RECT 1380.985 1158.895 1381.315 1158.910 ;
        RECT 1380.065 1062.650 1380.395 1062.665 ;
        RECT 1380.985 1062.650 1381.315 1062.665 ;
        RECT 1380.065 1062.350 1381.315 1062.650 ;
        RECT 1380.065 1062.335 1380.395 1062.350 ;
        RECT 1380.985 1062.335 1381.315 1062.350 ;
        RECT 1380.065 966.090 1380.395 966.105 ;
        RECT 1380.985 966.090 1381.315 966.105 ;
        RECT 1380.065 965.790 1381.315 966.090 ;
        RECT 1380.065 965.775 1380.395 965.790 ;
        RECT 1380.985 965.775 1381.315 965.790 ;
        RECT 1380.065 917.810 1380.395 917.825 ;
        RECT 1380.985 917.810 1381.315 917.825 ;
        RECT 1380.065 917.510 1381.315 917.810 ;
        RECT 1380.065 917.495 1380.395 917.510 ;
        RECT 1380.985 917.495 1381.315 917.510 ;
        RECT 1380.065 869.530 1380.395 869.545 ;
        RECT 1380.985 869.530 1381.315 869.545 ;
        RECT 1380.065 869.230 1381.315 869.530 ;
        RECT 1380.065 869.215 1380.395 869.230 ;
        RECT 1380.985 869.215 1381.315 869.230 ;
        RECT 1380.065 821.250 1380.395 821.265 ;
        RECT 1380.985 821.250 1381.315 821.265 ;
        RECT 1380.065 820.950 1381.315 821.250 ;
        RECT 1380.065 820.935 1380.395 820.950 ;
        RECT 1380.985 820.935 1381.315 820.950 ;
        RECT 1380.065 724.690 1380.395 724.705 ;
        RECT 1380.985 724.690 1381.315 724.705 ;
        RECT 1380.065 724.390 1381.315 724.690 ;
        RECT 1380.065 724.375 1380.395 724.390 ;
        RECT 1380.985 724.375 1381.315 724.390 ;
        RECT 1380.065 628.130 1380.395 628.145 ;
        RECT 1380.985 628.130 1381.315 628.145 ;
        RECT 1380.065 627.830 1381.315 628.130 ;
        RECT 1380.065 627.815 1380.395 627.830 ;
        RECT 1380.985 627.815 1381.315 627.830 ;
        RECT 1380.065 580.530 1380.395 580.545 ;
        RECT 1379.390 580.230 1380.395 580.530 ;
        RECT 1379.390 579.850 1379.690 580.230 ;
        RECT 1380.065 580.215 1380.395 580.230 ;
        RECT 1380.065 579.850 1380.395 579.865 ;
        RECT 1379.390 579.550 1380.395 579.850 ;
        RECT 1380.065 579.535 1380.395 579.550 ;
        RECT 1380.065 531.570 1380.395 531.585 ;
        RECT 1380.985 531.570 1381.315 531.585 ;
        RECT 1380.065 531.270 1381.315 531.570 ;
        RECT 1380.065 531.255 1380.395 531.270 ;
        RECT 1380.985 531.255 1381.315 531.270 ;
        RECT 1380.065 483.970 1380.395 483.985 ;
        RECT 1379.390 483.670 1380.395 483.970 ;
        RECT 1379.390 483.290 1379.690 483.670 ;
        RECT 1380.065 483.655 1380.395 483.670 ;
        RECT 1380.065 483.290 1380.395 483.305 ;
        RECT 1379.390 482.990 1380.395 483.290 ;
        RECT 1380.065 482.975 1380.395 482.990 ;
        RECT 1380.065 435.010 1380.395 435.025 ;
        RECT 1380.985 435.010 1381.315 435.025 ;
        RECT 1380.065 434.710 1381.315 435.010 ;
        RECT 1380.065 434.695 1380.395 434.710 ;
        RECT 1380.985 434.695 1381.315 434.710 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 703.945 1335.945 704.115 1393.575 ;
      LAYER mcon ;
        RECT 703.945 1393.405 704.115 1393.575 ;
      LAYER met1 ;
        RECT 703.870 1393.560 704.190 1393.620 ;
        RECT 703.675 1393.420 704.190 1393.560 ;
        RECT 703.870 1393.360 704.190 1393.420 ;
        RECT 703.870 1336.100 704.190 1336.160 ;
        RECT 703.870 1335.960 704.385 1336.100 ;
        RECT 703.870 1335.900 704.190 1335.960 ;
        RECT 703.870 26.080 704.190 26.140 ;
        RECT 1400.310 26.080 1400.630 26.140 ;
        RECT 703.870 25.940 1400.630 26.080 ;
        RECT 703.870 25.880 704.190 25.940 ;
        RECT 1400.310 25.880 1400.630 25.940 ;
      LAYER via ;
        RECT 703.900 1393.360 704.160 1393.620 ;
        RECT 703.900 1335.900 704.160 1336.160 ;
        RECT 703.900 25.880 704.160 26.140 ;
        RECT 1400.340 25.880 1400.600 26.140 ;
      LAYER met2 ;
        RECT 703.890 2318.955 704.170 2319.325 ;
        RECT 703.960 1393.650 704.100 2318.955 ;
        RECT 703.900 1393.330 704.160 1393.650 ;
        RECT 703.900 1335.870 704.160 1336.190 ;
        RECT 703.960 26.170 704.100 1335.870 ;
        RECT 703.900 25.850 704.160 26.170 ;
        RECT 1400.340 25.850 1400.600 26.170 ;
        RECT 1400.400 2.400 1400.540 25.850 ;
        RECT 1400.190 -4.800 1400.750 2.400 ;
      LAYER via2 ;
        RECT 703.890 2319.000 704.170 2319.280 ;
      LAYER met3 ;
        RECT 703.865 2319.290 704.195 2319.305 ;
        RECT 715.810 2319.290 719.810 2319.295 ;
        RECT 703.865 2318.990 719.810 2319.290 ;
        RECT 703.865 2318.975 704.195 2318.990 ;
        RECT 715.810 2318.695 719.810 2318.990 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1726.525 19.465 1726.695 20.315 ;
      LAYER mcon ;
        RECT 1726.525 20.145 1726.695 20.315 ;
      LAYER met1 ;
        RECT 1771.070 1356.840 1771.390 1356.900 ;
        RECT 1772.450 1356.840 1772.770 1356.900 ;
        RECT 1771.070 1356.700 1772.770 1356.840 ;
        RECT 1771.070 1356.640 1771.390 1356.700 ;
        RECT 1772.450 1356.640 1772.770 1356.700 ;
        RECT 1748.990 1321.820 1749.310 1321.880 ;
        RECT 1771.070 1321.820 1771.390 1321.880 ;
        RECT 1748.990 1321.680 1771.390 1321.820 ;
        RECT 1748.990 1321.620 1749.310 1321.680 ;
        RECT 1771.070 1321.620 1771.390 1321.680 ;
        RECT 1418.250 20.300 1418.570 20.360 ;
        RECT 1726.465 20.300 1726.755 20.345 ;
        RECT 1418.250 20.160 1726.755 20.300 ;
        RECT 1418.250 20.100 1418.570 20.160 ;
        RECT 1726.465 20.115 1726.755 20.160 ;
        RECT 1726.465 19.620 1726.755 19.665 ;
        RECT 1748.990 19.620 1749.310 19.680 ;
        RECT 1726.465 19.480 1749.310 19.620 ;
        RECT 1726.465 19.435 1726.755 19.480 ;
        RECT 1748.990 19.420 1749.310 19.480 ;
      LAYER via ;
        RECT 1771.100 1356.640 1771.360 1356.900 ;
        RECT 1772.480 1356.640 1772.740 1356.900 ;
        RECT 1749.020 1321.620 1749.280 1321.880 ;
        RECT 1771.100 1321.620 1771.360 1321.880 ;
        RECT 1418.280 20.100 1418.540 20.360 ;
        RECT 1749.020 19.420 1749.280 19.680 ;
      LAYER met2 ;
        RECT 1772.470 1493.435 1772.750 1493.805 ;
        RECT 1772.540 1356.930 1772.680 1493.435 ;
        RECT 1771.100 1356.610 1771.360 1356.930 ;
        RECT 1772.480 1356.610 1772.740 1356.930 ;
        RECT 1771.160 1321.910 1771.300 1356.610 ;
        RECT 1749.020 1321.590 1749.280 1321.910 ;
        RECT 1771.100 1321.590 1771.360 1321.910 ;
        RECT 1418.280 20.070 1418.540 20.390 ;
        RECT 1418.340 2.400 1418.480 20.070 ;
        RECT 1749.080 19.710 1749.220 1321.590 ;
        RECT 1749.020 19.390 1749.280 19.710 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
      LAYER via2 ;
        RECT 1772.470 1493.480 1772.750 1493.760 ;
      LAYER met3 ;
        RECT 1755.835 1493.770 1759.835 1493.775 ;
        RECT 1772.445 1493.770 1772.775 1493.785 ;
        RECT 1755.835 1493.470 1772.775 1493.770 ;
        RECT 1755.835 1493.175 1759.835 1493.470 ;
        RECT 1772.445 1493.455 1772.775 1493.470 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1435.730 19.960 1436.050 20.020 ;
        RECT 1775.210 19.960 1775.530 20.020 ;
        RECT 1435.730 19.820 1775.530 19.960 ;
        RECT 1435.730 19.760 1436.050 19.820 ;
        RECT 1775.210 19.760 1775.530 19.820 ;
      LAYER via ;
        RECT 1435.760 19.760 1436.020 20.020 ;
        RECT 1775.240 19.760 1775.500 20.020 ;
      LAYER met2 ;
        RECT 1369.050 2380.155 1369.330 2380.525 ;
        RECT 1369.120 2377.880 1369.260 2380.155 ;
        RECT 1369.100 2373.880 1369.380 2377.880 ;
        RECT 1775.230 2370.635 1775.510 2371.005 ;
        RECT 1775.300 20.050 1775.440 2370.635 ;
        RECT 1435.760 19.730 1436.020 20.050 ;
        RECT 1775.240 19.730 1775.500 20.050 ;
        RECT 1435.820 2.400 1435.960 19.730 ;
        RECT 1435.610 -4.800 1436.170 2.400 ;
      LAYER via2 ;
        RECT 1369.050 2380.200 1369.330 2380.480 ;
        RECT 1775.230 2370.680 1775.510 2370.960 ;
      LAYER met3 ;
        RECT 1369.025 2380.500 1369.355 2380.505 ;
        RECT 1369.025 2380.490 1369.610 2380.500 ;
        RECT 1369.025 2380.190 1369.810 2380.490 ;
        RECT 1369.025 2380.180 1369.610 2380.190 ;
        RECT 1369.025 2380.175 1369.355 2380.180 ;
        RECT 1369.230 2370.970 1369.610 2370.980 ;
        RECT 1775.205 2370.970 1775.535 2370.985 ;
        RECT 1369.230 2370.670 1775.535 2370.970 ;
        RECT 1369.230 2370.660 1369.610 2370.670 ;
        RECT 1775.205 2370.655 1775.535 2370.670 ;
      LAYER via3 ;
        RECT 1369.260 2380.180 1369.580 2380.500 ;
        RECT 1369.260 2370.660 1369.580 2370.980 ;
      LAYER met4 ;
        RECT 1369.255 2380.175 1369.585 2380.505 ;
        RECT 1369.270 2370.985 1369.570 2380.175 ;
        RECT 1369.255 2370.655 1369.585 2370.985 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 703.025 1361.105 703.195 1393.575 ;
      LAYER mcon ;
        RECT 703.025 1393.405 703.195 1393.575 ;
      LAYER met1 ;
        RECT 702.950 2375.140 703.270 2375.200 ;
        RECT 736.990 2375.140 737.310 2375.200 ;
        RECT 702.950 2375.000 737.310 2375.140 ;
        RECT 702.950 2374.940 703.270 2375.000 ;
        RECT 736.990 2374.940 737.310 2375.000 ;
        RECT 702.950 1393.560 703.270 1393.620 ;
        RECT 702.755 1393.420 703.270 1393.560 ;
        RECT 702.950 1393.360 703.270 1393.420 ;
        RECT 702.950 1361.260 703.270 1361.320 ;
        RECT 702.755 1361.120 703.270 1361.260 ;
        RECT 702.950 1361.060 703.270 1361.120 ;
      LAYER via ;
        RECT 702.980 2374.940 703.240 2375.200 ;
        RECT 737.020 2374.940 737.280 2375.200 ;
        RECT 702.980 1393.360 703.240 1393.620 ;
        RECT 702.980 1361.060 703.240 1361.320 ;
      LAYER met2 ;
        RECT 702.980 2374.910 703.240 2375.230 ;
        RECT 737.020 2374.970 737.280 2375.230 ;
        RECT 738.900 2374.970 739.180 2377.880 ;
        RECT 737.020 2374.910 739.180 2374.970 ;
        RECT 703.040 1393.650 703.180 2374.910 ;
        RECT 737.080 2374.830 739.180 2374.910 ;
        RECT 738.900 2373.880 739.180 2374.830 ;
        RECT 702.980 1393.330 703.240 1393.650 ;
        RECT 702.980 1361.030 703.240 1361.350 ;
        RECT 703.040 16.165 703.180 1361.030 ;
        RECT 702.970 15.795 703.250 16.165 ;
        RECT 1453.690 15.795 1453.970 16.165 ;
        RECT 1453.760 2.400 1453.900 15.795 ;
        RECT 1453.550 -4.800 1454.110 2.400 ;
      LAYER via2 ;
        RECT 702.970 15.840 703.250 16.120 ;
        RECT 1453.690 15.840 1453.970 16.120 ;
      LAYER met3 ;
        RECT 702.945 16.130 703.275 16.145 ;
        RECT 1453.665 16.130 1453.995 16.145 ;
        RECT 702.945 15.830 1453.995 16.130 ;
        RECT 702.945 15.815 703.275 15.830 ;
        RECT 1453.665 15.815 1453.995 15.830 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1035.990 1311.280 1036.310 1311.340 ;
        RECT 1041.510 1311.280 1041.830 1311.340 ;
        RECT 1035.990 1311.140 1041.830 1311.280 ;
        RECT 1035.990 1311.080 1036.310 1311.140 ;
        RECT 1041.510 1311.080 1041.830 1311.140 ;
        RECT 1041.510 27.100 1041.830 27.160 ;
        RECT 1471.610 27.100 1471.930 27.160 ;
        RECT 1041.510 26.960 1471.930 27.100 ;
        RECT 1041.510 26.900 1041.830 26.960 ;
        RECT 1471.610 26.900 1471.930 26.960 ;
      LAYER via ;
        RECT 1036.020 1311.080 1036.280 1311.340 ;
        RECT 1041.540 1311.080 1041.800 1311.340 ;
        RECT 1041.540 26.900 1041.800 27.160 ;
        RECT 1471.640 26.900 1471.900 27.160 ;
      LAYER met2 ;
        RECT 1036.060 1323.135 1036.340 1327.135 ;
        RECT 1036.080 1311.370 1036.220 1323.135 ;
        RECT 1036.020 1311.050 1036.280 1311.370 ;
        RECT 1041.540 1311.050 1041.800 1311.370 ;
        RECT 1041.600 27.190 1041.740 1311.050 ;
        RECT 1041.540 26.870 1041.800 27.190 ;
        RECT 1471.640 26.870 1471.900 27.190 ;
        RECT 1471.700 2.400 1471.840 26.870 ;
        RECT 1471.490 -4.800 1472.050 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1490.010 26.080 1490.330 26.140 ;
        RECT 1531.870 26.080 1532.190 26.140 ;
        RECT 1490.010 25.940 1532.190 26.080 ;
        RECT 1490.010 25.880 1490.330 25.940 ;
        RECT 1531.870 25.880 1532.190 25.940 ;
      LAYER via ;
        RECT 1490.040 25.880 1490.300 26.140 ;
        RECT 1531.900 25.880 1532.160 26.140 ;
      LAYER met2 ;
        RECT 1533.780 1323.690 1534.060 1327.135 ;
        RECT 1531.960 1323.550 1534.060 1323.690 ;
        RECT 1531.960 26.170 1532.100 1323.550 ;
        RECT 1533.780 1323.135 1534.060 1323.550 ;
        RECT 1490.040 25.850 1490.300 26.170 ;
        RECT 1531.900 25.850 1532.160 26.170 ;
        RECT 1490.100 3.130 1490.240 25.850 ;
        RECT 1489.640 2.990 1490.240 3.130 ;
        RECT 1489.640 2.400 1489.780 2.990 ;
        RECT 1489.430 -4.800 1489.990 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1535.165 18.785 1535.335 20.655 ;
        RECT 1583.465 18.785 1583.635 20.655 ;
        RECT 1635.445 18.785 1635.615 20.655 ;
        RECT 1704.445 18.785 1704.615 20.655 ;
        RECT 1724.685 20.485 1727.155 20.655 ;
        RECT 1724.685 18.785 1724.855 20.485 ;
        RECT 1726.985 20.145 1727.155 20.485 ;
        RECT 1738.945 20.145 1739.115 21.675 ;
      LAYER mcon ;
        RECT 1738.945 21.505 1739.115 21.675 ;
        RECT 1535.165 20.485 1535.335 20.655 ;
        RECT 1583.465 20.485 1583.635 20.655 ;
        RECT 1635.445 20.485 1635.615 20.655 ;
        RECT 1704.445 20.485 1704.615 20.655 ;
      LAYER met1 ;
        RECT 1451.370 2378.200 1451.690 2378.260 ;
        RECT 1451.370 2378.060 1753.820 2378.200 ;
        RECT 1451.370 2378.000 1451.690 2378.060 ;
        RECT 1753.680 2377.860 1753.820 2378.060 ;
        RECT 1781.190 2377.860 1781.510 2377.920 ;
        RECT 1753.680 2377.720 1781.510 2377.860 ;
        RECT 1781.190 2377.660 1781.510 2377.720 ;
        RECT 1738.885 21.660 1739.175 21.705 ;
        RECT 1781.190 21.660 1781.510 21.720 ;
        RECT 1738.885 21.520 1781.510 21.660 ;
        RECT 1738.885 21.475 1739.175 21.520 ;
        RECT 1781.190 21.460 1781.510 21.520 ;
        RECT 1535.105 20.640 1535.395 20.685 ;
        RECT 1583.405 20.640 1583.695 20.685 ;
        RECT 1535.105 20.500 1583.695 20.640 ;
        RECT 1535.105 20.455 1535.395 20.500 ;
        RECT 1583.405 20.455 1583.695 20.500 ;
        RECT 1635.385 20.640 1635.675 20.685 ;
        RECT 1704.385 20.640 1704.675 20.685 ;
        RECT 1635.385 20.500 1704.675 20.640 ;
        RECT 1635.385 20.455 1635.675 20.500 ;
        RECT 1704.385 20.455 1704.675 20.500 ;
        RECT 1726.925 20.300 1727.215 20.345 ;
        RECT 1738.885 20.300 1739.175 20.345 ;
        RECT 1726.925 20.160 1739.175 20.300 ;
        RECT 1726.925 20.115 1727.215 20.160 ;
        RECT 1738.885 20.115 1739.175 20.160 ;
        RECT 1507.030 18.940 1507.350 19.000 ;
        RECT 1535.105 18.940 1535.395 18.985 ;
        RECT 1507.030 18.800 1535.395 18.940 ;
        RECT 1507.030 18.740 1507.350 18.800 ;
        RECT 1535.105 18.755 1535.395 18.800 ;
        RECT 1583.405 18.940 1583.695 18.985 ;
        RECT 1635.385 18.940 1635.675 18.985 ;
        RECT 1583.405 18.800 1635.675 18.940 ;
        RECT 1583.405 18.755 1583.695 18.800 ;
        RECT 1635.385 18.755 1635.675 18.800 ;
        RECT 1704.385 18.940 1704.675 18.985 ;
        RECT 1724.625 18.940 1724.915 18.985 ;
        RECT 1704.385 18.800 1724.915 18.940 ;
        RECT 1704.385 18.755 1704.675 18.800 ;
        RECT 1724.625 18.755 1724.915 18.800 ;
      LAYER via ;
        RECT 1451.400 2378.000 1451.660 2378.260 ;
        RECT 1781.220 2377.660 1781.480 2377.920 ;
        RECT 1781.220 21.460 1781.480 21.720 ;
        RECT 1507.060 18.740 1507.320 19.000 ;
      LAYER met2 ;
        RECT 1451.400 2377.970 1451.660 2378.290 ;
        RECT 1450.060 2377.690 1450.340 2377.880 ;
        RECT 1451.460 2377.690 1451.600 2377.970 ;
        RECT 1450.060 2377.550 1451.600 2377.690 ;
        RECT 1781.220 2377.630 1781.480 2377.950 ;
        RECT 1450.060 2373.880 1450.340 2377.550 ;
        RECT 1781.280 21.750 1781.420 2377.630 ;
        RECT 1781.220 21.430 1781.480 21.750 ;
        RECT 1507.060 18.710 1507.320 19.030 ;
        RECT 1507.120 2.400 1507.260 18.710 ;
        RECT 1506.910 -4.800 1507.470 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 707.090 1294.960 707.410 1295.020 ;
        RECT 718.590 1294.960 718.910 1295.020 ;
        RECT 707.090 1294.820 718.910 1294.960 ;
        RECT 707.090 1294.760 707.410 1294.820 ;
        RECT 718.590 1294.760 718.910 1294.820 ;
        RECT 704.330 20.640 704.650 20.700 ;
        RECT 707.090 20.640 707.410 20.700 ;
        RECT 704.330 20.500 707.410 20.640 ;
        RECT 704.330 20.440 704.650 20.500 ;
        RECT 707.090 20.440 707.410 20.500 ;
      LAYER via ;
        RECT 707.120 1294.760 707.380 1295.020 ;
        RECT 718.620 1294.760 718.880 1295.020 ;
        RECT 704.360 20.440 704.620 20.700 ;
        RECT 707.120 20.440 707.380 20.700 ;
      LAYER met2 ;
        RECT 718.660 1323.135 718.940 1327.135 ;
        RECT 718.680 1295.050 718.820 1323.135 ;
        RECT 707.120 1294.730 707.380 1295.050 ;
        RECT 718.620 1294.730 718.880 1295.050 ;
        RECT 707.180 20.730 707.320 1294.730 ;
        RECT 704.360 20.410 704.620 20.730 ;
        RECT 707.120 20.410 707.380 20.730 ;
        RECT 704.420 2.400 704.560 20.410 ;
        RECT 704.210 -4.800 704.770 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1524.970 27.440 1525.290 27.500 ;
        RECT 1758.650 27.440 1758.970 27.500 ;
        RECT 1524.970 27.300 1758.970 27.440 ;
        RECT 1524.970 27.240 1525.290 27.300 ;
        RECT 1758.650 27.240 1758.970 27.300 ;
      LAYER via ;
        RECT 1525.000 27.240 1525.260 27.500 ;
        RECT 1758.680 27.240 1758.940 27.500 ;
      LAYER met2 ;
        RECT 1758.670 2097.955 1758.950 2098.325 ;
        RECT 1758.740 1760.365 1758.880 2097.955 ;
        RECT 1758.670 1759.995 1758.950 1760.365 ;
        RECT 1758.670 1759.315 1758.950 1759.685 ;
        RECT 1758.740 27.530 1758.880 1759.315 ;
        RECT 1525.000 27.210 1525.260 27.530 ;
        RECT 1758.680 27.210 1758.940 27.530 ;
        RECT 1525.060 2.400 1525.200 27.210 ;
        RECT 1524.850 -4.800 1525.410 2.400 ;
      LAYER via2 ;
        RECT 1758.670 2098.000 1758.950 2098.280 ;
        RECT 1758.670 1760.040 1758.950 1760.320 ;
        RECT 1758.670 1759.360 1758.950 1759.640 ;
      LAYER met3 ;
        RECT 1755.835 2099.735 1759.835 2100.335 ;
        RECT 1758.430 2098.305 1758.730 2099.735 ;
        RECT 1758.430 2097.990 1758.975 2098.305 ;
        RECT 1758.645 2097.975 1758.975 2097.990 ;
        RECT 1758.645 1760.330 1758.975 1760.345 ;
        RECT 1758.430 1760.015 1758.975 1760.330 ;
        RECT 1758.430 1759.665 1758.730 1760.015 ;
        RECT 1758.430 1759.350 1758.975 1759.665 ;
        RECT 1758.645 1759.335 1758.975 1759.350 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 708.470 41.380 708.790 41.440 ;
        RECT 1542.910 41.380 1543.230 41.440 ;
        RECT 708.470 41.240 1543.230 41.380 ;
        RECT 708.470 41.180 708.790 41.240 ;
        RECT 1542.910 41.180 1543.230 41.240 ;
      LAYER via ;
        RECT 708.500 41.180 708.760 41.440 ;
        RECT 1542.940 41.180 1543.200 41.440 ;
      LAYER met2 ;
        RECT 708.490 1702.875 708.770 1703.245 ;
        RECT 708.560 41.470 708.700 1702.875 ;
        RECT 708.500 41.150 708.760 41.470 ;
        RECT 1542.940 41.150 1543.200 41.470 ;
        RECT 1543.000 2.400 1543.140 41.150 ;
        RECT 1542.790 -4.800 1543.350 2.400 ;
      LAYER via2 ;
        RECT 708.490 1702.920 708.770 1703.200 ;
      LAYER met3 ;
        RECT 708.465 1703.210 708.795 1703.225 ;
        RECT 715.810 1703.210 719.810 1703.215 ;
        RECT 708.465 1702.910 719.810 1703.210 ;
        RECT 708.465 1702.895 708.795 1702.910 ;
        RECT 715.810 1702.615 719.810 1702.910 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 775.630 1311.620 775.950 1311.680 ;
        RECT 779.310 1311.620 779.630 1311.680 ;
        RECT 775.630 1311.480 779.630 1311.620 ;
        RECT 775.630 1311.420 775.950 1311.480 ;
        RECT 779.310 1311.420 779.630 1311.480 ;
        RECT 779.310 25.060 779.630 25.120 ;
        RECT 1560.850 25.060 1561.170 25.120 ;
        RECT 779.310 24.920 1561.170 25.060 ;
        RECT 779.310 24.860 779.630 24.920 ;
        RECT 1560.850 24.860 1561.170 24.920 ;
      LAYER via ;
        RECT 775.660 1311.420 775.920 1311.680 ;
        RECT 779.340 1311.420 779.600 1311.680 ;
        RECT 779.340 24.860 779.600 25.120 ;
        RECT 1560.880 24.860 1561.140 25.120 ;
      LAYER met2 ;
        RECT 775.700 1323.135 775.980 1327.135 ;
        RECT 775.720 1311.710 775.860 1323.135 ;
        RECT 775.660 1311.390 775.920 1311.710 ;
        RECT 779.340 1311.390 779.600 1311.710 ;
        RECT 779.400 25.150 779.540 1311.390 ;
        RECT 779.340 24.830 779.600 25.150 ;
        RECT 1560.880 24.830 1561.140 25.150 ;
        RECT 1560.940 2.400 1561.080 24.830 ;
        RECT 1560.730 -4.800 1561.290 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1754.585 1605.905 1754.755 1628.515 ;
        RECT 1756.885 1484.185 1757.055 1524.475 ;
        RECT 1753.205 1242.445 1753.375 1245.335 ;
        RECT 1752.745 1193.825 1752.915 1241.935 ;
        RECT 1752.745 910.945 1752.915 931.855 ;
        RECT 1754.125 879.665 1754.295 903.975 ;
        RECT 1752.745 717.825 1752.915 765.935 ;
        RECT 1752.745 662.405 1752.915 669.715 ;
        RECT 1753.205 517.565 1753.375 565.335 ;
        RECT 1752.745 276.165 1752.915 324.275 ;
        RECT 1752.745 144.925 1752.915 207.315 ;
      LAYER mcon ;
        RECT 1754.585 1628.345 1754.755 1628.515 ;
        RECT 1756.885 1524.305 1757.055 1524.475 ;
        RECT 1753.205 1245.165 1753.375 1245.335 ;
        RECT 1752.745 1241.765 1752.915 1241.935 ;
        RECT 1752.745 931.685 1752.915 931.855 ;
        RECT 1754.125 903.805 1754.295 903.975 ;
        RECT 1752.745 765.765 1752.915 765.935 ;
        RECT 1752.745 669.545 1752.915 669.715 ;
        RECT 1753.205 565.165 1753.375 565.335 ;
        RECT 1752.745 324.105 1752.915 324.275 ;
        RECT 1752.745 207.145 1752.915 207.315 ;
      LAYER met1 ;
        RECT 1754.510 1805.980 1754.830 1806.040 ;
        RECT 1757.730 1805.980 1758.050 1806.040 ;
        RECT 1754.510 1805.840 1758.050 1805.980 ;
        RECT 1754.510 1805.780 1754.830 1805.840 ;
        RECT 1757.730 1805.780 1758.050 1805.840 ;
        RECT 1754.510 1628.500 1754.830 1628.560 ;
        RECT 1754.315 1628.360 1754.830 1628.500 ;
        RECT 1754.510 1628.300 1754.830 1628.360 ;
        RECT 1754.510 1606.060 1754.830 1606.120 ;
        RECT 1754.315 1605.920 1754.830 1606.060 ;
        RECT 1754.510 1605.860 1754.830 1605.920 ;
        RECT 1754.510 1524.460 1754.830 1524.520 ;
        RECT 1756.825 1524.460 1757.115 1524.505 ;
        RECT 1754.510 1524.320 1757.115 1524.460 ;
        RECT 1754.510 1524.260 1754.830 1524.320 ;
        RECT 1756.825 1524.275 1757.115 1524.320 ;
        RECT 1754.510 1484.340 1754.830 1484.400 ;
        RECT 1756.825 1484.340 1757.115 1484.385 ;
        RECT 1754.510 1484.200 1757.115 1484.340 ;
        RECT 1754.510 1484.140 1754.830 1484.200 ;
        RECT 1756.825 1484.155 1757.115 1484.200 ;
        RECT 1753.145 1245.320 1753.435 1245.365 ;
        RECT 1753.590 1245.320 1753.910 1245.380 ;
        RECT 1753.145 1245.180 1753.910 1245.320 ;
        RECT 1753.145 1245.135 1753.435 1245.180 ;
        RECT 1753.590 1245.120 1753.910 1245.180 ;
        RECT 1753.130 1242.600 1753.450 1242.660 ;
        RECT 1752.935 1242.460 1753.450 1242.600 ;
        RECT 1753.130 1242.400 1753.450 1242.460 ;
        RECT 1752.685 1241.920 1752.975 1241.965 ;
        RECT 1753.130 1241.920 1753.450 1241.980 ;
        RECT 1752.685 1241.780 1753.450 1241.920 ;
        RECT 1752.685 1241.735 1752.975 1241.780 ;
        RECT 1753.130 1241.720 1753.450 1241.780 ;
        RECT 1752.670 1193.980 1752.990 1194.040 ;
        RECT 1752.475 1193.840 1752.990 1193.980 ;
        RECT 1752.670 1193.780 1752.990 1193.840 ;
        RECT 1752.670 1014.460 1752.990 1014.520 ;
        RECT 1753.130 1014.460 1753.450 1014.520 ;
        RECT 1752.670 1014.320 1753.450 1014.460 ;
        RECT 1752.670 1014.260 1752.990 1014.320 ;
        RECT 1753.130 1014.260 1753.450 1014.320 ;
        RECT 1752.670 931.840 1752.990 931.900 ;
        RECT 1752.475 931.700 1752.990 931.840 ;
        RECT 1752.670 931.640 1752.990 931.700 ;
        RECT 1752.670 911.100 1752.990 911.160 ;
        RECT 1752.475 910.960 1752.990 911.100 ;
        RECT 1752.670 910.900 1752.990 910.960 ;
        RECT 1752.670 908.040 1752.990 908.100 ;
        RECT 1754.050 908.040 1754.370 908.100 ;
        RECT 1752.670 907.900 1754.370 908.040 ;
        RECT 1752.670 907.840 1752.990 907.900 ;
        RECT 1754.050 907.840 1754.370 907.900 ;
        RECT 1754.050 903.960 1754.370 904.020 ;
        RECT 1753.855 903.820 1754.370 903.960 ;
        RECT 1754.050 903.760 1754.370 903.820 ;
        RECT 1754.050 879.820 1754.370 879.880 ;
        RECT 1753.855 879.680 1754.370 879.820 ;
        RECT 1754.050 879.620 1754.370 879.680 ;
        RECT 1752.670 845.480 1752.990 845.540 ;
        RECT 1754.050 845.480 1754.370 845.540 ;
        RECT 1752.670 845.340 1754.370 845.480 ;
        RECT 1752.670 845.280 1752.990 845.340 ;
        RECT 1754.050 845.280 1754.370 845.340 ;
        RECT 1750.830 821.000 1751.150 821.060 ;
        RECT 1752.670 821.000 1752.990 821.060 ;
        RECT 1750.830 820.860 1752.990 821.000 ;
        RECT 1750.830 820.800 1751.150 820.860 ;
        RECT 1752.670 820.800 1752.990 820.860 ;
        RECT 1752.685 765.920 1752.975 765.965 ;
        RECT 1753.130 765.920 1753.450 765.980 ;
        RECT 1752.685 765.780 1753.450 765.920 ;
        RECT 1752.685 765.735 1752.975 765.780 ;
        RECT 1753.130 765.720 1753.450 765.780 ;
        RECT 1752.670 717.980 1752.990 718.040 ;
        RECT 1752.475 717.840 1752.990 717.980 ;
        RECT 1752.670 717.780 1752.990 717.840 ;
        RECT 1752.670 669.700 1752.990 669.760 ;
        RECT 1752.475 669.560 1752.990 669.700 ;
        RECT 1752.670 669.500 1752.990 669.560 ;
        RECT 1752.670 662.560 1752.990 662.620 ;
        RECT 1752.475 662.420 1752.990 662.560 ;
        RECT 1752.670 662.360 1752.990 662.420 ;
        RECT 1752.670 614.280 1752.990 614.340 ;
        RECT 1753.130 614.280 1753.450 614.340 ;
        RECT 1752.670 614.140 1753.450 614.280 ;
        RECT 1752.670 614.080 1752.990 614.140 ;
        RECT 1753.130 614.080 1753.450 614.140 ;
        RECT 1752.670 566.000 1752.990 566.060 ;
        RECT 1753.130 566.000 1753.450 566.060 ;
        RECT 1752.670 565.860 1753.450 566.000 ;
        RECT 1752.670 565.800 1752.990 565.860 ;
        RECT 1753.130 565.800 1753.450 565.860 ;
        RECT 1752.670 565.320 1752.990 565.380 ;
        RECT 1753.145 565.320 1753.435 565.365 ;
        RECT 1752.670 565.180 1753.435 565.320 ;
        RECT 1752.670 565.120 1752.990 565.180 ;
        RECT 1753.145 565.135 1753.435 565.180 ;
        RECT 1753.130 517.720 1753.450 517.780 ;
        RECT 1753.130 517.580 1753.645 517.720 ;
        RECT 1753.130 517.520 1753.450 517.580 ;
        RECT 1753.130 469.920 1753.450 470.180 ;
        RECT 1753.220 469.500 1753.360 469.920 ;
        RECT 1753.130 469.240 1753.450 469.500 ;
        RECT 1753.130 352.480 1753.450 352.540 ;
        RECT 1752.760 352.340 1753.450 352.480 ;
        RECT 1752.760 351.860 1752.900 352.340 ;
        RECT 1753.130 352.280 1753.450 352.340 ;
        RECT 1752.670 351.600 1752.990 351.860 ;
        RECT 1752.670 324.260 1752.990 324.320 ;
        RECT 1752.475 324.120 1752.990 324.260 ;
        RECT 1752.670 324.060 1752.990 324.120 ;
        RECT 1752.670 276.320 1752.990 276.380 ;
        RECT 1752.475 276.180 1752.990 276.320 ;
        RECT 1752.670 276.120 1752.990 276.180 ;
        RECT 1752.670 207.300 1752.990 207.360 ;
        RECT 1752.475 207.160 1752.990 207.300 ;
        RECT 1752.670 207.100 1752.990 207.160 ;
        RECT 1752.670 145.080 1752.990 145.140 ;
        RECT 1752.475 144.940 1752.990 145.080 ;
        RECT 1752.670 144.880 1752.990 144.940 ;
        RECT 1752.670 110.400 1752.990 110.460 ;
        RECT 1753.590 110.400 1753.910 110.460 ;
        RECT 1752.670 110.260 1753.910 110.400 ;
        RECT 1752.670 110.200 1752.990 110.260 ;
        RECT 1753.590 110.200 1753.910 110.260 ;
        RECT 1753.590 96.260 1753.910 96.520 ;
        RECT 1753.680 95.840 1753.820 96.260 ;
        RECT 1753.590 95.580 1753.910 95.840 ;
        RECT 1578.790 23.700 1579.110 23.760 ;
        RECT 1753.590 23.700 1753.910 23.760 ;
        RECT 1578.790 23.560 1753.910 23.700 ;
        RECT 1578.790 23.500 1579.110 23.560 ;
        RECT 1753.590 23.500 1753.910 23.560 ;
      LAYER via ;
        RECT 1754.540 1805.780 1754.800 1806.040 ;
        RECT 1757.760 1805.780 1758.020 1806.040 ;
        RECT 1754.540 1628.300 1754.800 1628.560 ;
        RECT 1754.540 1605.860 1754.800 1606.120 ;
        RECT 1754.540 1524.260 1754.800 1524.520 ;
        RECT 1754.540 1484.140 1754.800 1484.400 ;
        RECT 1753.620 1245.120 1753.880 1245.380 ;
        RECT 1753.160 1242.400 1753.420 1242.660 ;
        RECT 1753.160 1241.720 1753.420 1241.980 ;
        RECT 1752.700 1193.780 1752.960 1194.040 ;
        RECT 1752.700 1014.260 1752.960 1014.520 ;
        RECT 1753.160 1014.260 1753.420 1014.520 ;
        RECT 1752.700 931.640 1752.960 931.900 ;
        RECT 1752.700 910.900 1752.960 911.160 ;
        RECT 1752.700 907.840 1752.960 908.100 ;
        RECT 1754.080 907.840 1754.340 908.100 ;
        RECT 1754.080 903.760 1754.340 904.020 ;
        RECT 1754.080 879.620 1754.340 879.880 ;
        RECT 1752.700 845.280 1752.960 845.540 ;
        RECT 1754.080 845.280 1754.340 845.540 ;
        RECT 1750.860 820.800 1751.120 821.060 ;
        RECT 1752.700 820.800 1752.960 821.060 ;
        RECT 1753.160 765.720 1753.420 765.980 ;
        RECT 1752.700 717.780 1752.960 718.040 ;
        RECT 1752.700 669.500 1752.960 669.760 ;
        RECT 1752.700 662.360 1752.960 662.620 ;
        RECT 1752.700 614.080 1752.960 614.340 ;
        RECT 1753.160 614.080 1753.420 614.340 ;
        RECT 1752.700 565.800 1752.960 566.060 ;
        RECT 1753.160 565.800 1753.420 566.060 ;
        RECT 1752.700 565.120 1752.960 565.380 ;
        RECT 1753.160 517.520 1753.420 517.780 ;
        RECT 1753.160 469.920 1753.420 470.180 ;
        RECT 1753.160 469.240 1753.420 469.500 ;
        RECT 1753.160 352.280 1753.420 352.540 ;
        RECT 1752.700 351.600 1752.960 351.860 ;
        RECT 1752.700 324.060 1752.960 324.320 ;
        RECT 1752.700 276.120 1752.960 276.380 ;
        RECT 1752.700 207.100 1752.960 207.360 ;
        RECT 1752.700 144.880 1752.960 145.140 ;
        RECT 1752.700 110.200 1752.960 110.460 ;
        RECT 1753.620 110.200 1753.880 110.460 ;
        RECT 1753.620 96.260 1753.880 96.520 ;
        RECT 1753.620 95.580 1753.880 95.840 ;
        RECT 1578.820 23.500 1579.080 23.760 ;
        RECT 1753.620 23.500 1753.880 23.760 ;
      LAYER met2 ;
        RECT 1757.750 1832.075 1758.030 1832.445 ;
        RECT 1757.820 1806.070 1757.960 1832.075 ;
        RECT 1754.540 1805.980 1754.800 1806.070 ;
        RECT 1752.300 1805.840 1754.800 1805.980 ;
        RECT 1752.300 1784.050 1752.440 1805.840 ;
        RECT 1754.540 1805.750 1754.800 1805.840 ;
        RECT 1757.760 1805.750 1758.020 1806.070 ;
        RECT 1752.300 1783.910 1752.900 1784.050 ;
        RECT 1752.760 1782.690 1752.900 1783.910 ;
        RECT 1752.760 1782.550 1753.820 1782.690 ;
        RECT 1753.680 1758.890 1753.820 1782.550 ;
        RECT 1752.760 1758.750 1753.820 1758.890 ;
        RECT 1752.760 1752.090 1752.900 1758.750 ;
        RECT 1752.760 1751.950 1754.280 1752.090 ;
        RECT 1754.140 1705.170 1754.280 1751.950 ;
        RECT 1753.220 1705.030 1754.280 1705.170 ;
        RECT 1753.220 1628.500 1753.360 1705.030 ;
        RECT 1754.540 1628.500 1754.800 1628.590 ;
        RECT 1753.220 1628.360 1754.800 1628.500 ;
        RECT 1754.540 1628.270 1754.800 1628.360 ;
        RECT 1754.540 1605.890 1754.800 1606.150 ;
        RECT 1753.220 1605.830 1754.800 1605.890 ;
        RECT 1753.220 1605.750 1754.740 1605.830 ;
        RECT 1753.220 1582.770 1753.360 1605.750 ;
        RECT 1753.220 1582.630 1753.820 1582.770 ;
        RECT 1753.680 1524.460 1753.820 1582.630 ;
        RECT 1754.540 1524.460 1754.800 1524.550 ;
        RECT 1753.680 1524.320 1754.800 1524.460 ;
        RECT 1754.540 1524.230 1754.800 1524.320 ;
        RECT 1754.540 1484.170 1754.800 1484.430 ;
        RECT 1753.220 1484.110 1754.800 1484.170 ;
        RECT 1753.220 1484.030 1754.740 1484.110 ;
        RECT 1753.220 1293.770 1753.360 1484.030 ;
        RECT 1753.220 1293.630 1753.820 1293.770 ;
        RECT 1753.680 1245.410 1753.820 1293.630 ;
        RECT 1753.620 1245.090 1753.880 1245.410 ;
        RECT 1753.160 1242.370 1753.420 1242.690 ;
        RECT 1753.220 1242.010 1753.360 1242.370 ;
        RECT 1753.160 1241.690 1753.420 1242.010 ;
        RECT 1752.700 1193.750 1752.960 1194.070 ;
        RECT 1752.760 1104.165 1752.900 1193.750 ;
        RECT 1752.690 1103.795 1752.970 1104.165 ;
        RECT 1753.150 1103.115 1753.430 1103.485 ;
        RECT 1753.220 1014.550 1753.360 1103.115 ;
        RECT 1752.700 1014.230 1752.960 1014.550 ;
        RECT 1753.160 1014.230 1753.420 1014.550 ;
        RECT 1752.760 931.930 1752.900 1014.230 ;
        RECT 1752.700 931.610 1752.960 931.930 ;
        RECT 1752.700 910.870 1752.960 911.190 ;
        RECT 1752.760 908.130 1752.900 910.870 ;
        RECT 1752.700 907.810 1752.960 908.130 ;
        RECT 1754.080 907.810 1754.340 908.130 ;
        RECT 1754.140 904.050 1754.280 907.810 ;
        RECT 1754.080 903.730 1754.340 904.050 ;
        RECT 1754.080 879.590 1754.340 879.910 ;
        RECT 1754.140 845.570 1754.280 879.590 ;
        RECT 1752.700 845.250 1752.960 845.570 ;
        RECT 1754.080 845.250 1754.340 845.570 ;
        RECT 1752.760 821.090 1752.900 845.250 ;
        RECT 1750.860 820.770 1751.120 821.090 ;
        RECT 1752.700 820.770 1752.960 821.090 ;
        RECT 1750.920 766.205 1751.060 820.770 ;
        RECT 1750.850 765.835 1751.130 766.205 ;
        RECT 1753.150 765.835 1753.430 766.205 ;
        RECT 1753.160 765.690 1753.420 765.835 ;
        RECT 1752.700 717.750 1752.960 718.070 ;
        RECT 1752.760 669.790 1752.900 717.750 ;
        RECT 1752.700 669.470 1752.960 669.790 ;
        RECT 1752.700 662.330 1752.960 662.650 ;
        RECT 1752.760 614.370 1752.900 662.330 ;
        RECT 1752.700 614.050 1752.960 614.370 ;
        RECT 1753.160 614.050 1753.420 614.370 ;
        RECT 1753.220 566.090 1753.360 614.050 ;
        RECT 1752.700 565.770 1752.960 566.090 ;
        RECT 1753.160 565.770 1753.420 566.090 ;
        RECT 1752.760 565.410 1752.900 565.770 ;
        RECT 1752.700 565.090 1752.960 565.410 ;
        RECT 1753.160 517.490 1753.420 517.810 ;
        RECT 1753.220 470.210 1753.360 517.490 ;
        RECT 1753.160 469.890 1753.420 470.210 ;
        RECT 1753.160 469.210 1753.420 469.530 ;
        RECT 1753.220 352.570 1753.360 469.210 ;
        RECT 1753.160 352.250 1753.420 352.570 ;
        RECT 1752.700 351.570 1752.960 351.890 ;
        RECT 1752.760 324.350 1752.900 351.570 ;
        RECT 1752.700 324.030 1752.960 324.350 ;
        RECT 1752.700 276.090 1752.960 276.410 ;
        RECT 1752.760 207.390 1752.900 276.090 ;
        RECT 1752.700 207.070 1752.960 207.390 ;
        RECT 1752.700 144.850 1752.960 145.170 ;
        RECT 1752.760 110.490 1752.900 144.850 ;
        RECT 1752.700 110.170 1752.960 110.490 ;
        RECT 1753.620 110.170 1753.880 110.490 ;
        RECT 1753.680 96.550 1753.820 110.170 ;
        RECT 1753.620 96.230 1753.880 96.550 ;
        RECT 1753.620 95.550 1753.880 95.870 ;
        RECT 1753.680 23.790 1753.820 95.550 ;
        RECT 1578.820 23.470 1579.080 23.790 ;
        RECT 1753.620 23.470 1753.880 23.790 ;
        RECT 1578.880 2.400 1579.020 23.470 ;
        RECT 1578.670 -4.800 1579.230 2.400 ;
      LAYER via2 ;
        RECT 1757.750 1832.120 1758.030 1832.400 ;
        RECT 1752.690 1103.840 1752.970 1104.120 ;
        RECT 1753.150 1103.160 1753.430 1103.440 ;
        RECT 1750.850 765.880 1751.130 766.160 ;
        RECT 1753.150 765.880 1753.430 766.160 ;
      LAYER met3 ;
        RECT 1755.835 1834.535 1759.835 1835.135 ;
        RECT 1757.510 1832.425 1757.810 1834.535 ;
        RECT 1757.510 1832.110 1758.055 1832.425 ;
        RECT 1757.725 1832.095 1758.055 1832.110 ;
        RECT 1752.665 1104.130 1752.995 1104.145 ;
        RECT 1752.665 1103.815 1753.210 1104.130 ;
        RECT 1752.910 1103.465 1753.210 1103.815 ;
        RECT 1752.910 1103.150 1753.455 1103.465 ;
        RECT 1753.125 1103.135 1753.455 1103.150 ;
        RECT 1750.825 766.170 1751.155 766.185 ;
        RECT 1753.125 766.170 1753.455 766.185 ;
        RECT 1750.825 765.870 1753.455 766.170 ;
        RECT 1750.825 765.855 1751.155 765.870 ;
        RECT 1753.125 765.855 1753.455 765.870 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1479.450 2380.155 1479.730 2380.525 ;
        RECT 1479.520 2377.880 1479.660 2380.155 ;
        RECT 1479.500 2373.880 1479.780 2377.880 ;
        RECT 1596.290 13.755 1596.570 14.125 ;
        RECT 1596.360 2.400 1596.500 13.755 ;
        RECT 1596.150 -4.800 1596.710 2.400 ;
      LAYER via2 ;
        RECT 1479.450 2380.200 1479.730 2380.480 ;
        RECT 1596.290 13.800 1596.570 14.080 ;
      LAYER met3 ;
        RECT 1479.425 2380.490 1479.755 2380.505 ;
        RECT 1745.510 2380.490 1745.890 2380.500 ;
        RECT 1479.425 2380.190 1745.890 2380.490 ;
        RECT 1479.425 2380.175 1479.755 2380.190 ;
        RECT 1745.510 2380.180 1745.890 2380.190 ;
        RECT 1596.265 14.090 1596.595 14.105 ;
        RECT 1745.510 14.090 1745.890 14.100 ;
        RECT 1596.265 13.790 1745.890 14.090 ;
        RECT 1596.265 13.775 1596.595 13.790 ;
        RECT 1745.510 13.780 1745.890 13.790 ;
      LAYER via3 ;
        RECT 1745.540 2380.180 1745.860 2380.500 ;
        RECT 1745.540 13.780 1745.860 14.100 ;
      LAYER met4 ;
        RECT 1745.535 2380.175 1745.865 2380.505 ;
        RECT 1745.550 14.105 1745.850 2380.175 ;
        RECT 1745.535 13.775 1745.865 14.105 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1613.825 862.665 1613.995 910.435 ;
        RECT 1613.825 766.105 1613.995 814.215 ;
        RECT 1613.825 669.545 1613.995 717.655 ;
        RECT 1613.825 572.645 1613.995 620.755 ;
        RECT 1613.825 476.085 1613.995 524.195 ;
        RECT 1613.825 379.525 1613.995 427.635 ;
        RECT 1613.825 282.965 1613.995 331.075 ;
        RECT 1613.825 186.405 1613.995 234.515 ;
        RECT 1613.825 89.845 1613.995 137.955 ;
        RECT 1613.365 48.705 1613.535 62.475 ;
        RECT 1614.285 17.425 1614.455 48.195 ;
      LAYER mcon ;
        RECT 1613.825 910.265 1613.995 910.435 ;
        RECT 1613.825 814.045 1613.995 814.215 ;
        RECT 1613.825 717.485 1613.995 717.655 ;
        RECT 1613.825 620.585 1613.995 620.755 ;
        RECT 1613.825 524.025 1613.995 524.195 ;
        RECT 1613.825 427.465 1613.995 427.635 ;
        RECT 1613.825 330.905 1613.995 331.075 ;
        RECT 1613.825 234.345 1613.995 234.515 ;
        RECT 1613.825 137.785 1613.995 137.955 ;
        RECT 1613.365 62.305 1613.535 62.475 ;
        RECT 1614.285 48.025 1614.455 48.195 ;
      LAYER met1 ;
        RECT 1692.870 2392.140 1693.190 2392.200 ;
        RECT 1782.110 2392.140 1782.430 2392.200 ;
        RECT 1692.870 2392.000 1782.430 2392.140 ;
        RECT 1692.870 2391.940 1693.190 2392.000 ;
        RECT 1782.110 2391.940 1782.430 2392.000 ;
        RECT 1782.110 1327.260 1782.430 1327.320 ;
        RECT 1613.840 1327.120 1782.430 1327.260 ;
        RECT 1613.840 1326.640 1613.980 1327.120 ;
        RECT 1782.110 1327.060 1782.430 1327.120 ;
        RECT 1613.750 1326.380 1614.070 1326.640 ;
        RECT 1612.830 1249.060 1613.150 1249.120 ;
        RECT 1613.750 1249.060 1614.070 1249.120 ;
        RECT 1612.830 1248.920 1614.070 1249.060 ;
        RECT 1612.830 1248.860 1613.150 1248.920 ;
        RECT 1613.750 1248.860 1614.070 1248.920 ;
        RECT 1612.830 1152.500 1613.150 1152.560 ;
        RECT 1613.750 1152.500 1614.070 1152.560 ;
        RECT 1612.830 1152.360 1614.070 1152.500 ;
        RECT 1612.830 1152.300 1613.150 1152.360 ;
        RECT 1613.750 1152.300 1614.070 1152.360 ;
        RECT 1612.830 1007.320 1613.150 1007.380 ;
        RECT 1613.750 1007.320 1614.070 1007.380 ;
        RECT 1612.830 1007.180 1614.070 1007.320 ;
        RECT 1612.830 1007.120 1613.150 1007.180 ;
        RECT 1613.750 1007.120 1614.070 1007.180 ;
        RECT 1613.750 910.420 1614.070 910.480 ;
        RECT 1613.555 910.280 1614.070 910.420 ;
        RECT 1613.750 910.220 1614.070 910.280 ;
        RECT 1613.750 862.820 1614.070 862.880 ;
        RECT 1613.555 862.680 1614.070 862.820 ;
        RECT 1613.750 862.620 1614.070 862.680 ;
        RECT 1613.750 814.200 1614.070 814.260 ;
        RECT 1613.555 814.060 1614.070 814.200 ;
        RECT 1613.750 814.000 1614.070 814.060 ;
        RECT 1613.750 766.260 1614.070 766.320 ;
        RECT 1613.555 766.120 1614.070 766.260 ;
        RECT 1613.750 766.060 1614.070 766.120 ;
        RECT 1613.750 717.640 1614.070 717.700 ;
        RECT 1613.555 717.500 1614.070 717.640 ;
        RECT 1613.750 717.440 1614.070 717.500 ;
        RECT 1613.750 669.700 1614.070 669.760 ;
        RECT 1613.555 669.560 1614.070 669.700 ;
        RECT 1613.750 669.500 1614.070 669.560 ;
        RECT 1613.750 620.740 1614.070 620.800 ;
        RECT 1613.555 620.600 1614.070 620.740 ;
        RECT 1613.750 620.540 1614.070 620.600 ;
        RECT 1613.750 572.800 1614.070 572.860 ;
        RECT 1613.555 572.660 1614.070 572.800 ;
        RECT 1613.750 572.600 1614.070 572.660 ;
        RECT 1613.750 524.180 1614.070 524.240 ;
        RECT 1613.555 524.040 1614.070 524.180 ;
        RECT 1613.750 523.980 1614.070 524.040 ;
        RECT 1613.750 476.240 1614.070 476.300 ;
        RECT 1613.555 476.100 1614.070 476.240 ;
        RECT 1613.750 476.040 1614.070 476.100 ;
        RECT 1613.750 427.620 1614.070 427.680 ;
        RECT 1613.555 427.480 1614.070 427.620 ;
        RECT 1613.750 427.420 1614.070 427.480 ;
        RECT 1613.750 379.680 1614.070 379.740 ;
        RECT 1613.555 379.540 1614.070 379.680 ;
        RECT 1613.750 379.480 1614.070 379.540 ;
        RECT 1613.750 331.060 1614.070 331.120 ;
        RECT 1613.555 330.920 1614.070 331.060 ;
        RECT 1613.750 330.860 1614.070 330.920 ;
        RECT 1613.750 283.120 1614.070 283.180 ;
        RECT 1613.555 282.980 1614.070 283.120 ;
        RECT 1613.750 282.920 1614.070 282.980 ;
        RECT 1613.750 234.500 1614.070 234.560 ;
        RECT 1613.555 234.360 1614.070 234.500 ;
        RECT 1613.750 234.300 1614.070 234.360 ;
        RECT 1613.750 186.560 1614.070 186.620 ;
        RECT 1613.555 186.420 1614.070 186.560 ;
        RECT 1613.750 186.360 1614.070 186.420 ;
        RECT 1613.750 137.940 1614.070 138.000 ;
        RECT 1613.555 137.800 1614.070 137.940 ;
        RECT 1613.750 137.740 1614.070 137.800 ;
        RECT 1613.750 90.000 1614.070 90.060 ;
        RECT 1613.555 89.860 1614.070 90.000 ;
        RECT 1613.750 89.800 1614.070 89.860 ;
        RECT 1613.305 62.460 1613.595 62.505 ;
        RECT 1613.750 62.460 1614.070 62.520 ;
        RECT 1613.305 62.320 1614.070 62.460 ;
        RECT 1613.305 62.275 1613.595 62.320 ;
        RECT 1613.750 62.260 1614.070 62.320 ;
        RECT 1613.290 48.860 1613.610 48.920 ;
        RECT 1613.095 48.720 1613.610 48.860 ;
        RECT 1613.290 48.660 1613.610 48.720 ;
        RECT 1613.290 48.180 1613.610 48.240 ;
        RECT 1614.225 48.180 1614.515 48.225 ;
        RECT 1613.290 48.040 1614.515 48.180 ;
        RECT 1613.290 47.980 1613.610 48.040 ;
        RECT 1614.225 47.995 1614.515 48.040 ;
        RECT 1614.210 17.580 1614.530 17.640 ;
        RECT 1614.015 17.440 1614.530 17.580 ;
        RECT 1614.210 17.380 1614.530 17.440 ;
      LAYER via ;
        RECT 1692.900 2391.940 1693.160 2392.200 ;
        RECT 1782.140 2391.940 1782.400 2392.200 ;
        RECT 1782.140 1327.060 1782.400 1327.320 ;
        RECT 1613.780 1326.380 1614.040 1326.640 ;
        RECT 1612.860 1248.860 1613.120 1249.120 ;
        RECT 1613.780 1248.860 1614.040 1249.120 ;
        RECT 1612.860 1152.300 1613.120 1152.560 ;
        RECT 1613.780 1152.300 1614.040 1152.560 ;
        RECT 1612.860 1007.120 1613.120 1007.380 ;
        RECT 1613.780 1007.120 1614.040 1007.380 ;
        RECT 1613.780 910.220 1614.040 910.480 ;
        RECT 1613.780 862.620 1614.040 862.880 ;
        RECT 1613.780 814.000 1614.040 814.260 ;
        RECT 1613.780 766.060 1614.040 766.320 ;
        RECT 1613.780 717.440 1614.040 717.700 ;
        RECT 1613.780 669.500 1614.040 669.760 ;
        RECT 1613.780 620.540 1614.040 620.800 ;
        RECT 1613.780 572.600 1614.040 572.860 ;
        RECT 1613.780 523.980 1614.040 524.240 ;
        RECT 1613.780 476.040 1614.040 476.300 ;
        RECT 1613.780 427.420 1614.040 427.680 ;
        RECT 1613.780 379.480 1614.040 379.740 ;
        RECT 1613.780 330.860 1614.040 331.120 ;
        RECT 1613.780 282.920 1614.040 283.180 ;
        RECT 1613.780 234.300 1614.040 234.560 ;
        RECT 1613.780 186.360 1614.040 186.620 ;
        RECT 1613.780 137.740 1614.040 138.000 ;
        RECT 1613.780 89.800 1614.040 90.060 ;
        RECT 1613.780 62.260 1614.040 62.520 ;
        RECT 1613.320 48.660 1613.580 48.920 ;
        RECT 1613.320 47.980 1613.580 48.240 ;
        RECT 1614.240 17.380 1614.500 17.640 ;
      LAYER met2 ;
        RECT 1692.900 2391.910 1693.160 2392.230 ;
        RECT 1782.140 2391.910 1782.400 2392.230 ;
        RECT 1692.960 2377.880 1693.100 2391.910 ;
        RECT 1692.940 2373.880 1693.220 2377.880 ;
        RECT 1782.200 1327.350 1782.340 2391.910 ;
        RECT 1782.140 1327.030 1782.400 1327.350 ;
        RECT 1613.780 1326.350 1614.040 1326.670 ;
        RECT 1613.840 1297.285 1613.980 1326.350 ;
        RECT 1612.850 1296.915 1613.130 1297.285 ;
        RECT 1613.770 1296.915 1614.050 1297.285 ;
        RECT 1612.920 1249.150 1613.060 1296.915 ;
        RECT 1612.860 1248.830 1613.120 1249.150 ;
        RECT 1613.780 1248.830 1614.040 1249.150 ;
        RECT 1613.840 1200.725 1613.980 1248.830 ;
        RECT 1612.850 1200.355 1613.130 1200.725 ;
        RECT 1613.770 1200.355 1614.050 1200.725 ;
        RECT 1612.920 1152.590 1613.060 1200.355 ;
        RECT 1612.860 1152.270 1613.120 1152.590 ;
        RECT 1613.780 1152.270 1614.040 1152.590 ;
        RECT 1613.840 1104.165 1613.980 1152.270 ;
        RECT 1612.850 1103.795 1613.130 1104.165 ;
        RECT 1613.770 1103.795 1614.050 1104.165 ;
        RECT 1612.920 1055.885 1613.060 1103.795 ;
        RECT 1612.850 1055.515 1613.130 1055.885 ;
        RECT 1613.770 1055.515 1614.050 1055.885 ;
        RECT 1613.840 1007.410 1613.980 1055.515 ;
        RECT 1612.860 1007.090 1613.120 1007.410 ;
        RECT 1613.780 1007.090 1614.040 1007.410 ;
        RECT 1612.920 959.325 1613.060 1007.090 ;
        RECT 1612.850 958.955 1613.130 959.325 ;
        RECT 1613.770 958.955 1614.050 959.325 ;
        RECT 1613.840 910.510 1613.980 958.955 ;
        RECT 1613.780 910.190 1614.040 910.510 ;
        RECT 1613.780 862.590 1614.040 862.910 ;
        RECT 1613.840 814.290 1613.980 862.590 ;
        RECT 1613.780 813.970 1614.040 814.290 ;
        RECT 1613.780 766.030 1614.040 766.350 ;
        RECT 1613.840 717.730 1613.980 766.030 ;
        RECT 1613.780 717.410 1614.040 717.730 ;
        RECT 1613.780 669.470 1614.040 669.790 ;
        RECT 1613.840 620.830 1613.980 669.470 ;
        RECT 1613.780 620.510 1614.040 620.830 ;
        RECT 1613.780 572.570 1614.040 572.890 ;
        RECT 1613.840 524.270 1613.980 572.570 ;
        RECT 1613.780 523.950 1614.040 524.270 ;
        RECT 1613.780 476.010 1614.040 476.330 ;
        RECT 1613.840 427.710 1613.980 476.010 ;
        RECT 1613.780 427.390 1614.040 427.710 ;
        RECT 1613.780 379.450 1614.040 379.770 ;
        RECT 1613.840 331.150 1613.980 379.450 ;
        RECT 1613.780 330.830 1614.040 331.150 ;
        RECT 1613.780 282.890 1614.040 283.210 ;
        RECT 1613.840 234.590 1613.980 282.890 ;
        RECT 1613.780 234.270 1614.040 234.590 ;
        RECT 1613.780 186.330 1614.040 186.650 ;
        RECT 1613.840 138.030 1613.980 186.330 ;
        RECT 1613.780 137.710 1614.040 138.030 ;
        RECT 1613.780 89.770 1614.040 90.090 ;
        RECT 1613.840 62.550 1613.980 89.770 ;
        RECT 1613.780 62.230 1614.040 62.550 ;
        RECT 1613.320 48.630 1613.580 48.950 ;
        RECT 1613.380 48.270 1613.520 48.630 ;
        RECT 1613.320 47.950 1613.580 48.270 ;
        RECT 1614.240 17.350 1614.500 17.670 ;
        RECT 1614.300 2.400 1614.440 17.350 ;
        RECT 1614.090 -4.800 1614.650 2.400 ;
      LAYER via2 ;
        RECT 1612.850 1296.960 1613.130 1297.240 ;
        RECT 1613.770 1296.960 1614.050 1297.240 ;
        RECT 1612.850 1200.400 1613.130 1200.680 ;
        RECT 1613.770 1200.400 1614.050 1200.680 ;
        RECT 1612.850 1103.840 1613.130 1104.120 ;
        RECT 1613.770 1103.840 1614.050 1104.120 ;
        RECT 1612.850 1055.560 1613.130 1055.840 ;
        RECT 1613.770 1055.560 1614.050 1055.840 ;
        RECT 1612.850 959.000 1613.130 959.280 ;
        RECT 1613.770 959.000 1614.050 959.280 ;
      LAYER met3 ;
        RECT 1612.825 1297.250 1613.155 1297.265 ;
        RECT 1613.745 1297.250 1614.075 1297.265 ;
        RECT 1612.825 1296.950 1614.075 1297.250 ;
        RECT 1612.825 1296.935 1613.155 1296.950 ;
        RECT 1613.745 1296.935 1614.075 1296.950 ;
        RECT 1612.825 1200.690 1613.155 1200.705 ;
        RECT 1613.745 1200.690 1614.075 1200.705 ;
        RECT 1612.825 1200.390 1614.075 1200.690 ;
        RECT 1612.825 1200.375 1613.155 1200.390 ;
        RECT 1613.745 1200.375 1614.075 1200.390 ;
        RECT 1612.825 1104.130 1613.155 1104.145 ;
        RECT 1613.745 1104.130 1614.075 1104.145 ;
        RECT 1612.825 1103.830 1614.075 1104.130 ;
        RECT 1612.825 1103.815 1613.155 1103.830 ;
        RECT 1613.745 1103.815 1614.075 1103.830 ;
        RECT 1612.825 1055.850 1613.155 1055.865 ;
        RECT 1613.745 1055.850 1614.075 1055.865 ;
        RECT 1612.825 1055.550 1614.075 1055.850 ;
        RECT 1612.825 1055.535 1613.155 1055.550 ;
        RECT 1613.745 1055.535 1614.075 1055.550 ;
        RECT 1612.825 959.290 1613.155 959.305 ;
        RECT 1613.745 959.290 1614.075 959.305 ;
        RECT 1612.825 958.990 1614.075 959.290 ;
        RECT 1612.825 958.975 1613.155 958.990 ;
        RECT 1613.745 958.975 1614.075 958.990 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1755.890 2277.220 1756.210 2277.280 ;
        RECT 1756.810 2277.220 1757.130 2277.280 ;
        RECT 1755.890 2277.080 1757.130 2277.220 ;
        RECT 1755.890 2277.020 1756.210 2277.080 ;
        RECT 1756.810 2277.020 1757.130 2277.080 ;
        RECT 1755.890 1342.220 1756.210 1342.280 ;
        RECT 1759.110 1342.220 1759.430 1342.280 ;
        RECT 1755.890 1342.080 1759.430 1342.220 ;
        RECT 1755.890 1342.020 1756.210 1342.080 ;
        RECT 1759.110 1342.020 1759.430 1342.080 ;
        RECT 1634.910 1293.940 1635.230 1294.000 ;
        RECT 1759.110 1293.940 1759.430 1294.000 ;
        RECT 1634.910 1293.800 1759.430 1293.940 ;
        RECT 1634.910 1293.740 1635.230 1293.800 ;
        RECT 1759.110 1293.740 1759.430 1293.800 ;
        RECT 1632.150 20.640 1632.470 20.700 ;
        RECT 1634.910 20.640 1635.230 20.700 ;
        RECT 1632.150 20.500 1635.230 20.640 ;
        RECT 1632.150 20.440 1632.470 20.500 ;
        RECT 1634.910 20.440 1635.230 20.500 ;
      LAYER via ;
        RECT 1755.920 2277.020 1756.180 2277.280 ;
        RECT 1756.840 2277.020 1757.100 2277.280 ;
        RECT 1755.920 1342.020 1756.180 1342.280 ;
        RECT 1759.140 1342.020 1759.400 1342.280 ;
        RECT 1634.940 1293.740 1635.200 1294.000 ;
        RECT 1759.140 1293.740 1759.400 1294.000 ;
        RECT 1632.180 20.440 1632.440 20.700 ;
        RECT 1634.940 20.440 1635.200 20.700 ;
      LAYER met2 ;
        RECT 1756.830 2277.475 1757.110 2277.845 ;
        RECT 1756.900 2277.310 1757.040 2277.475 ;
        RECT 1755.920 2276.990 1756.180 2277.310 ;
        RECT 1756.840 2276.990 1757.100 2277.310 ;
        RECT 1755.980 1342.310 1756.120 2276.990 ;
        RECT 1755.920 1341.990 1756.180 1342.310 ;
        RECT 1759.140 1341.990 1759.400 1342.310 ;
        RECT 1759.200 1294.030 1759.340 1341.990 ;
        RECT 1634.940 1293.710 1635.200 1294.030 ;
        RECT 1759.140 1293.710 1759.400 1294.030 ;
        RECT 1635.000 20.730 1635.140 1293.710 ;
        RECT 1632.180 20.410 1632.440 20.730 ;
        RECT 1634.940 20.410 1635.200 20.730 ;
        RECT 1632.240 2.400 1632.380 20.410 ;
        RECT 1632.030 -4.800 1632.590 2.400 ;
      LAYER via2 ;
        RECT 1756.830 2277.520 1757.110 2277.800 ;
      LAYER met3 ;
        RECT 1755.835 2279.255 1759.835 2279.855 ;
        RECT 1756.590 2277.825 1756.890 2279.255 ;
        RECT 1756.590 2277.510 1757.135 2277.825 ;
        RECT 1756.805 2277.495 1757.135 2277.510 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1755.965 1476.705 1756.135 1499.315 ;
      LAYER mcon ;
        RECT 1755.965 1499.145 1756.135 1499.315 ;
      LAYER met1 ;
        RECT 1755.430 2311.900 1755.750 2311.960 ;
        RECT 1757.270 2311.900 1757.590 2311.960 ;
        RECT 1755.430 2311.760 1757.590 2311.900 ;
        RECT 1755.430 2311.700 1755.750 2311.760 ;
        RECT 1757.270 2311.700 1757.590 2311.760 ;
        RECT 1755.430 1499.300 1755.750 1499.360 ;
        RECT 1755.905 1499.300 1756.195 1499.345 ;
        RECT 1755.430 1499.160 1756.195 1499.300 ;
        RECT 1755.430 1499.100 1755.750 1499.160 ;
        RECT 1755.905 1499.115 1756.195 1499.160 ;
        RECT 1755.430 1476.860 1755.750 1476.920 ;
        RECT 1755.905 1476.860 1756.195 1476.905 ;
        RECT 1755.430 1476.720 1756.195 1476.860 ;
        RECT 1755.430 1476.660 1755.750 1476.720 ;
        RECT 1755.905 1476.675 1756.195 1476.720 ;
        RECT 1655.610 1308.900 1655.930 1308.960 ;
        RECT 1755.430 1308.900 1755.750 1308.960 ;
        RECT 1655.610 1308.760 1755.750 1308.900 ;
        RECT 1655.610 1308.700 1655.930 1308.760 ;
        RECT 1755.430 1308.700 1755.750 1308.760 ;
        RECT 1650.090 18.940 1650.410 19.000 ;
        RECT 1655.610 18.940 1655.930 19.000 ;
        RECT 1650.090 18.800 1655.930 18.940 ;
        RECT 1650.090 18.740 1650.410 18.800 ;
        RECT 1655.610 18.740 1655.930 18.800 ;
      LAYER via ;
        RECT 1755.460 2311.700 1755.720 2311.960 ;
        RECT 1757.300 2311.700 1757.560 2311.960 ;
        RECT 1755.460 1499.100 1755.720 1499.360 ;
        RECT 1755.460 1476.660 1755.720 1476.920 ;
        RECT 1655.640 1308.700 1655.900 1308.960 ;
        RECT 1755.460 1308.700 1755.720 1308.960 ;
        RECT 1650.120 18.740 1650.380 19.000 ;
        RECT 1655.640 18.740 1655.900 19.000 ;
      LAYER met2 ;
        RECT 1757.290 2312.155 1757.570 2312.525 ;
        RECT 1757.360 2311.990 1757.500 2312.155 ;
        RECT 1755.460 2311.670 1755.720 2311.990 ;
        RECT 1757.300 2311.670 1757.560 2311.990 ;
        RECT 1755.520 1499.390 1755.660 2311.670 ;
        RECT 1755.460 1499.070 1755.720 1499.390 ;
        RECT 1755.460 1476.630 1755.720 1476.950 ;
        RECT 1755.520 1308.990 1755.660 1476.630 ;
        RECT 1655.640 1308.670 1655.900 1308.990 ;
        RECT 1755.460 1308.670 1755.720 1308.990 ;
        RECT 1655.700 19.030 1655.840 1308.670 ;
        RECT 1650.120 18.710 1650.380 19.030 ;
        RECT 1655.640 18.710 1655.900 19.030 ;
        RECT 1650.180 2.400 1650.320 18.710 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
      LAYER via2 ;
        RECT 1757.290 2312.200 1757.570 2312.480 ;
      LAYER met3 ;
        RECT 1755.835 2313.255 1759.835 2313.855 ;
        RECT 1757.510 2312.505 1757.810 2313.255 ;
        RECT 1757.265 2312.190 1757.810 2312.505 ;
        RECT 1757.265 2312.175 1757.595 2312.190 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1600.410 26.080 1600.730 26.140 ;
        RECT 1668.030 26.080 1668.350 26.140 ;
        RECT 1600.410 25.940 1668.350 26.080 ;
        RECT 1600.410 25.880 1600.730 25.940 ;
        RECT 1668.030 25.880 1668.350 25.940 ;
      LAYER via ;
        RECT 1600.440 25.880 1600.700 26.140 ;
        RECT 1668.060 25.880 1668.320 26.140 ;
      LAYER met2 ;
        RECT 1597.260 1323.690 1597.540 1327.135 ;
        RECT 1597.260 1323.550 1600.640 1323.690 ;
        RECT 1597.260 1323.135 1597.540 1323.550 ;
        RECT 1600.500 26.170 1600.640 1323.550 ;
        RECT 1600.440 25.850 1600.700 26.170 ;
        RECT 1668.060 25.850 1668.320 26.170 ;
        RECT 1668.120 2.400 1668.260 25.850 ;
        RECT 1667.910 -4.800 1668.470 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1684.205 338.045 1684.375 386.155 ;
        RECT 1684.205 241.485 1684.375 289.595 ;
        RECT 1683.745 131.665 1683.915 179.435 ;
        RECT 1684.205 34.425 1684.375 82.875 ;
      LAYER mcon ;
        RECT 1684.205 385.985 1684.375 386.155 ;
        RECT 1684.205 289.425 1684.375 289.595 ;
        RECT 1683.745 179.265 1683.915 179.435 ;
        RECT 1684.205 82.705 1684.375 82.875 ;
      LAYER met1 ;
        RECT 1684.590 1256.200 1684.910 1256.260 ;
        RECT 1688.270 1256.200 1688.590 1256.260 ;
        RECT 1684.590 1256.060 1688.590 1256.200 ;
        RECT 1684.590 1256.000 1684.910 1256.060 ;
        RECT 1688.270 1256.000 1688.590 1256.060 ;
        RECT 1683.210 1159.300 1683.530 1159.360 ;
        RECT 1684.590 1159.300 1684.910 1159.360 ;
        RECT 1683.210 1159.160 1684.910 1159.300 ;
        RECT 1683.210 1159.100 1683.530 1159.160 ;
        RECT 1684.590 1159.100 1684.910 1159.160 ;
        RECT 1683.210 1062.740 1683.530 1062.800 ;
        RECT 1684.590 1062.740 1684.910 1062.800 ;
        RECT 1683.210 1062.600 1684.910 1062.740 ;
        RECT 1683.210 1062.540 1683.530 1062.600 ;
        RECT 1684.590 1062.540 1684.910 1062.600 ;
        RECT 1683.210 966.180 1683.530 966.240 ;
        RECT 1684.590 966.180 1684.910 966.240 ;
        RECT 1683.210 966.040 1684.910 966.180 ;
        RECT 1683.210 965.980 1683.530 966.040 ;
        RECT 1684.590 965.980 1684.910 966.040 ;
        RECT 1684.130 717.640 1684.450 717.700 ;
        RECT 1684.590 717.640 1684.910 717.700 ;
        RECT 1684.130 717.500 1684.910 717.640 ;
        RECT 1684.130 717.440 1684.450 717.500 ;
        RECT 1684.590 717.440 1684.910 717.500 ;
        RECT 1684.145 386.140 1684.435 386.185 ;
        RECT 1684.590 386.140 1684.910 386.200 ;
        RECT 1684.145 386.000 1684.910 386.140 ;
        RECT 1684.145 385.955 1684.435 386.000 ;
        RECT 1684.590 385.940 1684.910 386.000 ;
        RECT 1684.130 338.200 1684.450 338.260 ;
        RECT 1683.935 338.060 1684.450 338.200 ;
        RECT 1684.130 338.000 1684.450 338.060 ;
        RECT 1683.670 303.520 1683.990 303.580 ;
        RECT 1684.590 303.520 1684.910 303.580 ;
        RECT 1683.670 303.380 1684.910 303.520 ;
        RECT 1683.670 303.320 1683.990 303.380 ;
        RECT 1684.590 303.320 1684.910 303.380 ;
        RECT 1684.145 289.580 1684.435 289.625 ;
        RECT 1684.590 289.580 1684.910 289.640 ;
        RECT 1684.145 289.440 1684.910 289.580 ;
        RECT 1684.145 289.395 1684.435 289.440 ;
        RECT 1684.590 289.380 1684.910 289.440 ;
        RECT 1684.130 241.640 1684.450 241.700 ;
        RECT 1683.935 241.500 1684.450 241.640 ;
        RECT 1684.130 241.440 1684.450 241.500 ;
        RECT 1683.670 206.960 1683.990 207.020 ;
        RECT 1684.590 206.960 1684.910 207.020 ;
        RECT 1683.670 206.820 1684.910 206.960 ;
        RECT 1683.670 206.760 1683.990 206.820 ;
        RECT 1684.590 206.760 1684.910 206.820 ;
        RECT 1683.685 179.420 1683.975 179.465 ;
        RECT 1684.590 179.420 1684.910 179.480 ;
        RECT 1683.685 179.280 1684.910 179.420 ;
        RECT 1683.685 179.235 1683.975 179.280 ;
        RECT 1684.590 179.220 1684.910 179.280 ;
        RECT 1683.670 131.820 1683.990 131.880 ;
        RECT 1683.475 131.680 1683.990 131.820 ;
        RECT 1683.670 131.620 1683.990 131.680 ;
        RECT 1683.670 131.140 1683.990 131.200 ;
        RECT 1684.130 131.140 1684.450 131.200 ;
        RECT 1683.670 131.000 1684.450 131.140 ;
        RECT 1683.670 130.940 1683.990 131.000 ;
        RECT 1684.130 130.940 1684.450 131.000 ;
        RECT 1684.130 82.860 1684.450 82.920 ;
        RECT 1683.935 82.720 1684.450 82.860 ;
        RECT 1684.130 82.660 1684.450 82.720 ;
        RECT 1684.130 34.580 1684.450 34.640 ;
        RECT 1683.935 34.440 1684.450 34.580 ;
        RECT 1684.130 34.380 1684.450 34.440 ;
        RECT 1685.510 2.960 1685.830 3.020 ;
        RECT 1685.970 2.960 1686.290 3.020 ;
        RECT 1685.510 2.820 1686.290 2.960 ;
        RECT 1685.510 2.760 1685.830 2.820 ;
        RECT 1685.970 2.760 1686.290 2.820 ;
      LAYER via ;
        RECT 1684.620 1256.000 1684.880 1256.260 ;
        RECT 1688.300 1256.000 1688.560 1256.260 ;
        RECT 1683.240 1159.100 1683.500 1159.360 ;
        RECT 1684.620 1159.100 1684.880 1159.360 ;
        RECT 1683.240 1062.540 1683.500 1062.800 ;
        RECT 1684.620 1062.540 1684.880 1062.800 ;
        RECT 1683.240 965.980 1683.500 966.240 ;
        RECT 1684.620 965.980 1684.880 966.240 ;
        RECT 1684.160 717.440 1684.420 717.700 ;
        RECT 1684.620 717.440 1684.880 717.700 ;
        RECT 1684.620 385.940 1684.880 386.200 ;
        RECT 1684.160 338.000 1684.420 338.260 ;
        RECT 1683.700 303.320 1683.960 303.580 ;
        RECT 1684.620 303.320 1684.880 303.580 ;
        RECT 1684.620 289.380 1684.880 289.640 ;
        RECT 1684.160 241.440 1684.420 241.700 ;
        RECT 1683.700 206.760 1683.960 207.020 ;
        RECT 1684.620 206.760 1684.880 207.020 ;
        RECT 1684.620 179.220 1684.880 179.480 ;
        RECT 1683.700 131.620 1683.960 131.880 ;
        RECT 1683.700 130.940 1683.960 131.200 ;
        RECT 1684.160 130.940 1684.420 131.200 ;
        RECT 1684.160 82.660 1684.420 82.920 ;
        RECT 1684.160 34.380 1684.420 34.640 ;
        RECT 1685.540 2.760 1685.800 3.020 ;
        RECT 1686.000 2.760 1686.260 3.020 ;
      LAYER met2 ;
        RECT 1690.180 1323.690 1690.460 1327.135 ;
        RECT 1688.360 1323.550 1690.460 1323.690 ;
        RECT 1688.360 1256.290 1688.500 1323.550 ;
        RECT 1690.180 1323.135 1690.460 1323.550 ;
        RECT 1684.620 1255.970 1684.880 1256.290 ;
        RECT 1688.300 1255.970 1688.560 1256.290 ;
        RECT 1684.680 1221.010 1684.820 1255.970 ;
        RECT 1684.220 1220.870 1684.820 1221.010 ;
        RECT 1684.220 1207.525 1684.360 1220.870 ;
        RECT 1683.230 1207.155 1683.510 1207.525 ;
        RECT 1684.150 1207.155 1684.430 1207.525 ;
        RECT 1683.300 1159.390 1683.440 1207.155 ;
        RECT 1683.240 1159.070 1683.500 1159.390 ;
        RECT 1684.620 1159.070 1684.880 1159.390 ;
        RECT 1684.680 1124.450 1684.820 1159.070 ;
        RECT 1684.220 1124.310 1684.820 1124.450 ;
        RECT 1684.220 1110.965 1684.360 1124.310 ;
        RECT 1683.230 1110.595 1683.510 1110.965 ;
        RECT 1684.150 1110.595 1684.430 1110.965 ;
        RECT 1683.300 1062.830 1683.440 1110.595 ;
        RECT 1683.240 1062.510 1683.500 1062.830 ;
        RECT 1684.620 1062.510 1684.880 1062.830 ;
        RECT 1684.680 1027.890 1684.820 1062.510 ;
        RECT 1684.220 1027.750 1684.820 1027.890 ;
        RECT 1684.220 1014.405 1684.360 1027.750 ;
        RECT 1683.230 1014.035 1683.510 1014.405 ;
        RECT 1684.150 1014.035 1684.430 1014.405 ;
        RECT 1683.300 966.270 1683.440 1014.035 ;
        RECT 1683.240 965.950 1683.500 966.270 ;
        RECT 1684.620 965.950 1684.880 966.270 ;
        RECT 1684.680 931.330 1684.820 965.950 ;
        RECT 1684.220 931.190 1684.820 931.330 ;
        RECT 1684.220 917.730 1684.360 931.190 ;
        RECT 1684.220 917.590 1684.820 917.730 ;
        RECT 1684.680 834.770 1684.820 917.590 ;
        RECT 1684.220 834.630 1684.820 834.770 ;
        RECT 1684.220 796.690 1684.360 834.630 ;
        RECT 1684.220 796.550 1684.820 796.690 ;
        RECT 1684.680 738.210 1684.820 796.550 ;
        RECT 1684.220 738.070 1684.820 738.210 ;
        RECT 1684.220 717.730 1684.360 738.070 ;
        RECT 1684.160 717.410 1684.420 717.730 ;
        RECT 1684.620 717.410 1684.880 717.730 ;
        RECT 1684.680 651.850 1684.820 717.410 ;
        RECT 1684.220 651.710 1684.820 651.850 ;
        RECT 1684.220 603.570 1684.360 651.710 ;
        RECT 1683.300 603.430 1684.360 603.570 ;
        RECT 1683.300 579.885 1683.440 603.430 ;
        RECT 1683.230 579.515 1683.510 579.885 ;
        RECT 1684.610 579.515 1684.890 579.885 ;
        RECT 1684.680 545.090 1684.820 579.515 ;
        RECT 1684.220 544.950 1684.820 545.090 ;
        RECT 1684.220 507.010 1684.360 544.950 ;
        RECT 1683.300 506.870 1684.360 507.010 ;
        RECT 1683.300 483.325 1683.440 506.870 ;
        RECT 1683.230 482.955 1683.510 483.325 ;
        RECT 1684.610 482.955 1684.890 483.325 ;
        RECT 1684.680 448.530 1684.820 482.955 ;
        RECT 1684.220 448.390 1684.820 448.530 ;
        RECT 1684.220 410.450 1684.360 448.390 ;
        RECT 1684.220 410.310 1685.280 410.450 ;
        RECT 1685.140 386.650 1685.280 410.310 ;
        RECT 1684.680 386.510 1685.280 386.650 ;
        RECT 1684.680 386.230 1684.820 386.510 ;
        RECT 1684.620 385.910 1684.880 386.230 ;
        RECT 1684.160 337.970 1684.420 338.290 ;
        RECT 1684.220 303.690 1684.360 337.970 ;
        RECT 1683.760 303.610 1684.360 303.690 ;
        RECT 1683.700 303.550 1684.360 303.610 ;
        RECT 1683.700 303.290 1683.960 303.550 ;
        RECT 1684.620 303.290 1684.880 303.610 ;
        RECT 1684.680 289.670 1684.820 303.290 ;
        RECT 1684.620 289.350 1684.880 289.670 ;
        RECT 1684.160 241.410 1684.420 241.730 ;
        RECT 1684.220 207.130 1684.360 241.410 ;
        RECT 1683.760 207.050 1684.360 207.130 ;
        RECT 1683.700 206.990 1684.360 207.050 ;
        RECT 1683.700 206.730 1683.960 206.990 ;
        RECT 1684.620 206.730 1684.880 207.050 ;
        RECT 1684.680 179.510 1684.820 206.730 ;
        RECT 1684.620 179.190 1684.880 179.510 ;
        RECT 1683.700 131.590 1683.960 131.910 ;
        RECT 1683.760 131.230 1683.900 131.590 ;
        RECT 1683.700 130.910 1683.960 131.230 ;
        RECT 1684.160 130.910 1684.420 131.230 ;
        RECT 1684.220 82.950 1684.360 130.910 ;
        RECT 1684.160 82.630 1684.420 82.950 ;
        RECT 1684.160 34.525 1684.420 34.670 ;
        RECT 1684.150 34.155 1684.430 34.525 ;
        RECT 1685.990 34.155 1686.270 34.525 ;
        RECT 1686.060 3.050 1686.200 34.155 ;
        RECT 1685.540 2.730 1685.800 3.050 ;
        RECT 1686.000 2.730 1686.260 3.050 ;
        RECT 1685.600 2.400 1685.740 2.730 ;
        RECT 1685.390 -4.800 1685.950 2.400 ;
      LAYER via2 ;
        RECT 1683.230 1207.200 1683.510 1207.480 ;
        RECT 1684.150 1207.200 1684.430 1207.480 ;
        RECT 1683.230 1110.640 1683.510 1110.920 ;
        RECT 1684.150 1110.640 1684.430 1110.920 ;
        RECT 1683.230 1014.080 1683.510 1014.360 ;
        RECT 1684.150 1014.080 1684.430 1014.360 ;
        RECT 1683.230 579.560 1683.510 579.840 ;
        RECT 1684.610 579.560 1684.890 579.840 ;
        RECT 1683.230 483.000 1683.510 483.280 ;
        RECT 1684.610 483.000 1684.890 483.280 ;
        RECT 1684.150 34.200 1684.430 34.480 ;
        RECT 1685.990 34.200 1686.270 34.480 ;
      LAYER met3 ;
        RECT 1683.205 1207.490 1683.535 1207.505 ;
        RECT 1684.125 1207.490 1684.455 1207.505 ;
        RECT 1683.205 1207.190 1684.455 1207.490 ;
        RECT 1683.205 1207.175 1683.535 1207.190 ;
        RECT 1684.125 1207.175 1684.455 1207.190 ;
        RECT 1683.205 1110.930 1683.535 1110.945 ;
        RECT 1684.125 1110.930 1684.455 1110.945 ;
        RECT 1683.205 1110.630 1684.455 1110.930 ;
        RECT 1683.205 1110.615 1683.535 1110.630 ;
        RECT 1684.125 1110.615 1684.455 1110.630 ;
        RECT 1683.205 1014.370 1683.535 1014.385 ;
        RECT 1684.125 1014.370 1684.455 1014.385 ;
        RECT 1683.205 1014.070 1684.455 1014.370 ;
        RECT 1683.205 1014.055 1683.535 1014.070 ;
        RECT 1684.125 1014.055 1684.455 1014.070 ;
        RECT 1683.205 579.850 1683.535 579.865 ;
        RECT 1684.585 579.850 1684.915 579.865 ;
        RECT 1683.205 579.550 1684.915 579.850 ;
        RECT 1683.205 579.535 1683.535 579.550 ;
        RECT 1684.585 579.535 1684.915 579.550 ;
        RECT 1683.205 483.290 1683.535 483.305 ;
        RECT 1684.585 483.290 1684.915 483.305 ;
        RECT 1683.205 482.990 1684.915 483.290 ;
        RECT 1683.205 482.975 1683.535 482.990 ;
        RECT 1684.585 482.975 1684.915 482.990 ;
        RECT 1684.125 34.490 1684.455 34.505 ;
        RECT 1685.965 34.490 1686.295 34.505 ;
        RECT 1684.125 34.190 1686.295 34.490 ;
        RECT 1684.125 34.175 1684.455 34.190 ;
        RECT 1685.965 34.175 1686.295 34.190 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 722.270 53.280 722.590 53.340 ;
        RECT 1449.070 53.280 1449.390 53.340 ;
        RECT 722.270 53.140 1449.390 53.280 ;
        RECT 722.270 53.080 722.590 53.140 ;
        RECT 1449.070 53.080 1449.390 53.140 ;
      LAYER via ;
        RECT 722.300 53.080 722.560 53.340 ;
        RECT 1449.100 53.080 1449.360 53.340 ;
      LAYER met2 ;
        RECT 1452.820 1323.690 1453.100 1327.135 ;
        RECT 1449.160 1323.550 1453.100 1323.690 ;
        RECT 1449.160 53.370 1449.300 1323.550 ;
        RECT 1452.820 1323.135 1453.100 1323.550 ;
        RECT 722.300 53.050 722.560 53.370 ;
        RECT 1449.100 53.050 1449.360 53.370 ;
        RECT 722.360 2.400 722.500 53.050 ;
        RECT 722.150 -4.800 722.710 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 704.865 1518.865 705.035 1597.575 ;
        RECT 704.865 1308.065 705.035 1393.575 ;
      LAYER mcon ;
        RECT 704.865 1597.405 705.035 1597.575 ;
        RECT 704.865 1393.405 705.035 1393.575 ;
      LAYER met1 ;
        RECT 704.790 1616.600 705.110 1616.660 ;
        RECT 712.150 1616.600 712.470 1616.660 ;
        RECT 704.790 1616.460 712.470 1616.600 ;
        RECT 704.790 1616.400 705.110 1616.460 ;
        RECT 712.150 1616.400 712.470 1616.460 ;
        RECT 704.790 1597.560 705.110 1597.620 ;
        RECT 704.595 1597.420 705.110 1597.560 ;
        RECT 704.790 1597.360 705.110 1597.420 ;
        RECT 704.790 1519.020 705.110 1519.080 ;
        RECT 704.595 1518.880 705.110 1519.020 ;
        RECT 704.790 1518.820 705.110 1518.880 ;
        RECT 704.790 1393.560 705.110 1393.620 ;
        RECT 704.595 1393.420 705.110 1393.560 ;
        RECT 704.790 1393.360 705.110 1393.420 ;
        RECT 704.805 1308.220 705.095 1308.265 ;
        RECT 1697.470 1308.220 1697.790 1308.280 ;
        RECT 704.805 1308.080 1697.790 1308.220 ;
        RECT 704.805 1308.035 705.095 1308.080 ;
        RECT 1697.470 1308.020 1697.790 1308.080 ;
        RECT 1697.470 37.980 1697.790 38.040 ;
        RECT 1703.450 37.980 1703.770 38.040 ;
        RECT 1697.470 37.840 1703.770 37.980 ;
        RECT 1697.470 37.780 1697.790 37.840 ;
        RECT 1703.450 37.780 1703.770 37.840 ;
      LAYER via ;
        RECT 704.820 1616.400 705.080 1616.660 ;
        RECT 712.180 1616.400 712.440 1616.660 ;
        RECT 704.820 1597.360 705.080 1597.620 ;
        RECT 704.820 1518.820 705.080 1519.080 ;
        RECT 704.820 1393.360 705.080 1393.620 ;
        RECT 1697.500 1308.020 1697.760 1308.280 ;
        RECT 1697.500 37.780 1697.760 38.040 ;
        RECT 1703.480 37.780 1703.740 38.040 ;
      LAYER met2 ;
        RECT 712.170 1660.715 712.450 1661.085 ;
        RECT 712.240 1616.690 712.380 1660.715 ;
        RECT 704.820 1616.370 705.080 1616.690 ;
        RECT 712.180 1616.370 712.440 1616.690 ;
        RECT 704.880 1597.650 705.020 1616.370 ;
        RECT 704.820 1597.330 705.080 1597.650 ;
        RECT 704.820 1518.790 705.080 1519.110 ;
        RECT 704.880 1393.650 705.020 1518.790 ;
        RECT 704.820 1393.330 705.080 1393.650 ;
        RECT 1697.500 1307.990 1697.760 1308.310 ;
        RECT 1697.560 38.070 1697.700 1307.990 ;
        RECT 1697.500 37.750 1697.760 38.070 ;
        RECT 1703.480 37.750 1703.740 38.070 ;
        RECT 1703.540 2.400 1703.680 37.750 ;
        RECT 1703.330 -4.800 1703.890 2.400 ;
      LAYER via2 ;
        RECT 712.170 1660.760 712.450 1661.040 ;
      LAYER met3 ;
        RECT 712.145 1661.050 712.475 1661.065 ;
        RECT 715.810 1661.050 719.810 1661.055 ;
        RECT 712.145 1660.750 719.810 1661.050 ;
        RECT 712.145 1660.735 712.475 1660.750 ;
        RECT 715.810 1660.455 719.810 1660.750 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1752.745 2377.535 1752.915 2378.895 ;
        RECT 1752.745 2377.365 1755.675 2377.535 ;
      LAYER mcon ;
        RECT 1752.745 2378.725 1752.915 2378.895 ;
        RECT 1755.505 2377.365 1755.675 2377.535 ;
      LAYER met1 ;
        RECT 1502.430 2378.880 1502.750 2378.940 ;
        RECT 1752.685 2378.880 1752.975 2378.925 ;
        RECT 1502.430 2378.740 1752.975 2378.880 ;
        RECT 1502.430 2378.680 1502.750 2378.740 ;
        RECT 1752.685 2378.695 1752.975 2378.740 ;
        RECT 1755.445 2377.520 1755.735 2377.565 ;
        RECT 1780.270 2377.520 1780.590 2377.580 ;
        RECT 1755.445 2377.380 1780.590 2377.520 ;
        RECT 1755.445 2377.335 1755.735 2377.380 ;
        RECT 1780.270 2377.320 1780.590 2377.380 ;
        RECT 1721.390 15.200 1721.710 15.260 ;
        RECT 1779.810 15.200 1780.130 15.260 ;
        RECT 1721.390 15.060 1780.130 15.200 ;
        RECT 1721.390 15.000 1721.710 15.060 ;
        RECT 1779.810 15.000 1780.130 15.060 ;
      LAYER via ;
        RECT 1502.460 2378.680 1502.720 2378.940 ;
        RECT 1780.300 2377.320 1780.560 2377.580 ;
        RECT 1721.420 15.000 1721.680 15.260 ;
        RECT 1779.840 15.000 1780.100 15.260 ;
      LAYER met2 ;
        RECT 1502.460 2378.650 1502.720 2378.970 ;
        RECT 1502.520 2377.880 1502.660 2378.650 ;
        RECT 1502.500 2373.880 1502.780 2377.880 ;
        RECT 1780.300 2377.290 1780.560 2377.610 ;
        RECT 1780.360 22.170 1780.500 2377.290 ;
        RECT 1779.900 22.030 1780.500 22.170 ;
        RECT 1779.900 15.290 1780.040 22.030 ;
        RECT 1721.420 14.970 1721.680 15.290 ;
        RECT 1779.840 14.970 1780.100 15.290 ;
        RECT 1721.480 2.400 1721.620 14.970 ;
        RECT 1721.270 -4.800 1721.830 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1745.310 1326.580 1745.630 1326.640 ;
        RECT 1756.810 1326.580 1757.130 1326.640 ;
        RECT 1745.310 1326.440 1757.130 1326.580 ;
        RECT 1745.310 1326.380 1745.630 1326.440 ;
        RECT 1756.810 1326.380 1757.130 1326.440 ;
        RECT 1739.330 20.300 1739.650 20.360 ;
        RECT 1745.310 20.300 1745.630 20.360 ;
        RECT 1739.330 20.160 1745.630 20.300 ;
        RECT 1739.330 20.100 1739.650 20.160 ;
        RECT 1745.310 20.100 1745.630 20.160 ;
      LAYER via ;
        RECT 1745.340 1326.380 1745.600 1326.640 ;
        RECT 1756.840 1326.380 1757.100 1326.640 ;
        RECT 1739.360 20.100 1739.620 20.360 ;
        RECT 1745.340 20.100 1745.600 20.360 ;
      LAYER met2 ;
        RECT 1756.830 1327.515 1757.110 1327.885 ;
        RECT 1756.900 1326.670 1757.040 1327.515 ;
        RECT 1745.340 1326.350 1745.600 1326.670 ;
        RECT 1756.840 1326.350 1757.100 1326.670 ;
        RECT 1745.400 20.390 1745.540 1326.350 ;
        RECT 1739.360 20.070 1739.620 20.390 ;
        RECT 1745.340 20.070 1745.600 20.390 ;
        RECT 1739.420 2.400 1739.560 20.070 ;
        RECT 1739.210 -4.800 1739.770 2.400 ;
      LAYER via2 ;
        RECT 1756.830 1327.560 1757.110 1327.840 ;
      LAYER met3 ;
        RECT 1755.835 1329.975 1759.835 1330.575 ;
        RECT 1756.590 1327.865 1756.890 1329.975 ;
        RECT 1756.590 1327.550 1757.135 1327.865 ;
        RECT 1756.805 1327.535 1757.135 1327.550 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 709.390 40.020 709.710 40.080 ;
        RECT 1756.810 40.020 1757.130 40.080 ;
        RECT 709.390 39.880 1757.130 40.020 ;
        RECT 709.390 39.820 709.710 39.880 ;
        RECT 1756.810 39.820 1757.130 39.880 ;
      LAYER via ;
        RECT 709.420 39.820 709.680 40.080 ;
        RECT 1756.840 39.820 1757.100 40.080 ;
      LAYER met2 ;
        RECT 709.410 1976.235 709.690 1976.605 ;
        RECT 709.480 40.110 709.620 1976.235 ;
        RECT 709.420 39.790 709.680 40.110 ;
        RECT 1756.840 39.790 1757.100 40.110 ;
        RECT 1756.900 2.400 1757.040 39.790 ;
        RECT 1756.690 -4.800 1757.250 2.400 ;
      LAYER via2 ;
        RECT 709.410 1976.280 709.690 1976.560 ;
      LAYER met3 ;
        RECT 709.385 1976.570 709.715 1976.585 ;
        RECT 715.810 1976.570 719.810 1976.575 ;
        RECT 709.385 1976.270 719.810 1976.570 ;
        RECT 709.385 1976.255 709.715 1976.270 ;
        RECT 715.810 1975.975 719.810 1976.270 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1774.825 2.805 1774.995 48.195 ;
      LAYER mcon ;
        RECT 1774.825 48.025 1774.995 48.195 ;
      LAYER met1 ;
        RECT 1773.370 2378.880 1773.690 2378.940 ;
        RECT 1753.220 2378.740 1773.690 2378.880 ;
        RECT 1472.990 2378.540 1473.310 2378.600 ;
        RECT 1753.220 2378.540 1753.360 2378.740 ;
        RECT 1773.370 2378.680 1773.690 2378.740 ;
        RECT 1472.990 2378.400 1753.360 2378.540 ;
        RECT 1472.990 2378.340 1473.310 2378.400 ;
        RECT 1773.370 61.440 1773.690 61.500 ;
        RECT 1776.130 61.440 1776.450 61.500 ;
        RECT 1773.370 61.300 1776.450 61.440 ;
        RECT 1773.370 61.240 1773.690 61.300 ;
        RECT 1776.130 61.240 1776.450 61.300 ;
        RECT 1774.765 48.180 1775.055 48.225 ;
        RECT 1776.130 48.180 1776.450 48.240 ;
        RECT 1774.765 48.040 1776.450 48.180 ;
        RECT 1774.765 47.995 1775.055 48.040 ;
        RECT 1776.130 47.980 1776.450 48.040 ;
        RECT 1774.750 2.960 1775.070 3.020 ;
        RECT 1774.555 2.820 1775.070 2.960 ;
        RECT 1774.750 2.760 1775.070 2.820 ;
      LAYER via ;
        RECT 1473.020 2378.340 1473.280 2378.600 ;
        RECT 1773.400 2378.680 1773.660 2378.940 ;
        RECT 1773.400 61.240 1773.660 61.500 ;
        RECT 1776.160 61.240 1776.420 61.500 ;
        RECT 1776.160 47.980 1776.420 48.240 ;
        RECT 1774.780 2.760 1775.040 3.020 ;
      LAYER met2 ;
        RECT 1773.400 2378.650 1773.660 2378.970 ;
        RECT 1473.020 2378.310 1473.280 2378.630 ;
        RECT 1473.080 2377.880 1473.220 2378.310 ;
        RECT 1473.060 2373.880 1473.340 2377.880 ;
        RECT 1773.460 61.530 1773.600 2378.650 ;
        RECT 1773.400 61.210 1773.660 61.530 ;
        RECT 1776.160 61.210 1776.420 61.530 ;
        RECT 1776.220 48.270 1776.360 61.210 ;
        RECT 1776.160 47.950 1776.420 48.270 ;
        RECT 1774.780 2.730 1775.040 3.050 ;
        RECT 1774.840 2.400 1774.980 2.730 ;
        RECT 1774.630 -4.800 1775.190 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1792.765 2.805 1792.935 25.415 ;
      LAYER mcon ;
        RECT 1792.765 25.245 1792.935 25.415 ;
      LAYER met1 ;
        RECT 716.750 1307.880 717.070 1307.940 ;
        RECT 1788.090 1307.880 1788.410 1307.940 ;
        RECT 716.750 1307.740 1788.410 1307.880 ;
        RECT 716.750 1307.680 717.070 1307.740 ;
        RECT 1788.090 1307.680 1788.410 1307.740 ;
        RECT 1788.090 25.400 1788.410 25.460 ;
        RECT 1792.705 25.400 1792.995 25.445 ;
        RECT 1788.090 25.260 1792.995 25.400 ;
        RECT 1788.090 25.200 1788.410 25.260 ;
        RECT 1792.705 25.215 1792.995 25.260 ;
        RECT 1792.690 2.960 1793.010 3.020 ;
        RECT 1792.495 2.820 1793.010 2.960 ;
        RECT 1792.690 2.760 1793.010 2.820 ;
      LAYER via ;
        RECT 716.780 1307.680 717.040 1307.940 ;
        RECT 1788.120 1307.680 1788.380 1307.940 ;
        RECT 1788.120 25.200 1788.380 25.460 ;
        RECT 1792.720 2.760 1792.980 3.020 ;
      LAYER met2 ;
        RECT 716.770 1444.475 717.050 1444.845 ;
        RECT 716.840 1307.970 716.980 1444.475 ;
        RECT 716.780 1307.650 717.040 1307.970 ;
        RECT 1788.120 1307.650 1788.380 1307.970 ;
        RECT 1788.180 25.490 1788.320 1307.650 ;
        RECT 1788.120 25.170 1788.380 25.490 ;
        RECT 1792.720 2.730 1792.980 3.050 ;
        RECT 1792.780 2.400 1792.920 2.730 ;
        RECT 1792.570 -4.800 1793.130 2.400 ;
      LAYER via2 ;
        RECT 716.770 1444.520 717.050 1444.800 ;
      LAYER met3 ;
        RECT 715.810 1446.935 719.810 1447.535 ;
        RECT 716.990 1444.825 717.290 1446.935 ;
        RECT 716.745 1444.510 717.290 1444.825 ;
        RECT 716.745 1444.495 717.075 1444.510 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1372.710 26.760 1373.030 26.820 ;
        RECT 1810.630 26.760 1810.950 26.820 ;
        RECT 1372.710 26.620 1810.950 26.760 ;
        RECT 1372.710 26.560 1373.030 26.620 ;
        RECT 1810.630 26.560 1810.950 26.620 ;
      LAYER via ;
        RECT 1372.740 26.560 1373.000 26.820 ;
        RECT 1810.660 26.560 1810.920 26.820 ;
      LAYER met2 ;
        RECT 1371.860 1323.690 1372.140 1327.135 ;
        RECT 1371.860 1323.550 1372.940 1323.690 ;
        RECT 1371.860 1323.135 1372.140 1323.550 ;
        RECT 1372.800 26.850 1372.940 1323.550 ;
        RECT 1372.740 26.530 1373.000 26.850 ;
        RECT 1810.660 26.530 1810.920 26.850 ;
        RECT 1810.720 2.400 1810.860 26.530 ;
        RECT 1810.510 -4.800 1811.070 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1772.910 1718.260 1773.230 1718.320 ;
        RECT 1829.030 1718.260 1829.350 1718.320 ;
        RECT 1772.910 1718.120 1829.350 1718.260 ;
        RECT 1772.910 1718.060 1773.230 1718.120 ;
        RECT 1829.030 1718.060 1829.350 1718.120 ;
      LAYER via ;
        RECT 1772.940 1718.060 1773.200 1718.320 ;
        RECT 1829.060 1718.060 1829.320 1718.320 ;
      LAYER met2 ;
        RECT 1772.930 1724.635 1773.210 1725.005 ;
        RECT 1773.000 1718.350 1773.140 1724.635 ;
        RECT 1772.940 1718.030 1773.200 1718.350 ;
        RECT 1829.060 1718.030 1829.320 1718.350 ;
        RECT 1829.120 17.410 1829.260 1718.030 ;
        RECT 1828.660 17.270 1829.260 17.410 ;
        RECT 1828.660 2.400 1828.800 17.270 ;
        RECT 1828.450 -4.800 1829.010 2.400 ;
      LAYER via2 ;
        RECT 1772.930 1724.680 1773.210 1724.960 ;
      LAYER met3 ;
        RECT 1755.835 1724.970 1759.835 1724.975 ;
        RECT 1772.905 1724.970 1773.235 1724.985 ;
        RECT 1755.835 1724.670 1773.235 1724.970 ;
        RECT 1755.835 1724.375 1759.835 1724.670 ;
        RECT 1772.905 1724.655 1773.235 1724.670 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 728.270 1307.795 728.550 1308.165 ;
        RECT 728.340 19.565 728.480 1307.795 ;
        RECT 728.270 19.195 728.550 19.565 ;
        RECT 1846.070 19.195 1846.350 19.565 ;
        RECT 1846.140 2.400 1846.280 19.195 ;
        RECT 1845.930 -4.800 1846.490 2.400 ;
      LAYER via2 ;
        RECT 728.270 1307.840 728.550 1308.120 ;
        RECT 728.270 19.240 728.550 19.520 ;
        RECT 1846.070 19.240 1846.350 19.520 ;
      LAYER met3 ;
        RECT 707.750 2345.130 708.130 2345.140 ;
        RECT 715.810 2345.130 719.810 2345.135 ;
        RECT 707.750 2344.830 719.810 2345.130 ;
        RECT 707.750 2344.820 708.130 2344.830 ;
        RECT 715.810 2344.535 719.810 2344.830 ;
        RECT 707.750 1308.130 708.130 1308.140 ;
        RECT 728.245 1308.130 728.575 1308.145 ;
        RECT 707.750 1307.830 728.575 1308.130 ;
        RECT 707.750 1307.820 708.130 1307.830 ;
        RECT 728.245 1307.815 728.575 1307.830 ;
        RECT 728.245 19.530 728.575 19.545 ;
        RECT 1846.045 19.530 1846.375 19.545 ;
        RECT 728.245 19.230 1846.375 19.530 ;
        RECT 728.245 19.215 728.575 19.230 ;
        RECT 1846.045 19.215 1846.375 19.230 ;
      LAYER via3 ;
        RECT 707.780 2344.820 708.100 2345.140 ;
        RECT 707.780 1307.820 708.100 1308.140 ;
      LAYER met4 ;
        RECT 707.775 2344.815 708.105 2345.145 ;
        RECT 707.790 1308.145 708.090 2344.815 ;
        RECT 707.775 1307.815 708.105 1308.145 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1864.065 2.805 1864.235 16.235 ;
      LAYER mcon ;
        RECT 1864.065 16.065 1864.235 16.235 ;
      LAYER met1 ;
        RECT 1863.070 1307.540 1863.390 1307.600 ;
        RECT 720.520 1307.400 1863.390 1307.540 ;
        RECT 715.370 1307.200 715.690 1307.260 ;
        RECT 720.520 1307.200 720.660 1307.400 ;
        RECT 1863.070 1307.340 1863.390 1307.400 ;
        RECT 715.370 1307.060 720.660 1307.200 ;
        RECT 715.370 1307.000 715.690 1307.060 ;
        RECT 1863.070 16.220 1863.390 16.280 ;
        RECT 1864.005 16.220 1864.295 16.265 ;
        RECT 1863.070 16.080 1864.295 16.220 ;
        RECT 1863.070 16.020 1863.390 16.080 ;
        RECT 1864.005 16.035 1864.295 16.080 ;
        RECT 1863.990 2.960 1864.310 3.020 ;
        RECT 1863.795 2.820 1864.310 2.960 ;
        RECT 1863.990 2.760 1864.310 2.820 ;
      LAYER via ;
        RECT 715.400 1307.000 715.660 1307.260 ;
        RECT 1863.100 1307.340 1863.360 1307.600 ;
        RECT 1863.100 16.020 1863.360 16.280 ;
        RECT 1864.020 2.760 1864.280 3.020 ;
      LAYER met2 ;
        RECT 715.390 2140.115 715.670 2140.485 ;
        RECT 715.460 1307.290 715.600 2140.115 ;
        RECT 1863.100 1307.310 1863.360 1307.630 ;
        RECT 715.400 1306.970 715.660 1307.290 ;
        RECT 1863.160 16.310 1863.300 1307.310 ;
        RECT 1863.100 15.990 1863.360 16.310 ;
        RECT 1864.020 2.730 1864.280 3.050 ;
        RECT 1864.080 2.400 1864.220 2.730 ;
        RECT 1863.870 -4.800 1864.430 2.400 ;
      LAYER via2 ;
        RECT 715.390 2140.160 715.670 2140.440 ;
      LAYER met3 ;
        RECT 715.365 2140.450 715.695 2140.465 ;
        RECT 715.365 2140.150 716.370 2140.450 ;
        RECT 715.365 2140.135 715.695 2140.150 ;
        RECT 716.070 2139.775 716.370 2140.150 ;
        RECT 715.810 2139.175 719.810 2139.775 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1757.270 2028.000 1757.590 2028.060 ;
        RECT 1758.190 2028.000 1758.510 2028.060 ;
        RECT 1757.270 2027.860 1758.510 2028.000 ;
        RECT 1757.270 2027.800 1757.590 2027.860 ;
        RECT 1758.190 2027.800 1758.510 2027.860 ;
        RECT 1758.190 1774.360 1758.510 1774.420 ;
        RECT 1759.110 1774.360 1759.430 1774.420 ;
        RECT 1758.190 1774.220 1759.430 1774.360 ;
        RECT 1758.190 1774.160 1758.510 1774.220 ;
        RECT 1759.110 1774.160 1759.430 1774.220 ;
        RECT 740.210 18.260 740.530 18.320 ;
        RECT 744.810 18.260 745.130 18.320 ;
        RECT 740.210 18.120 745.130 18.260 ;
        RECT 740.210 18.060 740.530 18.120 ;
        RECT 744.810 18.060 745.130 18.120 ;
      LAYER via ;
        RECT 1757.300 2027.800 1757.560 2028.060 ;
        RECT 1758.220 2027.800 1758.480 2028.060 ;
        RECT 1758.220 1774.160 1758.480 1774.420 ;
        RECT 1759.140 1774.160 1759.400 1774.420 ;
        RECT 740.240 18.060 740.500 18.320 ;
        RECT 744.840 18.060 745.100 18.320 ;
      LAYER met2 ;
        RECT 1758.670 2354.315 1758.950 2354.685 ;
        RECT 1758.740 2318.645 1758.880 2354.315 ;
        RECT 1758.670 2318.275 1758.950 2318.645 ;
        RECT 1756.830 2307.395 1757.110 2307.765 ;
        RECT 1756.900 2283.285 1757.040 2307.395 ;
        RECT 1756.830 2282.915 1757.110 2283.285 ;
        RECT 1757.290 2097.275 1757.570 2097.645 ;
        RECT 1757.360 2054.805 1757.500 2097.275 ;
        RECT 1757.290 2054.435 1757.570 2054.805 ;
        RECT 1757.290 2042.875 1757.570 2043.245 ;
        RECT 1757.360 2028.090 1757.500 2042.875 ;
        RECT 1757.300 2027.770 1757.560 2028.090 ;
        RECT 1758.220 2027.770 1758.480 2028.090 ;
        RECT 1758.280 1997.005 1758.420 2027.770 ;
        RECT 1758.210 1996.635 1758.490 1997.005 ;
        RECT 1757.290 1964.675 1757.570 1965.045 ;
        RECT 1757.360 1867.805 1757.500 1964.675 ;
        RECT 1757.290 1867.435 1757.570 1867.805 ;
        RECT 1758.210 1840.915 1758.490 1841.285 ;
        RECT 1758.280 1774.450 1758.420 1840.915 ;
        RECT 1758.220 1774.130 1758.480 1774.450 ;
        RECT 1759.140 1774.130 1759.400 1774.450 ;
        RECT 1759.200 1746.085 1759.340 1774.130 ;
        RECT 1759.130 1745.715 1759.410 1746.085 ;
        RECT 1757.750 1665.475 1758.030 1665.845 ;
        RECT 1757.820 1663.805 1757.960 1665.475 ;
        RECT 1757.750 1663.435 1758.030 1663.805 ;
        RECT 1758.210 1608.355 1758.490 1608.725 ;
        RECT 1758.280 1602.605 1758.420 1608.355 ;
        RECT 1758.210 1602.235 1758.490 1602.605 ;
        RECT 1765.570 1556.675 1765.850 1557.045 ;
        RECT 1765.640 1513.525 1765.780 1556.675 ;
        RECT 1765.570 1513.155 1765.850 1513.525 ;
        RECT 744.830 1302.355 745.110 1302.725 ;
        RECT 744.900 18.350 745.040 1302.355 ;
        RECT 740.240 18.030 740.500 18.350 ;
        RECT 744.840 18.030 745.100 18.350 ;
        RECT 740.300 2.400 740.440 18.030 ;
        RECT 740.090 -4.800 740.650 2.400 ;
      LAYER via2 ;
        RECT 1758.670 2354.360 1758.950 2354.640 ;
        RECT 1758.670 2318.320 1758.950 2318.600 ;
        RECT 1756.830 2307.440 1757.110 2307.720 ;
        RECT 1756.830 2282.960 1757.110 2283.240 ;
        RECT 1757.290 2097.320 1757.570 2097.600 ;
        RECT 1757.290 2054.480 1757.570 2054.760 ;
        RECT 1757.290 2042.920 1757.570 2043.200 ;
        RECT 1758.210 1996.680 1758.490 1996.960 ;
        RECT 1757.290 1964.720 1757.570 1965.000 ;
        RECT 1757.290 1867.480 1757.570 1867.760 ;
        RECT 1758.210 1840.960 1758.490 1841.240 ;
        RECT 1759.130 1745.760 1759.410 1746.040 ;
        RECT 1757.750 1665.520 1758.030 1665.800 ;
        RECT 1757.750 1663.480 1758.030 1663.760 ;
        RECT 1758.210 1608.400 1758.490 1608.680 ;
        RECT 1758.210 1602.280 1758.490 1602.560 ;
        RECT 1765.570 1556.720 1765.850 1557.000 ;
        RECT 1765.570 1513.200 1765.850 1513.480 ;
        RECT 744.830 1302.400 745.110 1302.680 ;
      LAYER met3 ;
        RECT 1755.835 2356.775 1759.835 2357.375 ;
        RECT 1758.430 2354.665 1758.730 2356.775 ;
        RECT 1758.430 2354.350 1758.975 2354.665 ;
        RECT 1758.645 2354.335 1758.975 2354.350 ;
        RECT 1756.550 2318.610 1756.930 2318.620 ;
        RECT 1758.645 2318.610 1758.975 2318.625 ;
        RECT 1756.550 2318.310 1758.975 2318.610 ;
        RECT 1756.550 2318.300 1756.930 2318.310 ;
        RECT 1758.645 2318.295 1758.975 2318.310 ;
        RECT 1756.550 2309.090 1756.930 2309.100 ;
        RECT 1756.550 2308.780 1757.120 2309.090 ;
        RECT 1756.820 2307.745 1757.120 2308.780 ;
        RECT 1756.805 2307.415 1757.135 2307.745 ;
        RECT 1756.805 2283.260 1757.135 2283.265 ;
        RECT 1756.550 2283.250 1757.135 2283.260 ;
        RECT 1756.350 2282.950 1757.135 2283.250 ;
        RECT 1756.550 2282.940 1757.135 2282.950 ;
        RECT 1756.805 2282.935 1757.135 2282.940 ;
        RECT 1756.550 2188.420 1756.930 2188.740 ;
        RECT 1756.590 2186.700 1756.890 2188.420 ;
        RECT 1756.550 2186.380 1756.930 2186.700 ;
        RECT 1757.265 2097.610 1757.595 2097.625 ;
        RECT 1758.390 2097.610 1758.770 2097.620 ;
        RECT 1757.265 2097.310 1758.770 2097.610 ;
        RECT 1757.265 2097.295 1757.595 2097.310 ;
        RECT 1758.390 2097.300 1758.770 2097.310 ;
        RECT 1756.550 2054.770 1756.930 2054.780 ;
        RECT 1757.265 2054.770 1757.595 2054.785 ;
        RECT 1756.550 2054.470 1757.595 2054.770 ;
        RECT 1756.550 2054.460 1756.930 2054.470 ;
        RECT 1757.265 2054.455 1757.595 2054.470 ;
        RECT 1756.550 2043.210 1756.930 2043.220 ;
        RECT 1757.265 2043.210 1757.595 2043.225 ;
        RECT 1756.550 2042.910 1757.595 2043.210 ;
        RECT 1756.550 2042.900 1756.930 2042.910 ;
        RECT 1757.265 2042.895 1757.595 2042.910 ;
        RECT 1756.550 1996.970 1756.930 1996.980 ;
        RECT 1758.185 1996.970 1758.515 1996.985 ;
        RECT 1756.550 1996.670 1758.515 1996.970 ;
        RECT 1756.550 1996.660 1756.930 1996.670 ;
        RECT 1758.185 1996.655 1758.515 1996.670 ;
        RECT 1756.550 1965.010 1756.930 1965.020 ;
        RECT 1757.265 1965.010 1757.595 1965.025 ;
        RECT 1756.550 1964.710 1757.595 1965.010 ;
        RECT 1756.550 1964.700 1756.930 1964.710 ;
        RECT 1757.265 1964.695 1757.595 1964.710 ;
        RECT 1756.550 1867.770 1756.930 1867.780 ;
        RECT 1757.265 1867.770 1757.595 1867.785 ;
        RECT 1756.550 1867.470 1757.595 1867.770 ;
        RECT 1756.550 1867.460 1756.930 1867.470 ;
        RECT 1757.265 1867.455 1757.595 1867.470 ;
        RECT 1756.550 1841.620 1756.930 1841.940 ;
        RECT 1756.590 1841.250 1756.890 1841.620 ;
        RECT 1758.185 1841.250 1758.515 1841.265 ;
        RECT 1756.590 1840.950 1758.515 1841.250 ;
        RECT 1758.185 1840.935 1758.515 1840.950 ;
        RECT 1756.550 1746.050 1756.930 1746.060 ;
        RECT 1759.105 1746.050 1759.435 1746.065 ;
        RECT 1756.550 1745.750 1759.435 1746.050 ;
        RECT 1756.550 1745.740 1756.930 1745.750 ;
        RECT 1759.105 1745.735 1759.435 1745.750 ;
        RECT 1757.470 1705.930 1757.850 1705.940 ;
        RECT 1756.590 1705.630 1757.850 1705.930 ;
        RECT 1756.590 1704.580 1756.890 1705.630 ;
        RECT 1757.470 1705.620 1757.850 1705.630 ;
        RECT 1756.550 1704.260 1756.930 1704.580 ;
        RECT 1756.550 1665.810 1756.930 1665.820 ;
        RECT 1757.725 1665.810 1758.055 1665.825 ;
        RECT 1756.550 1665.510 1758.055 1665.810 ;
        RECT 1756.550 1665.500 1756.930 1665.510 ;
        RECT 1757.725 1665.495 1758.055 1665.510 ;
        RECT 1756.550 1663.770 1756.930 1663.780 ;
        RECT 1757.725 1663.770 1758.055 1663.785 ;
        RECT 1756.550 1663.470 1758.055 1663.770 ;
        RECT 1756.550 1663.460 1756.930 1663.470 ;
        RECT 1757.725 1663.455 1758.055 1663.470 ;
        RECT 1756.550 1608.690 1756.930 1608.700 ;
        RECT 1758.185 1608.690 1758.515 1608.705 ;
        RECT 1756.550 1608.390 1758.515 1608.690 ;
        RECT 1756.550 1608.380 1756.930 1608.390 ;
        RECT 1758.185 1608.375 1758.515 1608.390 ;
        RECT 1756.550 1602.570 1756.930 1602.580 ;
        RECT 1758.185 1602.570 1758.515 1602.585 ;
        RECT 1756.550 1602.270 1758.515 1602.570 ;
        RECT 1756.550 1602.260 1756.930 1602.270 ;
        RECT 1758.185 1602.255 1758.515 1602.270 ;
        RECT 1756.550 1557.010 1756.930 1557.020 ;
        RECT 1765.545 1557.010 1765.875 1557.025 ;
        RECT 1756.550 1556.710 1765.875 1557.010 ;
        RECT 1756.550 1556.700 1756.930 1556.710 ;
        RECT 1765.545 1556.695 1765.875 1556.710 ;
        RECT 1756.550 1513.490 1756.930 1513.500 ;
        RECT 1765.545 1513.490 1765.875 1513.505 ;
        RECT 1756.550 1513.190 1765.875 1513.490 ;
        RECT 1756.550 1513.180 1756.930 1513.190 ;
        RECT 1765.545 1513.175 1765.875 1513.190 ;
        RECT 1756.550 1413.530 1756.930 1413.540 ;
        RECT 1764.830 1413.530 1765.210 1413.540 ;
        RECT 1756.550 1413.230 1765.210 1413.530 ;
        RECT 1756.550 1413.220 1756.930 1413.230 ;
        RECT 1764.830 1413.220 1765.210 1413.230 ;
        RECT 1756.550 1361.170 1756.930 1361.180 ;
        RECT 1764.830 1361.170 1765.210 1361.180 ;
        RECT 1756.550 1360.870 1765.210 1361.170 ;
        RECT 1756.550 1360.860 1756.930 1360.870 ;
        RECT 1764.830 1360.860 1765.210 1360.870 ;
        RECT 744.805 1302.690 745.135 1302.705 ;
        RECT 1756.550 1302.690 1756.930 1302.700 ;
        RECT 744.805 1302.390 1756.930 1302.690 ;
        RECT 744.805 1302.375 745.135 1302.390 ;
        RECT 1756.550 1302.380 1756.930 1302.390 ;
      LAYER via3 ;
        RECT 1756.580 2318.300 1756.900 2318.620 ;
        RECT 1756.580 2308.780 1756.900 2309.100 ;
        RECT 1756.580 2282.940 1756.900 2283.260 ;
        RECT 1756.580 2188.420 1756.900 2188.740 ;
        RECT 1756.580 2186.380 1756.900 2186.700 ;
        RECT 1758.420 2097.300 1758.740 2097.620 ;
        RECT 1756.580 2054.460 1756.900 2054.780 ;
        RECT 1756.580 2042.900 1756.900 2043.220 ;
        RECT 1756.580 1996.660 1756.900 1996.980 ;
        RECT 1756.580 1964.700 1756.900 1965.020 ;
        RECT 1756.580 1867.460 1756.900 1867.780 ;
        RECT 1756.580 1841.620 1756.900 1841.940 ;
        RECT 1756.580 1745.740 1756.900 1746.060 ;
        RECT 1757.500 1705.620 1757.820 1705.940 ;
        RECT 1756.580 1704.260 1756.900 1704.580 ;
        RECT 1756.580 1665.500 1756.900 1665.820 ;
        RECT 1756.580 1663.460 1756.900 1663.780 ;
        RECT 1756.580 1608.380 1756.900 1608.700 ;
        RECT 1756.580 1602.260 1756.900 1602.580 ;
        RECT 1756.580 1556.700 1756.900 1557.020 ;
        RECT 1756.580 1513.180 1756.900 1513.500 ;
        RECT 1756.580 1413.220 1756.900 1413.540 ;
        RECT 1764.860 1413.220 1765.180 1413.540 ;
        RECT 1756.580 1360.860 1756.900 1361.180 ;
        RECT 1764.860 1360.860 1765.180 1361.180 ;
        RECT 1756.580 1302.380 1756.900 1302.700 ;
      LAYER met4 ;
        RECT 1756.575 2318.295 1756.905 2318.625 ;
        RECT 1756.590 2309.105 1756.890 2318.295 ;
        RECT 1756.575 2308.775 1756.905 2309.105 ;
        RECT 1756.575 2282.935 1756.905 2283.265 ;
        RECT 1756.590 2188.745 1756.890 2282.935 ;
        RECT 1756.575 2188.415 1756.905 2188.745 ;
        RECT 1756.575 2186.375 1756.905 2186.705 ;
        RECT 1756.590 2133.650 1756.890 2186.375 ;
        RECT 1756.590 2133.350 1758.730 2133.650 ;
        RECT 1758.430 2097.625 1758.730 2133.350 ;
        RECT 1758.415 2097.295 1758.745 2097.625 ;
        RECT 1756.575 2054.455 1756.905 2054.785 ;
        RECT 1756.590 2043.225 1756.890 2054.455 ;
        RECT 1756.575 2042.895 1756.905 2043.225 ;
        RECT 1756.575 1996.655 1756.905 1996.985 ;
        RECT 1756.590 1965.025 1756.890 1996.655 ;
        RECT 1756.575 1964.695 1756.905 1965.025 ;
        RECT 1756.575 1867.455 1756.905 1867.785 ;
        RECT 1756.590 1841.945 1756.890 1867.455 ;
        RECT 1756.575 1841.615 1756.905 1841.945 ;
        RECT 1756.575 1745.735 1756.905 1746.065 ;
        RECT 1756.590 1724.290 1756.890 1745.735 ;
        RECT 1756.590 1723.990 1757.810 1724.290 ;
        RECT 1757.510 1705.945 1757.810 1723.990 ;
        RECT 1757.495 1705.615 1757.825 1705.945 ;
        RECT 1756.575 1704.255 1756.905 1704.585 ;
        RECT 1756.590 1665.825 1756.890 1704.255 ;
        RECT 1756.575 1665.495 1756.905 1665.825 ;
        RECT 1756.575 1663.455 1756.905 1663.785 ;
        RECT 1756.590 1608.705 1756.890 1663.455 ;
        RECT 1756.575 1608.375 1756.905 1608.705 ;
        RECT 1756.575 1602.255 1756.905 1602.585 ;
        RECT 1756.590 1557.025 1756.890 1602.255 ;
        RECT 1756.575 1556.695 1756.905 1557.025 ;
        RECT 1756.575 1513.175 1756.905 1513.505 ;
        RECT 1756.590 1413.545 1756.890 1513.175 ;
        RECT 1756.575 1413.215 1756.905 1413.545 ;
        RECT 1764.855 1413.215 1765.185 1413.545 ;
        RECT 1764.870 1361.185 1765.170 1413.215 ;
        RECT 1756.575 1360.855 1756.905 1361.185 ;
        RECT 1764.855 1360.855 1765.185 1361.185 ;
        RECT 1756.590 1302.705 1756.890 1360.855 ;
        RECT 1756.575 1302.375 1756.905 1302.705 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1876.945 2263.125 1877.115 2311.575 ;
        RECT 1876.945 2166.905 1877.115 2214.675 ;
        RECT 1877.405 2070.005 1877.575 2118.115 ;
        RECT 1877.405 1973.445 1877.575 2021.555 ;
        RECT 1877.405 1876.885 1877.575 1924.995 ;
        RECT 1876.945 1780.325 1877.115 1828.435 ;
        RECT 1877.405 1683.765 1877.575 1731.535 ;
        RECT 1876.945 1587.205 1877.115 1635.315 ;
        RECT 1876.945 1490.645 1877.115 1538.755 ;
        RECT 1876.945 620.925 1877.115 669.375 ;
        RECT 1876.945 524.365 1877.115 572.475 ;
        RECT 1877.405 427.805 1877.575 475.915 ;
        RECT 1876.945 331.245 1877.115 379.355 ;
        RECT 1876.945 234.685 1877.115 282.795 ;
        RECT 1876.945 138.125 1877.115 186.235 ;
        RECT 1882.005 2.805 1882.175 41.395 ;
      LAYER mcon ;
        RECT 1876.945 2311.405 1877.115 2311.575 ;
        RECT 1876.945 2214.505 1877.115 2214.675 ;
        RECT 1877.405 2117.945 1877.575 2118.115 ;
        RECT 1877.405 2021.385 1877.575 2021.555 ;
        RECT 1877.405 1924.825 1877.575 1924.995 ;
        RECT 1876.945 1828.265 1877.115 1828.435 ;
        RECT 1877.405 1731.365 1877.575 1731.535 ;
        RECT 1876.945 1635.145 1877.115 1635.315 ;
        RECT 1876.945 1538.585 1877.115 1538.755 ;
        RECT 1876.945 669.205 1877.115 669.375 ;
        RECT 1876.945 572.305 1877.115 572.475 ;
        RECT 1877.405 475.745 1877.575 475.915 ;
        RECT 1876.945 379.185 1877.115 379.355 ;
        RECT 1876.945 282.625 1877.115 282.795 ;
        RECT 1876.945 186.065 1877.115 186.235 ;
        RECT 1882.005 41.225 1882.175 41.395 ;
      LAYER met1 ;
        RECT 1364.890 2377.180 1365.210 2377.240 ;
        RECT 1877.790 2377.180 1878.110 2377.240 ;
        RECT 1364.890 2377.040 1878.110 2377.180 ;
        RECT 1364.890 2376.980 1365.210 2377.040 ;
        RECT 1877.790 2376.980 1878.110 2377.040 ;
        RECT 1876.870 2311.560 1877.190 2311.620 ;
        RECT 1876.870 2311.420 1877.385 2311.560 ;
        RECT 1876.870 2311.360 1877.190 2311.420 ;
        RECT 1876.870 2263.280 1877.190 2263.340 ;
        RECT 1876.870 2263.140 1877.385 2263.280 ;
        RECT 1876.870 2263.080 1877.190 2263.140 ;
        RECT 1876.870 2214.660 1877.190 2214.720 ;
        RECT 1876.870 2214.520 1877.385 2214.660 ;
        RECT 1876.870 2214.460 1877.190 2214.520 ;
        RECT 1876.870 2167.060 1877.190 2167.120 ;
        RECT 1876.870 2166.920 1877.385 2167.060 ;
        RECT 1876.870 2166.860 1877.190 2166.920 ;
        RECT 1876.870 2118.100 1877.190 2118.160 ;
        RECT 1877.345 2118.100 1877.635 2118.145 ;
        RECT 1876.870 2117.960 1877.635 2118.100 ;
        RECT 1876.870 2117.900 1877.190 2117.960 ;
        RECT 1877.345 2117.915 1877.635 2117.960 ;
        RECT 1876.870 2070.160 1877.190 2070.220 ;
        RECT 1877.345 2070.160 1877.635 2070.205 ;
        RECT 1876.870 2070.020 1877.635 2070.160 ;
        RECT 1876.870 2069.960 1877.190 2070.020 ;
        RECT 1877.345 2069.975 1877.635 2070.020 ;
        RECT 1876.870 2021.540 1877.190 2021.600 ;
        RECT 1877.345 2021.540 1877.635 2021.585 ;
        RECT 1876.870 2021.400 1877.635 2021.540 ;
        RECT 1876.870 2021.340 1877.190 2021.400 ;
        RECT 1877.345 2021.355 1877.635 2021.400 ;
        RECT 1876.870 1973.600 1877.190 1973.660 ;
        RECT 1877.345 1973.600 1877.635 1973.645 ;
        RECT 1876.870 1973.460 1877.635 1973.600 ;
        RECT 1876.870 1973.400 1877.190 1973.460 ;
        RECT 1877.345 1973.415 1877.635 1973.460 ;
        RECT 1876.870 1924.980 1877.190 1925.040 ;
        RECT 1877.345 1924.980 1877.635 1925.025 ;
        RECT 1876.870 1924.840 1877.635 1924.980 ;
        RECT 1876.870 1924.780 1877.190 1924.840 ;
        RECT 1877.345 1924.795 1877.635 1924.840 ;
        RECT 1876.870 1877.040 1877.190 1877.100 ;
        RECT 1877.345 1877.040 1877.635 1877.085 ;
        RECT 1876.870 1876.900 1877.635 1877.040 ;
        RECT 1876.870 1876.840 1877.190 1876.900 ;
        RECT 1877.345 1876.855 1877.635 1876.900 ;
        RECT 1876.870 1828.420 1877.190 1828.480 ;
        RECT 1876.870 1828.280 1877.385 1828.420 ;
        RECT 1876.870 1828.220 1877.190 1828.280 ;
        RECT 1876.870 1780.480 1877.190 1780.540 ;
        RECT 1876.870 1780.340 1877.385 1780.480 ;
        RECT 1876.870 1780.280 1877.190 1780.340 ;
        RECT 1876.870 1731.520 1877.190 1731.580 ;
        RECT 1877.345 1731.520 1877.635 1731.565 ;
        RECT 1876.870 1731.380 1877.635 1731.520 ;
        RECT 1876.870 1731.320 1877.190 1731.380 ;
        RECT 1877.345 1731.335 1877.635 1731.380 ;
        RECT 1876.870 1683.920 1877.190 1683.980 ;
        RECT 1877.345 1683.920 1877.635 1683.965 ;
        RECT 1876.870 1683.780 1877.635 1683.920 ;
        RECT 1876.870 1683.720 1877.190 1683.780 ;
        RECT 1877.345 1683.735 1877.635 1683.780 ;
        RECT 1876.870 1635.300 1877.190 1635.360 ;
        RECT 1876.870 1635.160 1877.385 1635.300 ;
        RECT 1876.870 1635.100 1877.190 1635.160 ;
        RECT 1876.870 1587.360 1877.190 1587.420 ;
        RECT 1876.870 1587.220 1877.385 1587.360 ;
        RECT 1876.870 1587.160 1877.190 1587.220 ;
        RECT 1876.870 1538.740 1877.190 1538.800 ;
        RECT 1876.870 1538.600 1877.385 1538.740 ;
        RECT 1876.870 1538.540 1877.190 1538.600 ;
        RECT 1876.870 1490.800 1877.190 1490.860 ;
        RECT 1876.870 1490.660 1877.385 1490.800 ;
        RECT 1876.870 1490.600 1877.190 1490.660 ;
        RECT 1876.870 1393.900 1877.190 1393.960 ;
        RECT 1877.790 1393.900 1878.110 1393.960 ;
        RECT 1876.870 1393.760 1878.110 1393.900 ;
        RECT 1876.870 1393.700 1877.190 1393.760 ;
        RECT 1877.790 1393.700 1878.110 1393.760 ;
        RECT 1876.870 1297.340 1877.190 1297.400 ;
        RECT 1877.790 1297.340 1878.110 1297.400 ;
        RECT 1876.870 1297.200 1878.110 1297.340 ;
        RECT 1876.870 1297.140 1877.190 1297.200 ;
        RECT 1877.790 1297.140 1878.110 1297.200 ;
        RECT 1876.870 1200.780 1877.190 1200.840 ;
        RECT 1877.790 1200.780 1878.110 1200.840 ;
        RECT 1876.870 1200.640 1878.110 1200.780 ;
        RECT 1876.870 1200.580 1877.190 1200.640 ;
        RECT 1877.790 1200.580 1878.110 1200.640 ;
        RECT 1876.870 1104.220 1877.190 1104.280 ;
        RECT 1877.790 1104.220 1878.110 1104.280 ;
        RECT 1876.870 1104.080 1878.110 1104.220 ;
        RECT 1876.870 1104.020 1877.190 1104.080 ;
        RECT 1877.790 1104.020 1878.110 1104.080 ;
        RECT 1876.870 1055.400 1877.190 1055.660 ;
        RECT 1876.960 1055.260 1877.100 1055.400 ;
        RECT 1877.790 1055.260 1878.110 1055.320 ;
        RECT 1876.960 1055.120 1878.110 1055.260 ;
        RECT 1877.790 1055.060 1878.110 1055.120 ;
        RECT 1876.870 959.040 1877.190 959.100 ;
        RECT 1877.790 959.040 1878.110 959.100 ;
        RECT 1876.870 958.900 1878.110 959.040 ;
        RECT 1876.870 958.840 1877.190 958.900 ;
        RECT 1877.790 958.840 1878.110 958.900 ;
        RECT 1876.870 862.480 1877.190 862.540 ;
        RECT 1877.790 862.480 1878.110 862.540 ;
        RECT 1876.870 862.340 1878.110 862.480 ;
        RECT 1876.870 862.280 1877.190 862.340 ;
        RECT 1877.790 862.280 1878.110 862.340 ;
        RECT 1876.870 765.920 1877.190 765.980 ;
        RECT 1877.790 765.920 1878.110 765.980 ;
        RECT 1876.870 765.780 1878.110 765.920 ;
        RECT 1876.870 765.720 1877.190 765.780 ;
        RECT 1877.790 765.720 1878.110 765.780 ;
        RECT 1876.870 669.360 1877.190 669.420 ;
        RECT 1876.870 669.220 1877.385 669.360 ;
        RECT 1876.870 669.160 1877.190 669.220 ;
        RECT 1876.870 621.080 1877.190 621.140 ;
        RECT 1876.870 620.940 1877.385 621.080 ;
        RECT 1876.870 620.880 1877.190 620.940 ;
        RECT 1876.870 572.460 1877.190 572.520 ;
        RECT 1876.870 572.320 1877.385 572.460 ;
        RECT 1876.870 572.260 1877.190 572.320 ;
        RECT 1876.870 524.520 1877.190 524.580 ;
        RECT 1876.870 524.380 1877.385 524.520 ;
        RECT 1876.870 524.320 1877.190 524.380 ;
        RECT 1876.870 475.900 1877.190 475.960 ;
        RECT 1877.345 475.900 1877.635 475.945 ;
        RECT 1876.870 475.760 1877.635 475.900 ;
        RECT 1876.870 475.700 1877.190 475.760 ;
        RECT 1877.345 475.715 1877.635 475.760 ;
        RECT 1876.870 427.960 1877.190 428.020 ;
        RECT 1877.345 427.960 1877.635 428.005 ;
        RECT 1876.870 427.820 1877.635 427.960 ;
        RECT 1876.870 427.760 1877.190 427.820 ;
        RECT 1877.345 427.775 1877.635 427.820 ;
        RECT 1876.870 379.340 1877.190 379.400 ;
        RECT 1876.870 379.200 1877.385 379.340 ;
        RECT 1876.870 379.140 1877.190 379.200 ;
        RECT 1876.870 331.400 1877.190 331.460 ;
        RECT 1876.870 331.260 1877.385 331.400 ;
        RECT 1876.870 331.200 1877.190 331.260 ;
        RECT 1876.870 282.780 1877.190 282.840 ;
        RECT 1876.870 282.640 1877.385 282.780 ;
        RECT 1876.870 282.580 1877.190 282.640 ;
        RECT 1876.870 234.840 1877.190 234.900 ;
        RECT 1876.870 234.700 1877.385 234.840 ;
        RECT 1876.870 234.640 1877.190 234.700 ;
        RECT 1876.870 186.220 1877.190 186.280 ;
        RECT 1876.870 186.080 1877.385 186.220 ;
        RECT 1876.870 186.020 1877.190 186.080 ;
        RECT 1876.870 138.280 1877.190 138.340 ;
        RECT 1876.870 138.140 1877.385 138.280 ;
        RECT 1876.870 138.080 1877.190 138.140 ;
        RECT 1876.870 41.380 1877.190 41.440 ;
        RECT 1881.945 41.380 1882.235 41.425 ;
        RECT 1876.870 41.240 1882.235 41.380 ;
        RECT 1876.870 41.180 1877.190 41.240 ;
        RECT 1881.945 41.195 1882.235 41.240 ;
        RECT 1881.930 2.960 1882.250 3.020 ;
        RECT 1881.735 2.820 1882.250 2.960 ;
        RECT 1881.930 2.760 1882.250 2.820 ;
      LAYER via ;
        RECT 1364.920 2376.980 1365.180 2377.240 ;
        RECT 1877.820 2376.980 1878.080 2377.240 ;
        RECT 1876.900 2311.360 1877.160 2311.620 ;
        RECT 1876.900 2263.080 1877.160 2263.340 ;
        RECT 1876.900 2214.460 1877.160 2214.720 ;
        RECT 1876.900 2166.860 1877.160 2167.120 ;
        RECT 1876.900 2117.900 1877.160 2118.160 ;
        RECT 1876.900 2069.960 1877.160 2070.220 ;
        RECT 1876.900 2021.340 1877.160 2021.600 ;
        RECT 1876.900 1973.400 1877.160 1973.660 ;
        RECT 1876.900 1924.780 1877.160 1925.040 ;
        RECT 1876.900 1876.840 1877.160 1877.100 ;
        RECT 1876.900 1828.220 1877.160 1828.480 ;
        RECT 1876.900 1780.280 1877.160 1780.540 ;
        RECT 1876.900 1731.320 1877.160 1731.580 ;
        RECT 1876.900 1683.720 1877.160 1683.980 ;
        RECT 1876.900 1635.100 1877.160 1635.360 ;
        RECT 1876.900 1587.160 1877.160 1587.420 ;
        RECT 1876.900 1538.540 1877.160 1538.800 ;
        RECT 1876.900 1490.600 1877.160 1490.860 ;
        RECT 1876.900 1393.700 1877.160 1393.960 ;
        RECT 1877.820 1393.700 1878.080 1393.960 ;
        RECT 1876.900 1297.140 1877.160 1297.400 ;
        RECT 1877.820 1297.140 1878.080 1297.400 ;
        RECT 1876.900 1200.580 1877.160 1200.840 ;
        RECT 1877.820 1200.580 1878.080 1200.840 ;
        RECT 1876.900 1104.020 1877.160 1104.280 ;
        RECT 1877.820 1104.020 1878.080 1104.280 ;
        RECT 1876.900 1055.400 1877.160 1055.660 ;
        RECT 1877.820 1055.060 1878.080 1055.320 ;
        RECT 1876.900 958.840 1877.160 959.100 ;
        RECT 1877.820 958.840 1878.080 959.100 ;
        RECT 1876.900 862.280 1877.160 862.540 ;
        RECT 1877.820 862.280 1878.080 862.540 ;
        RECT 1876.900 765.720 1877.160 765.980 ;
        RECT 1877.820 765.720 1878.080 765.980 ;
        RECT 1876.900 669.160 1877.160 669.420 ;
        RECT 1876.900 620.880 1877.160 621.140 ;
        RECT 1876.900 572.260 1877.160 572.520 ;
        RECT 1876.900 524.320 1877.160 524.580 ;
        RECT 1876.900 475.700 1877.160 475.960 ;
        RECT 1876.900 427.760 1877.160 428.020 ;
        RECT 1876.900 379.140 1877.160 379.400 ;
        RECT 1876.900 331.200 1877.160 331.460 ;
        RECT 1876.900 282.580 1877.160 282.840 ;
        RECT 1876.900 234.640 1877.160 234.900 ;
        RECT 1876.900 186.020 1877.160 186.280 ;
        RECT 1876.900 138.080 1877.160 138.340 ;
        RECT 1876.900 41.180 1877.160 41.440 ;
        RECT 1881.960 2.760 1882.220 3.020 ;
      LAYER met2 ;
        RECT 1363.580 2377.010 1363.860 2377.880 ;
        RECT 1364.920 2377.010 1365.180 2377.270 ;
        RECT 1363.580 2376.950 1365.180 2377.010 ;
        RECT 1877.820 2376.950 1878.080 2377.270 ;
        RECT 1363.580 2376.870 1365.120 2376.950 ;
        RECT 1363.580 2373.880 1363.860 2376.870 ;
        RECT 1877.880 2360.125 1878.020 2376.950 ;
        RECT 1876.890 2359.755 1877.170 2360.125 ;
        RECT 1877.810 2359.755 1878.090 2360.125 ;
        RECT 1876.960 2311.650 1877.100 2359.755 ;
        RECT 1876.900 2311.330 1877.160 2311.650 ;
        RECT 1876.900 2263.050 1877.160 2263.370 ;
        RECT 1876.960 2214.750 1877.100 2263.050 ;
        RECT 1876.900 2214.430 1877.160 2214.750 ;
        RECT 1876.900 2166.830 1877.160 2167.150 ;
        RECT 1876.960 2118.190 1877.100 2166.830 ;
        RECT 1876.900 2117.870 1877.160 2118.190 ;
        RECT 1876.900 2069.930 1877.160 2070.250 ;
        RECT 1876.960 2021.630 1877.100 2069.930 ;
        RECT 1876.900 2021.310 1877.160 2021.630 ;
        RECT 1876.900 1973.370 1877.160 1973.690 ;
        RECT 1876.960 1925.070 1877.100 1973.370 ;
        RECT 1876.900 1924.750 1877.160 1925.070 ;
        RECT 1876.900 1876.810 1877.160 1877.130 ;
        RECT 1876.960 1828.510 1877.100 1876.810 ;
        RECT 1876.900 1828.190 1877.160 1828.510 ;
        RECT 1876.900 1780.250 1877.160 1780.570 ;
        RECT 1876.960 1731.610 1877.100 1780.250 ;
        RECT 1876.900 1731.290 1877.160 1731.610 ;
        RECT 1876.900 1683.690 1877.160 1684.010 ;
        RECT 1876.960 1635.390 1877.100 1683.690 ;
        RECT 1876.900 1635.070 1877.160 1635.390 ;
        RECT 1876.900 1587.130 1877.160 1587.450 ;
        RECT 1876.960 1538.830 1877.100 1587.130 ;
        RECT 1876.900 1538.510 1877.160 1538.830 ;
        RECT 1876.900 1490.570 1877.160 1490.890 ;
        RECT 1876.960 1442.125 1877.100 1490.570 ;
        RECT 1876.890 1441.755 1877.170 1442.125 ;
        RECT 1877.810 1441.755 1878.090 1442.125 ;
        RECT 1877.880 1393.990 1878.020 1441.755 ;
        RECT 1876.900 1393.670 1877.160 1393.990 ;
        RECT 1877.820 1393.670 1878.080 1393.990 ;
        RECT 1876.960 1345.565 1877.100 1393.670 ;
        RECT 1876.890 1345.195 1877.170 1345.565 ;
        RECT 1877.810 1345.195 1878.090 1345.565 ;
        RECT 1877.880 1297.430 1878.020 1345.195 ;
        RECT 1876.900 1297.110 1877.160 1297.430 ;
        RECT 1877.820 1297.110 1878.080 1297.430 ;
        RECT 1876.960 1249.005 1877.100 1297.110 ;
        RECT 1876.890 1248.635 1877.170 1249.005 ;
        RECT 1877.810 1248.635 1878.090 1249.005 ;
        RECT 1877.880 1200.870 1878.020 1248.635 ;
        RECT 1876.900 1200.550 1877.160 1200.870 ;
        RECT 1877.820 1200.550 1878.080 1200.870 ;
        RECT 1876.960 1152.445 1877.100 1200.550 ;
        RECT 1876.890 1152.075 1877.170 1152.445 ;
        RECT 1877.810 1152.075 1878.090 1152.445 ;
        RECT 1877.880 1104.310 1878.020 1152.075 ;
        RECT 1876.900 1103.990 1877.160 1104.310 ;
        RECT 1877.820 1103.990 1878.080 1104.310 ;
        RECT 1876.960 1055.690 1877.100 1103.990 ;
        RECT 1876.900 1055.370 1877.160 1055.690 ;
        RECT 1877.820 1055.030 1878.080 1055.350 ;
        RECT 1877.880 1007.605 1878.020 1055.030 ;
        RECT 1876.890 1007.235 1877.170 1007.605 ;
        RECT 1877.810 1007.235 1878.090 1007.605 ;
        RECT 1876.960 959.130 1877.100 1007.235 ;
        RECT 1876.900 958.810 1877.160 959.130 ;
        RECT 1877.820 958.810 1878.080 959.130 ;
        RECT 1877.880 911.045 1878.020 958.810 ;
        RECT 1876.890 910.675 1877.170 911.045 ;
        RECT 1877.810 910.675 1878.090 911.045 ;
        RECT 1876.960 862.570 1877.100 910.675 ;
        RECT 1876.900 862.250 1877.160 862.570 ;
        RECT 1877.820 862.250 1878.080 862.570 ;
        RECT 1877.880 814.485 1878.020 862.250 ;
        RECT 1876.890 814.115 1877.170 814.485 ;
        RECT 1877.810 814.115 1878.090 814.485 ;
        RECT 1876.960 766.010 1877.100 814.115 ;
        RECT 1876.900 765.690 1877.160 766.010 ;
        RECT 1877.820 765.690 1878.080 766.010 ;
        RECT 1877.880 717.925 1878.020 765.690 ;
        RECT 1876.890 717.555 1877.170 717.925 ;
        RECT 1877.810 717.555 1878.090 717.925 ;
        RECT 1876.960 669.450 1877.100 717.555 ;
        RECT 1876.900 669.130 1877.160 669.450 ;
        RECT 1876.900 620.850 1877.160 621.170 ;
        RECT 1876.960 572.550 1877.100 620.850 ;
        RECT 1876.900 572.230 1877.160 572.550 ;
        RECT 1876.900 524.290 1877.160 524.610 ;
        RECT 1876.960 475.990 1877.100 524.290 ;
        RECT 1876.900 475.670 1877.160 475.990 ;
        RECT 1876.900 427.730 1877.160 428.050 ;
        RECT 1876.960 379.430 1877.100 427.730 ;
        RECT 1876.900 379.110 1877.160 379.430 ;
        RECT 1876.900 331.170 1877.160 331.490 ;
        RECT 1876.960 282.870 1877.100 331.170 ;
        RECT 1876.900 282.550 1877.160 282.870 ;
        RECT 1876.900 234.610 1877.160 234.930 ;
        RECT 1876.960 186.310 1877.100 234.610 ;
        RECT 1876.900 185.990 1877.160 186.310 ;
        RECT 1876.900 138.050 1877.160 138.370 ;
        RECT 1876.960 86.090 1877.100 138.050 ;
        RECT 1876.960 85.950 1877.560 86.090 ;
        RECT 1877.420 41.890 1877.560 85.950 ;
        RECT 1876.960 41.750 1877.560 41.890 ;
        RECT 1876.960 41.470 1877.100 41.750 ;
        RECT 1876.900 41.150 1877.160 41.470 ;
        RECT 1881.960 2.730 1882.220 3.050 ;
        RECT 1882.020 2.400 1882.160 2.730 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
      LAYER via2 ;
        RECT 1876.890 2359.800 1877.170 2360.080 ;
        RECT 1877.810 2359.800 1878.090 2360.080 ;
        RECT 1876.890 1441.800 1877.170 1442.080 ;
        RECT 1877.810 1441.800 1878.090 1442.080 ;
        RECT 1876.890 1345.240 1877.170 1345.520 ;
        RECT 1877.810 1345.240 1878.090 1345.520 ;
        RECT 1876.890 1248.680 1877.170 1248.960 ;
        RECT 1877.810 1248.680 1878.090 1248.960 ;
        RECT 1876.890 1152.120 1877.170 1152.400 ;
        RECT 1877.810 1152.120 1878.090 1152.400 ;
        RECT 1876.890 1007.280 1877.170 1007.560 ;
        RECT 1877.810 1007.280 1878.090 1007.560 ;
        RECT 1876.890 910.720 1877.170 911.000 ;
        RECT 1877.810 910.720 1878.090 911.000 ;
        RECT 1876.890 814.160 1877.170 814.440 ;
        RECT 1877.810 814.160 1878.090 814.440 ;
        RECT 1876.890 717.600 1877.170 717.880 ;
        RECT 1877.810 717.600 1878.090 717.880 ;
      LAYER met3 ;
        RECT 1876.865 2360.090 1877.195 2360.105 ;
        RECT 1877.785 2360.090 1878.115 2360.105 ;
        RECT 1876.865 2359.790 1878.115 2360.090 ;
        RECT 1876.865 2359.775 1877.195 2359.790 ;
        RECT 1877.785 2359.775 1878.115 2359.790 ;
        RECT 1876.865 1442.090 1877.195 1442.105 ;
        RECT 1877.785 1442.090 1878.115 1442.105 ;
        RECT 1876.865 1441.790 1878.115 1442.090 ;
        RECT 1876.865 1441.775 1877.195 1441.790 ;
        RECT 1877.785 1441.775 1878.115 1441.790 ;
        RECT 1876.865 1345.530 1877.195 1345.545 ;
        RECT 1877.785 1345.530 1878.115 1345.545 ;
        RECT 1876.865 1345.230 1878.115 1345.530 ;
        RECT 1876.865 1345.215 1877.195 1345.230 ;
        RECT 1877.785 1345.215 1878.115 1345.230 ;
        RECT 1876.865 1248.970 1877.195 1248.985 ;
        RECT 1877.785 1248.970 1878.115 1248.985 ;
        RECT 1876.865 1248.670 1878.115 1248.970 ;
        RECT 1876.865 1248.655 1877.195 1248.670 ;
        RECT 1877.785 1248.655 1878.115 1248.670 ;
        RECT 1876.865 1152.410 1877.195 1152.425 ;
        RECT 1877.785 1152.410 1878.115 1152.425 ;
        RECT 1876.865 1152.110 1878.115 1152.410 ;
        RECT 1876.865 1152.095 1877.195 1152.110 ;
        RECT 1877.785 1152.095 1878.115 1152.110 ;
        RECT 1876.865 1007.570 1877.195 1007.585 ;
        RECT 1877.785 1007.570 1878.115 1007.585 ;
        RECT 1876.865 1007.270 1878.115 1007.570 ;
        RECT 1876.865 1007.255 1877.195 1007.270 ;
        RECT 1877.785 1007.255 1878.115 1007.270 ;
        RECT 1876.865 911.010 1877.195 911.025 ;
        RECT 1877.785 911.010 1878.115 911.025 ;
        RECT 1876.865 910.710 1878.115 911.010 ;
        RECT 1876.865 910.695 1877.195 910.710 ;
        RECT 1877.785 910.695 1878.115 910.710 ;
        RECT 1876.865 814.450 1877.195 814.465 ;
        RECT 1877.785 814.450 1878.115 814.465 ;
        RECT 1876.865 814.150 1878.115 814.450 ;
        RECT 1876.865 814.135 1877.195 814.150 ;
        RECT 1877.785 814.135 1878.115 814.150 ;
        RECT 1876.865 717.890 1877.195 717.905 ;
        RECT 1877.785 717.890 1878.115 717.905 ;
        RECT 1876.865 717.590 1878.115 717.890 ;
        RECT 1876.865 717.575 1877.195 717.590 ;
        RECT 1877.785 717.575 1878.115 717.590 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1539.230 1311.280 1539.550 1311.340 ;
        RECT 1545.210 1311.280 1545.530 1311.340 ;
        RECT 1539.230 1311.140 1545.530 1311.280 ;
        RECT 1539.230 1311.080 1539.550 1311.140 ;
        RECT 1545.210 1311.080 1545.530 1311.140 ;
        RECT 1545.210 27.100 1545.530 27.160 ;
        RECT 1899.870 27.100 1900.190 27.160 ;
        RECT 1545.210 26.960 1900.190 27.100 ;
        RECT 1545.210 26.900 1545.530 26.960 ;
        RECT 1899.870 26.900 1900.190 26.960 ;
      LAYER via ;
        RECT 1539.260 1311.080 1539.520 1311.340 ;
        RECT 1545.240 1311.080 1545.500 1311.340 ;
        RECT 1545.240 26.900 1545.500 27.160 ;
        RECT 1899.900 26.900 1900.160 27.160 ;
      LAYER met2 ;
        RECT 1539.300 1323.135 1539.580 1327.135 ;
        RECT 1539.320 1311.370 1539.460 1323.135 ;
        RECT 1539.260 1311.050 1539.520 1311.370 ;
        RECT 1545.240 1311.050 1545.500 1311.370 ;
        RECT 1545.300 27.190 1545.440 1311.050 ;
        RECT 1545.240 26.870 1545.500 27.190 ;
        RECT 1899.900 26.870 1900.160 27.190 ;
        RECT 1899.960 2.400 1900.100 26.870 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 708.930 86.600 709.250 86.660 ;
        RECT 1911.830 86.600 1912.150 86.660 ;
        RECT 708.930 86.460 1912.150 86.600 ;
        RECT 708.930 86.400 709.250 86.460 ;
        RECT 1911.830 86.400 1912.150 86.460 ;
        RECT 1911.830 37.640 1912.150 37.700 ;
        RECT 1917.810 37.640 1918.130 37.700 ;
        RECT 1911.830 37.500 1918.130 37.640 ;
        RECT 1911.830 37.440 1912.150 37.500 ;
        RECT 1917.810 37.440 1918.130 37.500 ;
      LAYER via ;
        RECT 708.960 86.400 709.220 86.660 ;
        RECT 1911.860 86.400 1912.120 86.660 ;
        RECT 1911.860 37.440 1912.120 37.700 ;
        RECT 1917.840 37.440 1918.100 37.700 ;
      LAYER met2 ;
        RECT 708.950 1814.395 709.230 1814.765 ;
        RECT 709.020 86.690 709.160 1814.395 ;
        RECT 708.960 86.370 709.220 86.690 ;
        RECT 1911.860 86.370 1912.120 86.690 ;
        RECT 1911.920 37.730 1912.060 86.370 ;
        RECT 1911.860 37.410 1912.120 37.730 ;
        RECT 1917.840 37.410 1918.100 37.730 ;
        RECT 1917.900 2.400 1918.040 37.410 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
      LAYER via2 ;
        RECT 708.950 1814.440 709.230 1814.720 ;
      LAYER met3 ;
        RECT 708.925 1814.730 709.255 1814.745 ;
        RECT 715.810 1814.730 719.810 1814.735 ;
        RECT 708.925 1814.430 719.810 1814.730 ;
        RECT 708.925 1814.415 709.255 1814.430 ;
        RECT 715.810 1814.135 719.810 1814.430 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1346.105 2375.325 1346.735 2375.495 ;
        RECT 1932.145 48.365 1932.315 96.475 ;
      LAYER mcon ;
        RECT 1346.565 2375.325 1346.735 2375.495 ;
        RECT 1932.145 96.305 1932.315 96.475 ;
      LAYER met1 ;
        RECT 815.650 2375.480 815.970 2375.540 ;
        RECT 1346.045 2375.480 1346.335 2375.525 ;
        RECT 815.650 2375.340 1346.335 2375.480 ;
        RECT 815.650 2375.280 815.970 2375.340 ;
        RECT 1346.045 2375.295 1346.335 2375.340 ;
        RECT 1346.505 2375.480 1346.795 2375.525 ;
        RECT 1932.070 2375.480 1932.390 2375.540 ;
        RECT 1346.505 2375.340 1932.390 2375.480 ;
        RECT 1346.505 2375.295 1346.795 2375.340 ;
        RECT 1932.070 2375.280 1932.390 2375.340 ;
        RECT 1932.070 96.460 1932.390 96.520 ;
        RECT 1932.070 96.320 1932.585 96.460 ;
        RECT 1932.070 96.260 1932.390 96.320 ;
        RECT 1932.085 48.520 1932.375 48.565 ;
        RECT 1935.290 48.520 1935.610 48.580 ;
        RECT 1932.085 48.380 1935.610 48.520 ;
        RECT 1932.085 48.335 1932.375 48.380 ;
        RECT 1935.290 48.320 1935.610 48.380 ;
      LAYER via ;
        RECT 815.680 2375.280 815.940 2375.540 ;
        RECT 1932.100 2375.280 1932.360 2375.540 ;
        RECT 1932.100 96.260 1932.360 96.520 ;
        RECT 1935.320 48.320 1935.580 48.580 ;
      LAYER met2 ;
        RECT 814.340 2375.650 814.620 2377.880 ;
        RECT 814.340 2375.570 815.880 2375.650 ;
        RECT 814.340 2375.510 815.940 2375.570 ;
        RECT 814.340 2373.880 814.620 2375.510 ;
        RECT 815.680 2375.250 815.940 2375.510 ;
        RECT 1932.100 2375.250 1932.360 2375.570 ;
        RECT 1932.160 96.550 1932.300 2375.250 ;
        RECT 1932.100 96.230 1932.360 96.550 ;
        RECT 1935.320 48.290 1935.580 48.610 ;
        RECT 1935.380 2.400 1935.520 48.290 ;
        RECT 1935.170 -4.800 1935.730 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1345.645 2375.665 1347.195 2375.835 ;
      LAYER mcon ;
        RECT 1347.025 2375.665 1347.195 2375.835 ;
      LAYER met1 ;
        RECT 937.090 2375.820 937.410 2375.880 ;
        RECT 1345.585 2375.820 1345.875 2375.865 ;
        RECT 937.090 2375.680 1345.875 2375.820 ;
        RECT 937.090 2375.620 937.410 2375.680 ;
        RECT 1345.585 2375.635 1345.875 2375.680 ;
        RECT 1346.965 2375.820 1347.255 2375.865 ;
        RECT 1953.230 2375.820 1953.550 2375.880 ;
        RECT 1346.965 2375.680 1953.550 2375.820 ;
        RECT 1346.965 2375.635 1347.255 2375.680 ;
        RECT 1953.230 2375.620 1953.550 2375.680 ;
      LAYER via ;
        RECT 937.120 2375.620 937.380 2375.880 ;
        RECT 1953.260 2375.620 1953.520 2375.880 ;
      LAYER met2 ;
        RECT 935.780 2375.650 936.060 2377.880 ;
        RECT 937.120 2375.650 937.380 2375.910 ;
        RECT 935.780 2375.590 937.380 2375.650 ;
        RECT 1953.260 2375.590 1953.520 2375.910 ;
        RECT 935.780 2375.510 937.320 2375.590 ;
        RECT 935.780 2373.880 936.060 2375.510 ;
        RECT 1953.320 2.400 1953.460 2375.590 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1111.430 1311.280 1111.750 1311.340 ;
        RECT 1117.410 1311.280 1117.730 1311.340 ;
        RECT 1111.430 1311.140 1117.730 1311.280 ;
        RECT 1111.430 1311.080 1111.750 1311.140 ;
        RECT 1117.410 1311.080 1117.730 1311.140 ;
        RECT 1117.410 24.720 1117.730 24.780 ;
        RECT 1971.170 24.720 1971.490 24.780 ;
        RECT 1117.410 24.580 1971.490 24.720 ;
        RECT 1117.410 24.520 1117.730 24.580 ;
        RECT 1971.170 24.520 1971.490 24.580 ;
      LAYER via ;
        RECT 1111.460 1311.080 1111.720 1311.340 ;
        RECT 1117.440 1311.080 1117.700 1311.340 ;
        RECT 1117.440 24.520 1117.700 24.780 ;
        RECT 1971.200 24.520 1971.460 24.780 ;
      LAYER met2 ;
        RECT 1111.500 1323.135 1111.780 1327.135 ;
        RECT 1111.520 1311.370 1111.660 1323.135 ;
        RECT 1111.460 1311.050 1111.720 1311.370 ;
        RECT 1117.440 1311.050 1117.700 1311.370 ;
        RECT 1117.500 24.810 1117.640 1311.050 ;
        RECT 1117.440 24.490 1117.700 24.810 ;
        RECT 1971.200 24.490 1971.460 24.810 ;
        RECT 1971.260 2.400 1971.400 24.490 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1987.345 1635.485 1987.515 1649.255 ;
        RECT 1987.345 1538.925 1987.515 1587.035 ;
        RECT 1987.345 1442.025 1987.515 1490.475 ;
        RECT 1987.345 862.665 1987.515 910.435 ;
        RECT 1987.345 766.105 1987.515 814.215 ;
        RECT 1987.345 669.545 1987.515 717.655 ;
        RECT 1987.345 572.645 1987.515 620.415 ;
        RECT 1987.345 476.085 1987.515 524.195 ;
        RECT 1987.345 379.525 1987.515 427.635 ;
        RECT 1987.345 282.965 1987.515 331.075 ;
        RECT 1987.345 186.405 1987.515 234.515 ;
      LAYER mcon ;
        RECT 1987.345 1649.085 1987.515 1649.255 ;
        RECT 1987.345 1586.865 1987.515 1587.035 ;
        RECT 1987.345 1490.305 1987.515 1490.475 ;
        RECT 1987.345 910.265 1987.515 910.435 ;
        RECT 1987.345 814.045 1987.515 814.215 ;
        RECT 1987.345 717.485 1987.515 717.655 ;
        RECT 1987.345 620.245 1987.515 620.415 ;
        RECT 1987.345 524.025 1987.515 524.195 ;
        RECT 1987.345 427.465 1987.515 427.635 ;
        RECT 1987.345 330.905 1987.515 331.075 ;
        RECT 1987.345 234.345 1987.515 234.515 ;
      LAYER met1 ;
        RECT 1772.910 1649.240 1773.230 1649.300 ;
        RECT 1987.285 1649.240 1987.575 1649.285 ;
        RECT 1772.910 1649.100 1987.575 1649.240 ;
        RECT 1772.910 1649.040 1773.230 1649.100 ;
        RECT 1987.285 1649.055 1987.575 1649.100 ;
        RECT 1987.270 1635.640 1987.590 1635.700 ;
        RECT 1987.075 1635.500 1987.590 1635.640 ;
        RECT 1987.270 1635.440 1987.590 1635.500 ;
        RECT 1987.270 1587.020 1987.590 1587.080 ;
        RECT 1987.075 1586.880 1987.590 1587.020 ;
        RECT 1987.270 1586.820 1987.590 1586.880 ;
        RECT 1987.270 1539.080 1987.590 1539.140 ;
        RECT 1987.075 1538.940 1987.590 1539.080 ;
        RECT 1987.270 1538.880 1987.590 1538.940 ;
        RECT 1987.270 1490.460 1987.590 1490.520 ;
        RECT 1987.075 1490.320 1987.590 1490.460 ;
        RECT 1987.270 1490.260 1987.590 1490.320 ;
        RECT 1987.270 1442.180 1987.590 1442.240 ;
        RECT 1987.075 1442.040 1987.590 1442.180 ;
        RECT 1987.270 1441.980 1987.590 1442.040 ;
        RECT 1987.270 1345.620 1987.590 1345.680 ;
        RECT 1988.190 1345.620 1988.510 1345.680 ;
        RECT 1987.270 1345.480 1988.510 1345.620 ;
        RECT 1987.270 1345.420 1987.590 1345.480 ;
        RECT 1988.190 1345.420 1988.510 1345.480 ;
        RECT 1987.270 1249.060 1987.590 1249.120 ;
        RECT 1988.190 1249.060 1988.510 1249.120 ;
        RECT 1987.270 1248.920 1988.510 1249.060 ;
        RECT 1987.270 1248.860 1987.590 1248.920 ;
        RECT 1988.190 1248.860 1988.510 1248.920 ;
        RECT 1987.270 1152.500 1987.590 1152.560 ;
        RECT 1988.190 1152.500 1988.510 1152.560 ;
        RECT 1987.270 1152.360 1988.510 1152.500 ;
        RECT 1987.270 1152.300 1987.590 1152.360 ;
        RECT 1988.190 1152.300 1988.510 1152.360 ;
        RECT 1987.270 1007.320 1987.590 1007.380 ;
        RECT 1988.190 1007.320 1988.510 1007.380 ;
        RECT 1987.270 1007.180 1988.510 1007.320 ;
        RECT 1987.270 1007.120 1987.590 1007.180 ;
        RECT 1988.190 1007.120 1988.510 1007.180 ;
        RECT 1987.270 910.420 1987.590 910.480 ;
        RECT 1987.075 910.280 1987.590 910.420 ;
        RECT 1987.270 910.220 1987.590 910.280 ;
        RECT 1987.270 862.820 1987.590 862.880 ;
        RECT 1987.075 862.680 1987.590 862.820 ;
        RECT 1987.270 862.620 1987.590 862.680 ;
        RECT 1987.270 814.200 1987.590 814.260 ;
        RECT 1987.075 814.060 1987.590 814.200 ;
        RECT 1987.270 814.000 1987.590 814.060 ;
        RECT 1987.270 766.260 1987.590 766.320 ;
        RECT 1987.075 766.120 1987.590 766.260 ;
        RECT 1987.270 766.060 1987.590 766.120 ;
        RECT 1987.270 717.640 1987.590 717.700 ;
        RECT 1987.075 717.500 1987.590 717.640 ;
        RECT 1987.270 717.440 1987.590 717.500 ;
        RECT 1987.270 669.700 1987.590 669.760 ;
        RECT 1987.075 669.560 1987.590 669.700 ;
        RECT 1987.270 669.500 1987.590 669.560 ;
        RECT 1987.270 620.400 1987.590 620.460 ;
        RECT 1987.075 620.260 1987.590 620.400 ;
        RECT 1987.270 620.200 1987.590 620.260 ;
        RECT 1987.270 572.800 1987.590 572.860 ;
        RECT 1987.075 572.660 1987.590 572.800 ;
        RECT 1987.270 572.600 1987.590 572.660 ;
        RECT 1987.270 524.180 1987.590 524.240 ;
        RECT 1987.075 524.040 1987.590 524.180 ;
        RECT 1987.270 523.980 1987.590 524.040 ;
        RECT 1987.270 476.240 1987.590 476.300 ;
        RECT 1987.075 476.100 1987.590 476.240 ;
        RECT 1987.270 476.040 1987.590 476.100 ;
        RECT 1987.270 427.620 1987.590 427.680 ;
        RECT 1987.075 427.480 1987.590 427.620 ;
        RECT 1987.270 427.420 1987.590 427.480 ;
        RECT 1987.270 379.680 1987.590 379.740 ;
        RECT 1987.075 379.540 1987.590 379.680 ;
        RECT 1987.270 379.480 1987.590 379.540 ;
        RECT 1987.270 331.060 1987.590 331.120 ;
        RECT 1987.075 330.920 1987.590 331.060 ;
        RECT 1987.270 330.860 1987.590 330.920 ;
        RECT 1987.270 283.120 1987.590 283.180 ;
        RECT 1987.075 282.980 1987.590 283.120 ;
        RECT 1987.270 282.920 1987.590 282.980 ;
        RECT 1987.270 234.500 1987.590 234.560 ;
        RECT 1987.075 234.360 1987.590 234.500 ;
        RECT 1987.270 234.300 1987.590 234.360 ;
        RECT 1987.270 186.560 1987.590 186.620 ;
        RECT 1987.075 186.420 1987.590 186.560 ;
        RECT 1987.270 186.360 1987.590 186.420 ;
        RECT 1987.270 137.940 1987.590 138.000 ;
        RECT 1988.650 137.940 1988.970 138.000 ;
        RECT 1987.270 137.800 1988.970 137.940 ;
        RECT 1987.270 137.740 1987.590 137.800 ;
        RECT 1988.650 137.740 1988.970 137.800 ;
        RECT 1989.110 47.980 1989.430 48.240 ;
        RECT 1989.200 47.560 1989.340 47.980 ;
        RECT 1989.110 47.300 1989.430 47.560 ;
      LAYER via ;
        RECT 1772.940 1649.040 1773.200 1649.300 ;
        RECT 1987.300 1635.440 1987.560 1635.700 ;
        RECT 1987.300 1586.820 1987.560 1587.080 ;
        RECT 1987.300 1538.880 1987.560 1539.140 ;
        RECT 1987.300 1490.260 1987.560 1490.520 ;
        RECT 1987.300 1441.980 1987.560 1442.240 ;
        RECT 1987.300 1345.420 1987.560 1345.680 ;
        RECT 1988.220 1345.420 1988.480 1345.680 ;
        RECT 1987.300 1248.860 1987.560 1249.120 ;
        RECT 1988.220 1248.860 1988.480 1249.120 ;
        RECT 1987.300 1152.300 1987.560 1152.560 ;
        RECT 1988.220 1152.300 1988.480 1152.560 ;
        RECT 1987.300 1007.120 1987.560 1007.380 ;
        RECT 1988.220 1007.120 1988.480 1007.380 ;
        RECT 1987.300 910.220 1987.560 910.480 ;
        RECT 1987.300 862.620 1987.560 862.880 ;
        RECT 1987.300 814.000 1987.560 814.260 ;
        RECT 1987.300 766.060 1987.560 766.320 ;
        RECT 1987.300 717.440 1987.560 717.700 ;
        RECT 1987.300 669.500 1987.560 669.760 ;
        RECT 1987.300 620.200 1987.560 620.460 ;
        RECT 1987.300 572.600 1987.560 572.860 ;
        RECT 1987.300 523.980 1987.560 524.240 ;
        RECT 1987.300 476.040 1987.560 476.300 ;
        RECT 1987.300 427.420 1987.560 427.680 ;
        RECT 1987.300 379.480 1987.560 379.740 ;
        RECT 1987.300 330.860 1987.560 331.120 ;
        RECT 1987.300 282.920 1987.560 283.180 ;
        RECT 1987.300 234.300 1987.560 234.560 ;
        RECT 1987.300 186.360 1987.560 186.620 ;
        RECT 1987.300 137.740 1987.560 138.000 ;
        RECT 1988.680 137.740 1988.940 138.000 ;
        RECT 1989.140 47.980 1989.400 48.240 ;
        RECT 1989.140 47.300 1989.400 47.560 ;
      LAYER met2 ;
        RECT 1772.930 1655.275 1773.210 1655.645 ;
        RECT 1773.000 1649.330 1773.140 1655.275 ;
        RECT 1772.940 1649.010 1773.200 1649.330 ;
        RECT 1987.300 1635.410 1987.560 1635.730 ;
        RECT 1987.360 1587.110 1987.500 1635.410 ;
        RECT 1987.300 1586.790 1987.560 1587.110 ;
        RECT 1987.300 1538.850 1987.560 1539.170 ;
        RECT 1987.360 1490.550 1987.500 1538.850 ;
        RECT 1987.300 1490.230 1987.560 1490.550 ;
        RECT 1987.300 1441.950 1987.560 1442.270 ;
        RECT 1987.360 1393.845 1987.500 1441.950 ;
        RECT 1987.290 1393.475 1987.570 1393.845 ;
        RECT 1988.210 1393.475 1988.490 1393.845 ;
        RECT 1988.280 1345.710 1988.420 1393.475 ;
        RECT 1987.300 1345.390 1987.560 1345.710 ;
        RECT 1988.220 1345.390 1988.480 1345.710 ;
        RECT 1987.360 1297.285 1987.500 1345.390 ;
        RECT 1987.290 1296.915 1987.570 1297.285 ;
        RECT 1988.210 1296.915 1988.490 1297.285 ;
        RECT 1988.280 1249.150 1988.420 1296.915 ;
        RECT 1987.300 1248.830 1987.560 1249.150 ;
        RECT 1988.220 1248.830 1988.480 1249.150 ;
        RECT 1987.360 1200.725 1987.500 1248.830 ;
        RECT 1987.290 1200.355 1987.570 1200.725 ;
        RECT 1988.210 1200.355 1988.490 1200.725 ;
        RECT 1988.280 1152.590 1988.420 1200.355 ;
        RECT 1987.300 1152.270 1987.560 1152.590 ;
        RECT 1988.220 1152.270 1988.480 1152.590 ;
        RECT 1987.360 1104.165 1987.500 1152.270 ;
        RECT 1987.290 1103.795 1987.570 1104.165 ;
        RECT 1988.210 1103.795 1988.490 1104.165 ;
        RECT 1988.280 1055.885 1988.420 1103.795 ;
        RECT 1987.290 1055.515 1987.570 1055.885 ;
        RECT 1988.210 1055.515 1988.490 1055.885 ;
        RECT 1987.360 1007.410 1987.500 1055.515 ;
        RECT 1987.300 1007.090 1987.560 1007.410 ;
        RECT 1988.220 1007.090 1988.480 1007.410 ;
        RECT 1988.280 959.325 1988.420 1007.090 ;
        RECT 1987.290 958.955 1987.570 959.325 ;
        RECT 1988.210 958.955 1988.490 959.325 ;
        RECT 1987.360 910.510 1987.500 958.955 ;
        RECT 1987.300 910.190 1987.560 910.510 ;
        RECT 1987.300 862.590 1987.560 862.910 ;
        RECT 1987.360 814.290 1987.500 862.590 ;
        RECT 1987.300 813.970 1987.560 814.290 ;
        RECT 1987.300 766.030 1987.560 766.350 ;
        RECT 1987.360 717.730 1987.500 766.030 ;
        RECT 1987.300 717.410 1987.560 717.730 ;
        RECT 1987.300 669.470 1987.560 669.790 ;
        RECT 1987.360 620.490 1987.500 669.470 ;
        RECT 1987.300 620.170 1987.560 620.490 ;
        RECT 1987.300 572.570 1987.560 572.890 ;
        RECT 1987.360 524.270 1987.500 572.570 ;
        RECT 1987.300 523.950 1987.560 524.270 ;
        RECT 1987.300 476.010 1987.560 476.330 ;
        RECT 1987.360 427.710 1987.500 476.010 ;
        RECT 1987.300 427.390 1987.560 427.710 ;
        RECT 1987.300 379.450 1987.560 379.770 ;
        RECT 1987.360 331.150 1987.500 379.450 ;
        RECT 1987.300 330.830 1987.560 331.150 ;
        RECT 1987.300 282.890 1987.560 283.210 ;
        RECT 1987.360 234.590 1987.500 282.890 ;
        RECT 1987.300 234.270 1987.560 234.590 ;
        RECT 1987.300 186.330 1987.560 186.650 ;
        RECT 1987.360 138.030 1987.500 186.330 ;
        RECT 1987.300 137.710 1987.560 138.030 ;
        RECT 1988.680 137.710 1988.940 138.030 ;
        RECT 1988.740 48.690 1988.880 137.710 ;
        RECT 1988.740 48.550 1989.340 48.690 ;
        RECT 1989.200 48.270 1989.340 48.550 ;
        RECT 1989.140 47.950 1989.400 48.270 ;
        RECT 1989.140 47.270 1989.400 47.590 ;
        RECT 1989.200 2.400 1989.340 47.270 ;
        RECT 1988.990 -4.800 1989.550 2.400 ;
      LAYER via2 ;
        RECT 1772.930 1655.320 1773.210 1655.600 ;
        RECT 1987.290 1393.520 1987.570 1393.800 ;
        RECT 1988.210 1393.520 1988.490 1393.800 ;
        RECT 1987.290 1296.960 1987.570 1297.240 ;
        RECT 1988.210 1296.960 1988.490 1297.240 ;
        RECT 1987.290 1200.400 1987.570 1200.680 ;
        RECT 1988.210 1200.400 1988.490 1200.680 ;
        RECT 1987.290 1103.840 1987.570 1104.120 ;
        RECT 1988.210 1103.840 1988.490 1104.120 ;
        RECT 1987.290 1055.560 1987.570 1055.840 ;
        RECT 1988.210 1055.560 1988.490 1055.840 ;
        RECT 1987.290 959.000 1987.570 959.280 ;
        RECT 1988.210 959.000 1988.490 959.280 ;
      LAYER met3 ;
        RECT 1755.835 1655.610 1759.835 1655.615 ;
        RECT 1772.905 1655.610 1773.235 1655.625 ;
        RECT 1755.835 1655.310 1773.235 1655.610 ;
        RECT 1755.835 1655.015 1759.835 1655.310 ;
        RECT 1772.905 1655.295 1773.235 1655.310 ;
        RECT 1987.265 1393.810 1987.595 1393.825 ;
        RECT 1988.185 1393.810 1988.515 1393.825 ;
        RECT 1987.265 1393.510 1988.515 1393.810 ;
        RECT 1987.265 1393.495 1987.595 1393.510 ;
        RECT 1988.185 1393.495 1988.515 1393.510 ;
        RECT 1987.265 1297.250 1987.595 1297.265 ;
        RECT 1988.185 1297.250 1988.515 1297.265 ;
        RECT 1987.265 1296.950 1988.515 1297.250 ;
        RECT 1987.265 1296.935 1987.595 1296.950 ;
        RECT 1988.185 1296.935 1988.515 1296.950 ;
        RECT 1987.265 1200.690 1987.595 1200.705 ;
        RECT 1988.185 1200.690 1988.515 1200.705 ;
        RECT 1987.265 1200.390 1988.515 1200.690 ;
        RECT 1987.265 1200.375 1987.595 1200.390 ;
        RECT 1988.185 1200.375 1988.515 1200.390 ;
        RECT 1987.265 1104.130 1987.595 1104.145 ;
        RECT 1988.185 1104.130 1988.515 1104.145 ;
        RECT 1987.265 1103.830 1988.515 1104.130 ;
        RECT 1987.265 1103.815 1987.595 1103.830 ;
        RECT 1988.185 1103.815 1988.515 1103.830 ;
        RECT 1987.265 1055.850 1987.595 1055.865 ;
        RECT 1988.185 1055.850 1988.515 1055.865 ;
        RECT 1987.265 1055.550 1988.515 1055.850 ;
        RECT 1987.265 1055.535 1987.595 1055.550 ;
        RECT 1988.185 1055.535 1988.515 1055.550 ;
        RECT 1987.265 959.290 1987.595 959.305 ;
        RECT 1988.185 959.290 1988.515 959.305 ;
        RECT 1987.265 958.990 1988.515 959.290 ;
        RECT 1987.265 958.975 1987.595 958.990 ;
        RECT 1988.185 958.975 1988.515 958.990 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1768.310 1387.100 1768.630 1387.160 ;
        RECT 2001.070 1387.100 2001.390 1387.160 ;
        RECT 1768.310 1386.960 2001.390 1387.100 ;
        RECT 1768.310 1386.900 1768.630 1386.960 ;
        RECT 2001.070 1386.900 2001.390 1386.960 ;
      LAYER via ;
        RECT 1768.340 1386.900 1768.600 1387.160 ;
        RECT 2001.100 1386.900 2001.360 1387.160 ;
      LAYER met2 ;
        RECT 1768.330 1390.075 1768.610 1390.445 ;
        RECT 1768.400 1387.190 1768.540 1390.075 ;
        RECT 1768.340 1386.870 1768.600 1387.190 ;
        RECT 2001.100 1386.870 2001.360 1387.190 ;
        RECT 2001.160 41.210 2001.300 1386.870 ;
        RECT 2001.160 41.070 2001.760 41.210 ;
        RECT 2001.620 19.450 2001.760 41.070 ;
        RECT 2001.620 19.310 2006.820 19.450 ;
        RECT 2006.680 2.400 2006.820 19.310 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
      LAYER via2 ;
        RECT 1768.330 1390.120 1768.610 1390.400 ;
      LAYER met3 ;
        RECT 1755.835 1390.410 1759.835 1390.415 ;
        RECT 1768.305 1390.410 1768.635 1390.425 ;
        RECT 1755.835 1390.110 1768.635 1390.410 ;
        RECT 1755.835 1389.815 1759.835 1390.110 ;
        RECT 1768.305 1390.095 1768.635 1390.110 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 692.445 1368.925 692.615 1393.575 ;
      LAYER mcon ;
        RECT 692.445 1393.405 692.615 1393.575 ;
      LAYER met1 ;
        RECT 692.370 1649.240 692.690 1649.300 ;
        RECT 707.550 1649.240 707.870 1649.300 ;
        RECT 692.370 1649.100 707.870 1649.240 ;
        RECT 692.370 1649.040 692.690 1649.100 ;
        RECT 707.550 1649.040 707.870 1649.100 ;
        RECT 692.370 1393.560 692.690 1393.620 ;
        RECT 692.370 1393.420 692.885 1393.560 ;
        RECT 692.370 1393.360 692.690 1393.420 ;
        RECT 692.370 1369.080 692.690 1369.140 ;
        RECT 692.175 1368.940 692.690 1369.080 ;
        RECT 692.370 1368.880 692.690 1368.940 ;
        RECT 692.830 17.240 693.150 17.300 ;
        RECT 2024.530 17.240 2024.850 17.300 ;
        RECT 692.830 17.100 2024.850 17.240 ;
        RECT 692.830 17.040 693.150 17.100 ;
        RECT 2024.530 17.040 2024.850 17.100 ;
      LAYER via ;
        RECT 692.400 1649.040 692.660 1649.300 ;
        RECT 707.580 1649.040 707.840 1649.300 ;
        RECT 692.400 1393.360 692.660 1393.620 ;
        RECT 692.400 1368.880 692.660 1369.140 ;
        RECT 692.860 17.040 693.120 17.300 ;
        RECT 2024.560 17.040 2024.820 17.300 ;
      LAYER met2 ;
        RECT 707.570 1651.195 707.850 1651.565 ;
        RECT 707.640 1649.330 707.780 1651.195 ;
        RECT 692.400 1649.010 692.660 1649.330 ;
        RECT 707.580 1649.010 707.840 1649.330 ;
        RECT 692.460 1393.650 692.600 1649.010 ;
        RECT 692.400 1393.330 692.660 1393.650 ;
        RECT 692.400 1368.850 692.660 1369.170 ;
        RECT 692.460 60.930 692.600 1368.850 ;
        RECT 692.460 60.790 693.060 60.930 ;
        RECT 692.920 17.330 693.060 60.790 ;
        RECT 692.860 17.010 693.120 17.330 ;
        RECT 2024.560 17.010 2024.820 17.330 ;
        RECT 2024.620 2.400 2024.760 17.010 ;
        RECT 2024.410 -4.800 2024.970 2.400 ;
      LAYER via2 ;
        RECT 707.570 1651.240 707.850 1651.520 ;
      LAYER met3 ;
        RECT 707.545 1651.530 707.875 1651.545 ;
        RECT 715.810 1651.530 719.810 1651.535 ;
        RECT 707.545 1651.230 719.810 1651.530 ;
        RECT 707.545 1651.215 707.875 1651.230 ;
        RECT 715.810 1650.935 719.810 1651.230 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1628.010 25.060 1628.330 25.120 ;
        RECT 2042.470 25.060 2042.790 25.120 ;
        RECT 1628.010 24.920 2042.790 25.060 ;
        RECT 1628.010 24.860 1628.330 24.920 ;
        RECT 2042.470 24.860 2042.790 24.920 ;
      LAYER via ;
        RECT 1628.040 24.860 1628.300 25.120 ;
        RECT 2042.500 24.860 2042.760 25.120 ;
      LAYER met2 ;
        RECT 1626.700 1323.690 1626.980 1327.135 ;
        RECT 1626.700 1323.550 1628.240 1323.690 ;
        RECT 1626.700 1323.135 1626.980 1323.550 ;
        RECT 1628.100 25.150 1628.240 1323.550 ;
        RECT 1628.040 24.830 1628.300 25.150 ;
        RECT 2042.500 24.830 2042.760 25.150 ;
        RECT 2042.560 2.400 2042.700 24.830 ;
        RECT 2042.350 -4.800 2042.910 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 758.685 628.065 758.855 676.175 ;
        RECT 758.685 282.965 758.855 331.075 ;
        RECT 758.685 186.405 758.855 234.515 ;
        RECT 757.765 61.965 757.935 137.955 ;
        RECT 757.765 2.805 757.935 48.195 ;
      LAYER mcon ;
        RECT 758.685 676.005 758.855 676.175 ;
        RECT 758.685 330.905 758.855 331.075 ;
        RECT 758.685 234.345 758.855 234.515 ;
        RECT 757.765 137.785 757.935 137.955 ;
        RECT 757.765 48.025 757.935 48.195 ;
      LAYER met1 ;
        RECT 758.610 869.620 758.930 869.680 ;
        RECT 759.070 869.620 759.390 869.680 ;
        RECT 758.610 869.480 759.390 869.620 ;
        RECT 758.610 869.420 758.930 869.480 ;
        RECT 759.070 869.420 759.390 869.480 ;
        RECT 758.610 676.160 758.930 676.220 ;
        RECT 758.415 676.020 758.930 676.160 ;
        RECT 758.610 675.960 758.930 676.020 ;
        RECT 758.610 628.220 758.930 628.280 ;
        RECT 758.415 628.080 758.930 628.220 ;
        RECT 758.610 628.020 758.930 628.080 ;
        RECT 758.610 339.020 758.930 339.280 ;
        RECT 758.700 338.260 758.840 339.020 ;
        RECT 758.610 338.000 758.930 338.260 ;
        RECT 758.610 331.060 758.930 331.120 ;
        RECT 758.415 330.920 758.930 331.060 ;
        RECT 758.610 330.860 758.930 330.920 ;
        RECT 758.610 283.120 758.930 283.180 ;
        RECT 758.415 282.980 758.930 283.120 ;
        RECT 758.610 282.920 758.930 282.980 ;
        RECT 758.610 242.460 758.930 242.720 ;
        RECT 758.700 241.700 758.840 242.460 ;
        RECT 758.610 241.440 758.930 241.700 ;
        RECT 758.610 234.500 758.930 234.560 ;
        RECT 758.415 234.360 758.930 234.500 ;
        RECT 758.610 234.300 758.930 234.360 ;
        RECT 758.610 186.560 758.930 186.620 ;
        RECT 758.415 186.420 758.930 186.560 ;
        RECT 758.610 186.360 758.930 186.420 ;
        RECT 757.705 137.940 757.995 137.985 ;
        RECT 758.610 137.940 758.930 138.000 ;
        RECT 757.705 137.800 758.930 137.940 ;
        RECT 757.705 137.755 757.995 137.800 ;
        RECT 758.610 137.740 758.930 137.800 ;
        RECT 757.690 62.120 758.010 62.180 ;
        RECT 757.495 61.980 758.010 62.120 ;
        RECT 757.690 61.920 758.010 61.980 ;
        RECT 757.690 48.180 758.010 48.240 ;
        RECT 757.495 48.040 758.010 48.180 ;
        RECT 757.690 47.980 758.010 48.040 ;
        RECT 757.690 2.960 758.010 3.020 ;
        RECT 757.495 2.820 758.010 2.960 ;
        RECT 757.690 2.760 758.010 2.820 ;
      LAYER via ;
        RECT 758.640 869.420 758.900 869.680 ;
        RECT 759.100 869.420 759.360 869.680 ;
        RECT 758.640 675.960 758.900 676.220 ;
        RECT 758.640 628.020 758.900 628.280 ;
        RECT 758.640 339.020 758.900 339.280 ;
        RECT 758.640 338.000 758.900 338.260 ;
        RECT 758.640 330.860 758.900 331.120 ;
        RECT 758.640 282.920 758.900 283.180 ;
        RECT 758.640 242.460 758.900 242.720 ;
        RECT 758.640 241.440 758.900 241.700 ;
        RECT 758.640 234.300 758.900 234.560 ;
        RECT 758.640 186.360 758.900 186.620 ;
        RECT 758.640 137.740 758.900 138.000 ;
        RECT 757.720 61.920 757.980 62.180 ;
        RECT 757.720 47.980 757.980 48.240 ;
        RECT 757.720 2.760 757.980 3.020 ;
      LAYER met2 ;
        RECT 758.630 1301.675 758.910 1302.045 ;
        RECT 758.700 917.730 758.840 1301.675 ;
        RECT 758.700 917.590 759.300 917.730 ;
        RECT 759.160 869.710 759.300 917.590 ;
        RECT 758.640 869.565 758.900 869.710 ;
        RECT 758.630 869.195 758.910 869.565 ;
        RECT 759.100 869.390 759.360 869.710 ;
        RECT 757.710 868.515 757.990 868.885 ;
        RECT 757.780 773.005 757.920 868.515 ;
        RECT 757.710 772.635 757.990 773.005 ;
        RECT 758.630 772.635 758.910 773.005 ;
        RECT 758.700 677.805 758.840 772.635 ;
        RECT 758.630 677.435 758.910 677.805 ;
        RECT 758.630 676.075 758.910 676.445 ;
        RECT 758.640 675.930 758.900 676.075 ;
        RECT 758.640 627.990 758.900 628.310 ;
        RECT 758.700 339.310 758.840 627.990 ;
        RECT 758.640 338.990 758.900 339.310 ;
        RECT 758.640 337.970 758.900 338.290 ;
        RECT 758.700 331.150 758.840 337.970 ;
        RECT 758.640 330.830 758.900 331.150 ;
        RECT 758.640 282.890 758.900 283.210 ;
        RECT 758.700 242.750 758.840 282.890 ;
        RECT 758.640 242.430 758.900 242.750 ;
        RECT 758.640 241.410 758.900 241.730 ;
        RECT 758.700 234.590 758.840 241.410 ;
        RECT 758.640 234.270 758.900 234.590 ;
        RECT 758.640 186.330 758.900 186.650 ;
        RECT 758.700 138.030 758.840 186.330 ;
        RECT 758.640 137.710 758.900 138.030 ;
        RECT 757.720 61.890 757.980 62.210 ;
        RECT 757.780 48.270 757.920 61.890 ;
        RECT 757.720 47.950 757.980 48.270 ;
        RECT 757.720 2.730 757.980 3.050 ;
        RECT 757.780 2.400 757.920 2.730 ;
        RECT 757.570 -4.800 758.130 2.400 ;
      LAYER via2 ;
        RECT 758.630 1301.720 758.910 1302.000 ;
        RECT 758.630 869.240 758.910 869.520 ;
        RECT 757.710 868.560 757.990 868.840 ;
        RECT 757.710 772.680 757.990 772.960 ;
        RECT 758.630 772.680 758.910 772.960 ;
        RECT 758.630 677.480 758.910 677.760 ;
        RECT 758.630 676.120 758.910 676.400 ;
      LAYER met3 ;
        RECT 1755.835 1938.490 1759.835 1938.495 ;
        RECT 1772.190 1938.490 1772.570 1938.500 ;
        RECT 1755.835 1938.190 1772.570 1938.490 ;
        RECT 1755.835 1937.895 1759.835 1938.190 ;
        RECT 1772.190 1938.180 1772.570 1938.190 ;
        RECT 758.605 1302.010 758.935 1302.025 ;
        RECT 1772.190 1302.010 1772.570 1302.020 ;
        RECT 758.605 1301.710 1772.570 1302.010 ;
        RECT 758.605 1301.695 758.935 1301.710 ;
        RECT 1772.190 1301.700 1772.570 1301.710 ;
        RECT 758.605 869.530 758.935 869.545 ;
        RECT 758.390 869.215 758.935 869.530 ;
        RECT 757.685 868.850 758.015 868.865 ;
        RECT 758.390 868.850 758.690 869.215 ;
        RECT 757.685 868.550 758.690 868.850 ;
        RECT 757.685 868.535 758.015 868.550 ;
        RECT 757.685 772.970 758.015 772.985 ;
        RECT 758.605 772.970 758.935 772.985 ;
        RECT 757.685 772.670 758.935 772.970 ;
        RECT 757.685 772.655 758.015 772.670 ;
        RECT 758.605 772.655 758.935 772.670 ;
        RECT 758.605 677.770 758.935 677.785 ;
        RECT 758.390 677.455 758.935 677.770 ;
        RECT 758.390 676.425 758.690 677.455 ;
        RECT 758.390 676.110 758.935 676.425 ;
        RECT 758.605 676.095 758.935 676.110 ;
      LAYER via3 ;
        RECT 1772.220 1938.180 1772.540 1938.500 ;
        RECT 1772.220 1301.700 1772.540 1302.020 ;
      LAYER met4 ;
        RECT 1772.215 1938.175 1772.545 1938.505 ;
        RECT 1772.230 1302.025 1772.530 1938.175 ;
        RECT 1772.215 1301.695 1772.545 1302.025 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1531.410 53.620 1531.730 53.680 ;
        RECT 2056.270 53.620 2056.590 53.680 ;
        RECT 1531.410 53.480 2056.590 53.620 ;
        RECT 1531.410 53.420 1531.730 53.480 ;
        RECT 2056.270 53.420 2056.590 53.480 ;
        RECT 2056.270 2.960 2056.590 3.020 ;
        RECT 2060.410 2.960 2060.730 3.020 ;
        RECT 2056.270 2.820 2060.730 2.960 ;
        RECT 2056.270 2.760 2056.590 2.820 ;
        RECT 2060.410 2.760 2060.730 2.820 ;
      LAYER via ;
        RECT 1531.440 53.420 1531.700 53.680 ;
        RECT 2056.300 53.420 2056.560 53.680 ;
        RECT 2056.300 2.760 2056.560 3.020 ;
        RECT 2060.440 2.760 2060.700 3.020 ;
      LAYER met2 ;
        RECT 1528.260 1323.690 1528.540 1327.135 ;
        RECT 1528.260 1323.550 1531.640 1323.690 ;
        RECT 1528.260 1323.135 1528.540 1323.550 ;
        RECT 1531.500 53.710 1531.640 1323.550 ;
        RECT 1531.440 53.390 1531.700 53.710 ;
        RECT 2056.300 53.390 2056.560 53.710 ;
        RECT 2056.360 3.050 2056.500 53.390 ;
        RECT 2056.300 2.730 2056.560 3.050 ;
        RECT 2060.440 2.730 2060.700 3.050 ;
        RECT 2060.500 2.400 2060.640 2.730 ;
        RECT 2060.290 -4.800 2060.850 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1713.110 1311.280 1713.430 1311.340 ;
        RECT 1717.710 1311.280 1718.030 1311.340 ;
        RECT 1713.110 1311.140 1718.030 1311.280 ;
        RECT 1713.110 1311.080 1713.430 1311.140 ;
        RECT 1717.710 1311.080 1718.030 1311.140 ;
        RECT 1717.710 26.080 1718.030 26.140 ;
        RECT 2078.350 26.080 2078.670 26.140 ;
        RECT 1717.710 25.940 2078.670 26.080 ;
        RECT 1717.710 25.880 1718.030 25.940 ;
        RECT 2078.350 25.880 2078.670 25.940 ;
      LAYER via ;
        RECT 1713.140 1311.080 1713.400 1311.340 ;
        RECT 1717.740 1311.080 1718.000 1311.340 ;
        RECT 1717.740 25.880 1718.000 26.140 ;
        RECT 2078.380 25.880 2078.640 26.140 ;
      LAYER met2 ;
        RECT 1713.180 1323.135 1713.460 1327.135 ;
        RECT 1713.200 1311.370 1713.340 1323.135 ;
        RECT 1713.140 1311.050 1713.400 1311.370 ;
        RECT 1717.740 1311.050 1718.000 1311.370 ;
        RECT 1717.800 26.170 1717.940 1311.050 ;
        RECT 1717.740 25.850 1718.000 26.170 ;
        RECT 2078.380 25.850 2078.640 26.170 ;
        RECT 2078.440 2.400 2078.580 25.850 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1771.070 2284.020 1771.390 2284.080 ;
        RECT 2090.770 2284.020 2091.090 2284.080 ;
        RECT 1771.070 2283.880 2091.090 2284.020 ;
        RECT 1771.070 2283.820 1771.390 2283.880 ;
        RECT 2090.770 2283.820 2091.090 2283.880 ;
      LAYER via ;
        RECT 1771.100 2283.820 1771.360 2284.080 ;
        RECT 2090.800 2283.820 2091.060 2284.080 ;
      LAYER met2 ;
        RECT 1771.090 2289.035 1771.370 2289.405 ;
        RECT 1771.160 2284.110 1771.300 2289.035 ;
        RECT 1771.100 2283.790 1771.360 2284.110 ;
        RECT 2090.800 2283.790 2091.060 2284.110 ;
        RECT 2090.860 24.720 2091.000 2283.790 ;
        RECT 2090.860 24.580 2096.060 24.720 ;
        RECT 2095.920 2.400 2096.060 24.580 ;
        RECT 2095.710 -4.800 2096.270 2.400 ;
      LAYER via2 ;
        RECT 1771.090 2289.080 1771.370 2289.360 ;
      LAYER met3 ;
        RECT 1755.835 2289.370 1759.835 2289.375 ;
        RECT 1771.065 2289.370 1771.395 2289.385 ;
        RECT 1755.835 2289.070 1771.395 2289.370 ;
        RECT 1755.835 2288.775 1759.835 2289.070 ;
        RECT 1771.065 2289.055 1771.395 2289.070 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1202.970 2376.160 1203.290 2376.220 ;
        RECT 2111.470 2376.160 2111.790 2376.220 ;
        RECT 1202.970 2376.020 2111.790 2376.160 ;
        RECT 1202.970 2375.960 1203.290 2376.020 ;
        RECT 2111.470 2375.960 2111.790 2376.020 ;
      LAYER via ;
        RECT 1203.000 2375.960 1203.260 2376.220 ;
        RECT 2111.500 2375.960 2111.760 2376.220 ;
      LAYER met2 ;
        RECT 1201.660 2376.330 1201.940 2377.880 ;
        RECT 1201.660 2376.250 1203.200 2376.330 ;
        RECT 1201.660 2376.190 1203.260 2376.250 ;
        RECT 1201.660 2373.880 1201.940 2376.190 ;
        RECT 1203.000 2375.930 1203.260 2376.190 ;
        RECT 2111.500 2375.930 2111.760 2376.250 ;
        RECT 2111.560 16.730 2111.700 2375.930 ;
        RECT 2111.560 16.590 2114.000 16.730 ;
        RECT 2113.860 2.400 2114.000 16.590 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 765.050 51.580 765.370 51.640 ;
        RECT 2125.730 51.580 2126.050 51.640 ;
        RECT 765.050 51.440 2126.050 51.580 ;
        RECT 765.050 51.380 765.370 51.440 ;
        RECT 2125.730 51.380 2126.050 51.440 ;
        RECT 2125.730 19.960 2126.050 20.020 ;
        RECT 2131.710 19.960 2132.030 20.020 ;
        RECT 2125.730 19.820 2132.030 19.960 ;
        RECT 2125.730 19.760 2126.050 19.820 ;
        RECT 2131.710 19.760 2132.030 19.820 ;
      LAYER via ;
        RECT 765.080 51.380 765.340 51.640 ;
        RECT 2125.760 51.380 2126.020 51.640 ;
        RECT 2125.760 19.760 2126.020 20.020 ;
        RECT 2131.740 19.760 2132.000 20.020 ;
      LAYER met2 ;
        RECT 764.660 1323.690 764.940 1327.135 ;
        RECT 764.660 1323.550 765.280 1323.690 ;
        RECT 764.660 1323.135 764.940 1323.550 ;
        RECT 765.140 51.670 765.280 1323.550 ;
        RECT 765.080 51.350 765.340 51.670 ;
        RECT 2125.760 51.350 2126.020 51.670 ;
        RECT 2125.820 20.050 2125.960 51.350 ;
        RECT 2125.760 19.730 2126.020 20.050 ;
        RECT 2131.740 19.730 2132.000 20.050 ;
        RECT 2131.800 2.400 2131.940 19.730 ;
        RECT 2131.590 -4.800 2132.150 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1310.610 52.940 1310.930 53.000 ;
        RECT 2145.970 52.940 2146.290 53.000 ;
        RECT 1310.610 52.800 2146.290 52.940 ;
        RECT 1310.610 52.740 1310.930 52.800 ;
        RECT 2145.970 52.740 2146.290 52.800 ;
      LAYER via ;
        RECT 1310.640 52.740 1310.900 53.000 ;
        RECT 2146.000 52.740 2146.260 53.000 ;
      LAYER met2 ;
        RECT 1308.380 1323.690 1308.660 1327.135 ;
        RECT 1308.380 1323.550 1310.840 1323.690 ;
        RECT 1308.380 1323.135 1308.660 1323.550 ;
        RECT 1310.700 53.030 1310.840 1323.550 ;
        RECT 1310.640 52.710 1310.900 53.030 ;
        RECT 2146.000 52.710 2146.260 53.030 ;
        RECT 2146.060 16.730 2146.200 52.710 ;
        RECT 2146.060 16.590 2149.880 16.730 ;
        RECT 2149.740 2.400 2149.880 16.590 ;
        RECT 2149.530 -4.800 2150.090 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1151.985 15.725 1152.155 18.275 ;
      LAYER mcon ;
        RECT 1151.985 18.105 1152.155 18.275 ;
      LAYER met1 ;
        RECT 1151.925 18.260 1152.215 18.305 ;
        RECT 2167.590 18.260 2167.910 18.320 ;
        RECT 1151.925 18.120 2167.910 18.260 ;
        RECT 1151.925 18.075 1152.215 18.120 ;
        RECT 2167.590 18.060 2167.910 18.120 ;
        RECT 1104.070 15.880 1104.390 15.940 ;
        RECT 1151.925 15.880 1152.215 15.925 ;
        RECT 1104.070 15.740 1152.215 15.880 ;
        RECT 1104.070 15.680 1104.390 15.740 ;
        RECT 1151.925 15.695 1152.215 15.740 ;
      LAYER via ;
        RECT 2167.620 18.060 2167.880 18.320 ;
        RECT 1104.100 15.680 1104.360 15.940 ;
      LAYER met2 ;
        RECT 1104.090 32.115 1104.370 32.485 ;
        RECT 1104.160 15.970 1104.300 32.115 ;
        RECT 2167.620 18.030 2167.880 18.350 ;
        RECT 1104.100 15.650 1104.360 15.970 ;
        RECT 2167.680 2.400 2167.820 18.030 ;
        RECT 2167.470 -4.800 2168.030 2.400 ;
      LAYER via2 ;
        RECT 1104.090 32.160 1104.370 32.440 ;
      LAYER met3 ;
        RECT 709.590 2267.610 709.970 2267.620 ;
        RECT 715.810 2267.610 719.810 2267.615 ;
        RECT 709.590 2267.310 719.810 2267.610 ;
        RECT 709.590 2267.300 709.970 2267.310 ;
        RECT 715.810 2267.015 719.810 2267.310 ;
        RECT 709.590 32.450 709.970 32.460 ;
        RECT 1104.065 32.450 1104.395 32.465 ;
        RECT 709.590 32.150 1104.395 32.450 ;
        RECT 709.590 32.140 709.970 32.150 ;
        RECT 1104.065 32.135 1104.395 32.150 ;
      LAYER via3 ;
        RECT 709.620 2267.300 709.940 2267.620 ;
        RECT 709.620 32.140 709.940 32.460 ;
      LAYER met4 ;
        RECT 709.615 2267.295 709.945 2267.625 ;
        RECT 709.630 32.465 709.930 2267.295 ;
        RECT 709.615 32.135 709.945 32.465 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 713.530 431.360 713.850 431.420 ;
        RECT 2180.470 431.360 2180.790 431.420 ;
        RECT 713.530 431.220 2180.790 431.360 ;
        RECT 713.530 431.160 713.850 431.220 ;
        RECT 2180.470 431.160 2180.790 431.220 ;
      LAYER via ;
        RECT 713.560 431.160 713.820 431.420 ;
        RECT 2180.500 431.160 2180.760 431.420 ;
      LAYER met2 ;
        RECT 713.550 1626.715 713.830 1627.085 ;
        RECT 713.620 431.450 713.760 1626.715 ;
        RECT 713.560 431.130 713.820 431.450 ;
        RECT 2180.500 431.130 2180.760 431.450 ;
        RECT 2180.560 24.210 2180.700 431.130 ;
        RECT 2180.560 24.070 2185.300 24.210 ;
        RECT 2185.160 2.400 2185.300 24.070 ;
        RECT 2184.950 -4.800 2185.510 2.400 ;
      LAYER via2 ;
        RECT 713.550 1626.760 713.830 1627.040 ;
      LAYER met3 ;
        RECT 713.525 1627.050 713.855 1627.065 ;
        RECT 715.810 1627.050 719.810 1627.055 ;
        RECT 713.525 1626.750 719.810 1627.050 ;
        RECT 713.525 1626.735 713.855 1626.750 ;
        RECT 715.810 1626.455 719.810 1626.750 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1517.610 62.120 1517.930 62.180 ;
        RECT 2201.170 62.120 2201.490 62.180 ;
        RECT 1517.610 61.980 2201.490 62.120 ;
        RECT 1517.610 61.920 1517.930 61.980 ;
        RECT 2201.170 61.920 2201.490 61.980 ;
      LAYER via ;
        RECT 1517.640 61.920 1517.900 62.180 ;
        RECT 2201.200 61.920 2201.460 62.180 ;
      LAYER met2 ;
        RECT 1516.300 1323.690 1516.580 1327.135 ;
        RECT 1516.300 1323.550 1517.840 1323.690 ;
        RECT 1516.300 1323.135 1516.580 1323.550 ;
        RECT 1517.700 62.210 1517.840 1323.550 ;
        RECT 1517.640 61.890 1517.900 62.210 ;
        RECT 2201.200 61.890 2201.460 62.210 ;
        RECT 2201.260 24.210 2201.400 61.890 ;
        RECT 2201.260 24.070 2203.240 24.210 ;
        RECT 2203.100 2.400 2203.240 24.070 ;
        RECT 2202.890 -4.800 2203.450 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1346.105 2374.645 1346.735 2374.815 ;
      LAYER mcon ;
        RECT 1346.565 2374.645 1346.735 2374.815 ;
      LAYER met1 ;
        RECT 988.610 2374.800 988.930 2374.860 ;
        RECT 1346.045 2374.800 1346.335 2374.845 ;
        RECT 988.610 2374.660 1346.335 2374.800 ;
        RECT 988.610 2374.600 988.930 2374.660 ;
        RECT 1346.045 2374.615 1346.335 2374.660 ;
        RECT 1346.505 2374.800 1346.795 2374.845 ;
        RECT 2215.430 2374.800 2215.750 2374.860 ;
        RECT 1346.505 2374.660 2215.750 2374.800 ;
        RECT 1346.505 2374.615 1346.795 2374.660 ;
        RECT 2215.430 2374.600 2215.750 2374.660 ;
      LAYER via ;
        RECT 988.640 2374.600 988.900 2374.860 ;
        RECT 2215.460 2374.600 2215.720 2374.860 ;
      LAYER met2 ;
        RECT 987.300 2374.970 987.580 2377.880 ;
        RECT 987.300 2374.890 988.840 2374.970 ;
        RECT 987.300 2374.830 988.900 2374.890 ;
        RECT 987.300 2373.880 987.580 2374.830 ;
        RECT 988.640 2374.570 988.900 2374.830 ;
        RECT 2215.460 2374.570 2215.720 2374.890 ;
        RECT 2215.520 16.730 2215.660 2374.570 ;
        RECT 2215.520 16.590 2221.180 16.730 ;
        RECT 2221.040 2.400 2221.180 16.590 ;
        RECT 2220.830 -4.800 2221.390 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 775.630 52.600 775.950 52.660 ;
        RECT 1677.230 52.600 1677.550 52.660 ;
        RECT 775.630 52.460 1677.550 52.600 ;
        RECT 775.630 52.400 775.950 52.460 ;
        RECT 1677.230 52.400 1677.550 52.460 ;
      LAYER via ;
        RECT 775.660 52.400 775.920 52.660 ;
        RECT 1677.260 52.400 1677.520 52.660 ;
      LAYER met2 ;
        RECT 1678.220 1323.690 1678.500 1327.135 ;
        RECT 1677.320 1323.550 1678.500 1323.690 ;
        RECT 1677.320 52.690 1677.460 1323.550 ;
        RECT 1678.220 1323.135 1678.500 1323.550 ;
        RECT 775.660 52.370 775.920 52.690 ;
        RECT 1677.260 52.370 1677.520 52.690 ;
        RECT 775.720 2.400 775.860 52.370 ;
        RECT 775.510 -4.800 776.070 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1345.645 2374.985 1347.195 2375.155 ;
      LAYER mcon ;
        RECT 1347.025 2374.985 1347.195 2375.155 ;
      LAYER met1 ;
        RECT 1116.490 2375.140 1116.810 2375.200 ;
        RECT 1345.585 2375.140 1345.875 2375.185 ;
        RECT 1116.490 2375.000 1345.875 2375.140 ;
        RECT 1116.490 2374.940 1116.810 2375.000 ;
        RECT 1345.585 2374.955 1345.875 2375.000 ;
        RECT 1346.965 2375.140 1347.255 2375.185 ;
        RECT 2235.670 2375.140 2235.990 2375.200 ;
        RECT 1346.965 2375.000 2235.990 2375.140 ;
        RECT 1346.965 2374.955 1347.255 2375.000 ;
        RECT 2235.670 2374.940 2235.990 2375.000 ;
      LAYER via ;
        RECT 1116.520 2374.940 1116.780 2375.200 ;
        RECT 2235.700 2374.940 2235.960 2375.200 ;
      LAYER met2 ;
        RECT 1115.180 2374.970 1115.460 2377.880 ;
        RECT 1116.520 2374.970 1116.780 2375.230 ;
        RECT 1115.180 2374.910 1116.780 2374.970 ;
        RECT 2235.700 2374.910 2235.960 2375.230 ;
        RECT 1115.180 2374.830 1116.720 2374.910 ;
        RECT 1115.180 2373.880 1115.460 2374.830 ;
        RECT 2235.760 16.730 2235.900 2374.910 ;
        RECT 2235.760 16.590 2239.120 16.730 ;
        RECT 2238.980 2.400 2239.120 16.590 ;
        RECT 2238.770 -4.800 2239.330 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1595.810 2376.500 1596.130 2376.560 ;
        RECT 2256.370 2376.500 2256.690 2376.560 ;
        RECT 1595.810 2376.360 2256.690 2376.500 ;
        RECT 1595.810 2376.300 1596.130 2376.360 ;
        RECT 2256.370 2376.300 2256.690 2376.360 ;
      LAYER via ;
        RECT 1595.840 2376.300 1596.100 2376.560 ;
        RECT 2256.400 2376.300 2256.660 2376.560 ;
      LAYER met2 ;
        RECT 1594.500 2376.330 1594.780 2377.880 ;
        RECT 1595.840 2376.330 1596.100 2376.590 ;
        RECT 1594.500 2376.270 1596.100 2376.330 ;
        RECT 2256.400 2376.270 2256.660 2376.590 ;
        RECT 1594.500 2376.190 1596.040 2376.270 ;
        RECT 1594.500 2373.880 1594.780 2376.190 ;
        RECT 2256.460 2.400 2256.600 2376.270 ;
        RECT 2256.250 -4.800 2256.810 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1147.770 18.260 1148.090 18.320 ;
        RECT 1151.450 18.260 1151.770 18.320 ;
        RECT 1147.770 18.120 1151.770 18.260 ;
        RECT 1147.770 18.060 1148.090 18.120 ;
        RECT 1151.450 18.060 1151.770 18.120 ;
      LAYER via ;
        RECT 1147.800 18.060 1148.060 18.320 ;
        RECT 1151.480 18.060 1151.740 18.320 ;
      LAYER met2 ;
        RECT 701.130 1591.355 701.410 1591.725 ;
        RECT 701.200 1393.845 701.340 1591.355 ;
        RECT 701.130 1393.475 701.410 1393.845 ;
        RECT 701.130 1390.755 701.410 1391.125 ;
        RECT 701.200 18.885 701.340 1390.755 ;
        RECT 701.130 18.515 701.410 18.885 ;
        RECT 1147.790 18.515 1148.070 18.885 ;
        RECT 1151.470 18.515 1151.750 18.885 ;
        RECT 1454.610 18.515 1454.890 18.885 ;
        RECT 1496.470 18.515 1496.750 18.885 ;
        RECT 2274.330 18.515 2274.610 18.885 ;
        RECT 1147.860 18.350 1148.000 18.515 ;
        RECT 1151.540 18.350 1151.680 18.515 ;
        RECT 1147.800 18.030 1148.060 18.350 ;
        RECT 1151.480 18.030 1151.740 18.350 ;
        RECT 1454.680 16.165 1454.820 18.515 ;
        RECT 1496.540 16.165 1496.680 18.515 ;
        RECT 1454.610 15.795 1454.890 16.165 ;
        RECT 1496.470 15.795 1496.750 16.165 ;
        RECT 2274.400 2.400 2274.540 18.515 ;
        RECT 2274.190 -4.800 2274.750 2.400 ;
      LAYER via2 ;
        RECT 701.130 1591.400 701.410 1591.680 ;
        RECT 701.130 1393.520 701.410 1393.800 ;
        RECT 701.130 1390.800 701.410 1391.080 ;
        RECT 701.130 18.560 701.410 18.840 ;
        RECT 1147.790 18.560 1148.070 18.840 ;
        RECT 1151.470 18.560 1151.750 18.840 ;
        RECT 1454.610 18.560 1454.890 18.840 ;
        RECT 1496.470 18.560 1496.750 18.840 ;
        RECT 2274.330 18.560 2274.610 18.840 ;
        RECT 1454.610 15.840 1454.890 16.120 ;
        RECT 1496.470 15.840 1496.750 16.120 ;
      LAYER met3 ;
        RECT 701.105 1591.690 701.435 1591.705 ;
        RECT 715.810 1591.690 719.810 1591.695 ;
        RECT 701.105 1591.390 719.810 1591.690 ;
        RECT 701.105 1591.375 701.435 1591.390 ;
        RECT 715.810 1591.095 719.810 1591.390 ;
        RECT 701.105 1393.810 701.435 1393.825 ;
        RECT 701.105 1393.495 701.650 1393.810 ;
        RECT 701.350 1391.105 701.650 1393.495 ;
        RECT 701.105 1390.790 701.650 1391.105 ;
        RECT 701.105 1390.775 701.435 1390.790 ;
        RECT 701.105 18.850 701.435 18.865 ;
        RECT 1147.765 18.850 1148.095 18.865 ;
        RECT 701.105 18.550 1148.095 18.850 ;
        RECT 701.105 18.535 701.435 18.550 ;
        RECT 1147.765 18.535 1148.095 18.550 ;
        RECT 1151.445 18.850 1151.775 18.865 ;
        RECT 1454.585 18.850 1454.915 18.865 ;
        RECT 1151.445 18.550 1454.915 18.850 ;
        RECT 1151.445 18.535 1151.775 18.550 ;
        RECT 1454.585 18.535 1454.915 18.550 ;
        RECT 1496.445 18.850 1496.775 18.865 ;
        RECT 2274.305 18.850 2274.635 18.865 ;
        RECT 1496.445 18.550 2274.635 18.850 ;
        RECT 1496.445 18.535 1496.775 18.550 ;
        RECT 2274.305 18.535 2274.635 18.550 ;
        RECT 1454.585 16.130 1454.915 16.145 ;
        RECT 1496.445 16.130 1496.775 16.145 ;
        RECT 1454.585 15.830 1496.775 16.130 ;
        RECT 1454.585 15.815 1454.915 15.830 ;
        RECT 1496.445 15.815 1496.775 15.830 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2290.890 888.235 2291.170 888.605 ;
        RECT 2290.960 24.210 2291.100 888.235 ;
        RECT 2290.960 24.070 2292.480 24.210 ;
        RECT 2292.340 2.400 2292.480 24.070 ;
        RECT 2292.130 -4.800 2292.690 2.400 ;
      LAYER via2 ;
        RECT 2290.890 888.280 2291.170 888.560 ;
      LAYER met3 ;
        RECT 706.830 1892.250 707.210 1892.260 ;
        RECT 715.810 1892.250 719.810 1892.255 ;
        RECT 706.830 1891.950 719.810 1892.250 ;
        RECT 706.830 1891.940 707.210 1891.950 ;
        RECT 715.810 1891.655 719.810 1891.950 ;
        RECT 706.830 888.570 707.210 888.580 ;
        RECT 2290.865 888.570 2291.195 888.585 ;
        RECT 706.830 888.270 2291.195 888.570 ;
        RECT 706.830 888.260 707.210 888.270 ;
        RECT 2290.865 888.255 2291.195 888.270 ;
      LAYER via3 ;
        RECT 706.860 1891.940 707.180 1892.260 ;
        RECT 706.860 888.260 707.180 888.580 ;
      LAYER met4 ;
        RECT 706.855 1891.935 707.185 1892.265 ;
        RECT 706.870 888.585 707.170 1891.935 ;
        RECT 706.855 888.255 707.185 888.585 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1124.310 61.100 1124.630 61.160 ;
        RECT 2304.670 61.100 2304.990 61.160 ;
        RECT 1124.310 60.960 2304.990 61.100 ;
        RECT 1124.310 60.900 1124.630 60.960 ;
        RECT 2304.670 60.900 2304.990 60.960 ;
      LAYER via ;
        RECT 1124.340 60.900 1124.600 61.160 ;
        RECT 2304.700 60.900 2304.960 61.160 ;
      LAYER met2 ;
        RECT 1123.460 1323.690 1123.740 1327.135 ;
        RECT 1123.460 1323.550 1124.540 1323.690 ;
        RECT 1123.460 1323.135 1123.740 1323.550 ;
        RECT 1124.400 61.190 1124.540 1323.550 ;
        RECT 1124.340 60.870 1124.600 61.190 ;
        RECT 2304.700 60.870 2304.960 61.190 ;
        RECT 2304.760 16.730 2304.900 60.870 ;
        RECT 2304.760 16.590 2310.420 16.730 ;
        RECT 2310.280 2.400 2310.420 16.590 ;
        RECT 2310.070 -4.800 2310.630 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 929.270 2379.900 929.590 2379.960 ;
        RECT 2325.370 2379.900 2325.690 2379.960 ;
        RECT 929.270 2379.760 2325.690 2379.900 ;
        RECT 929.270 2379.700 929.590 2379.760 ;
        RECT 2325.370 2379.700 2325.690 2379.760 ;
      LAYER via ;
        RECT 929.300 2379.700 929.560 2379.960 ;
        RECT 2325.400 2379.700 2325.660 2379.960 ;
      LAYER met2 ;
        RECT 929.300 2379.670 929.560 2379.990 ;
        RECT 2325.400 2379.670 2325.660 2379.990 ;
        RECT 929.360 2377.880 929.500 2379.670 ;
        RECT 929.340 2373.880 929.620 2377.880 ;
        RECT 2325.460 16.730 2325.600 2379.670 ;
        RECT 2325.460 16.590 2328.360 16.730 ;
        RECT 2328.220 2.400 2328.360 16.590 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1772.910 1504.400 1773.230 1504.460 ;
        RECT 2339.630 1504.400 2339.950 1504.460 ;
        RECT 1772.910 1504.260 2339.950 1504.400 ;
        RECT 1772.910 1504.200 1773.230 1504.260 ;
        RECT 2339.630 1504.200 2339.950 1504.260 ;
        RECT 2339.630 38.320 2339.950 38.380 ;
        RECT 2345.610 38.320 2345.930 38.380 ;
        RECT 2339.630 38.180 2345.930 38.320 ;
        RECT 2339.630 38.120 2339.950 38.180 ;
        RECT 2345.610 38.120 2345.930 38.180 ;
      LAYER via ;
        RECT 1772.940 1504.200 1773.200 1504.460 ;
        RECT 2339.660 1504.200 2339.920 1504.460 ;
        RECT 2339.660 38.120 2339.920 38.380 ;
        RECT 2345.640 38.120 2345.900 38.380 ;
      LAYER met2 ;
        RECT 1772.930 1509.755 1773.210 1510.125 ;
        RECT 1773.000 1504.490 1773.140 1509.755 ;
        RECT 1772.940 1504.170 1773.200 1504.490 ;
        RECT 2339.660 1504.170 2339.920 1504.490 ;
        RECT 2339.720 38.410 2339.860 1504.170 ;
        RECT 2339.660 38.090 2339.920 38.410 ;
        RECT 2345.640 38.090 2345.900 38.410 ;
        RECT 2345.700 2.400 2345.840 38.090 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
      LAYER via2 ;
        RECT 1772.930 1509.800 1773.210 1510.080 ;
      LAYER met3 ;
        RECT 1755.835 1510.090 1759.835 1510.095 ;
        RECT 1772.905 1510.090 1773.235 1510.105 ;
        RECT 1755.835 1509.790 1773.235 1510.090 ;
        RECT 1755.835 1509.495 1759.835 1509.790 ;
        RECT 1772.905 1509.775 1773.235 1509.790 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2363.625 2.805 2363.795 16.915 ;
      LAYER mcon ;
        RECT 2363.625 16.745 2363.795 16.915 ;
      LAYER met1 ;
        RECT 2359.870 16.900 2360.190 16.960 ;
        RECT 2363.565 16.900 2363.855 16.945 ;
        RECT 2359.870 16.760 2363.855 16.900 ;
        RECT 2359.870 16.700 2360.190 16.760 ;
        RECT 2363.565 16.715 2363.855 16.760 ;
        RECT 2363.550 2.960 2363.870 3.020 ;
        RECT 2363.355 2.820 2363.870 2.960 ;
        RECT 2363.550 2.760 2363.870 2.820 ;
      LAYER via ;
        RECT 2359.900 16.700 2360.160 16.960 ;
        RECT 2363.580 2.760 2363.840 3.020 ;
      LAYER met2 ;
        RECT 2359.890 1307.795 2360.170 1308.165 ;
        RECT 2359.960 16.990 2360.100 1307.795 ;
        RECT 2359.900 16.670 2360.160 16.990 ;
        RECT 2363.580 2.730 2363.840 3.050 ;
        RECT 2363.640 2.400 2363.780 2.730 ;
        RECT 2363.430 -4.800 2363.990 2.400 ;
      LAYER via2 ;
        RECT 2359.890 1307.840 2360.170 1308.120 ;
      LAYER met3 ;
        RECT 713.270 2181.930 713.650 2181.940 ;
        RECT 715.810 2181.930 719.810 2181.935 ;
        RECT 713.270 2181.630 719.810 2181.930 ;
        RECT 713.270 2181.620 713.650 2181.630 ;
        RECT 715.810 2181.335 719.810 2181.630 ;
        RECT 713.270 1309.490 713.650 1309.500 ;
        RECT 713.270 1309.190 731.090 1309.490 ;
        RECT 713.270 1309.180 713.650 1309.190 ;
        RECT 730.790 1308.130 731.090 1309.190 ;
        RECT 2359.865 1308.130 2360.195 1308.145 ;
        RECT 730.790 1307.830 2360.195 1308.130 ;
        RECT 2359.865 1307.815 2360.195 1307.830 ;
      LAYER via3 ;
        RECT 713.300 2181.620 713.620 2181.940 ;
        RECT 713.300 1309.180 713.620 1309.500 ;
      LAYER met4 ;
        RECT 713.295 2181.615 713.625 2181.945 ;
        RECT 713.310 1309.505 713.610 2181.615 ;
        RECT 713.295 1309.175 713.625 1309.505 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1424.230 1311.280 1424.550 1311.340 ;
        RECT 1427.910 1311.280 1428.230 1311.340 ;
        RECT 1424.230 1311.140 1428.230 1311.280 ;
        RECT 1424.230 1311.080 1424.550 1311.140 ;
        RECT 1427.910 1311.080 1428.230 1311.140 ;
        RECT 1427.910 61.780 1428.230 61.840 ;
        RECT 2381.490 61.780 2381.810 61.840 ;
        RECT 1427.910 61.640 2381.810 61.780 ;
        RECT 1427.910 61.580 1428.230 61.640 ;
        RECT 2381.490 61.580 2381.810 61.640 ;
      LAYER via ;
        RECT 1424.260 1311.080 1424.520 1311.340 ;
        RECT 1427.940 1311.080 1428.200 1311.340 ;
        RECT 1427.940 61.580 1428.200 61.840 ;
        RECT 2381.520 61.580 2381.780 61.840 ;
      LAYER met2 ;
        RECT 1424.300 1323.135 1424.580 1327.135 ;
        RECT 1424.320 1311.370 1424.460 1323.135 ;
        RECT 1424.260 1311.050 1424.520 1311.370 ;
        RECT 1427.940 1311.050 1428.200 1311.370 ;
        RECT 1428.000 61.870 1428.140 1311.050 ;
        RECT 1427.940 61.550 1428.200 61.870 ;
        RECT 2381.520 61.550 2381.780 61.870 ;
        RECT 2381.580 2.400 2381.720 61.550 ;
        RECT 2381.370 -4.800 2381.930 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1772.910 1960.000 1773.230 1960.060 ;
        RECT 2394.370 1960.000 2394.690 1960.060 ;
        RECT 1772.910 1959.860 2394.690 1960.000 ;
        RECT 1772.910 1959.800 1773.230 1959.860 ;
        RECT 2394.370 1959.800 2394.690 1959.860 ;
        RECT 2394.370 62.120 2394.690 62.180 ;
        RECT 2399.430 62.120 2399.750 62.180 ;
        RECT 2394.370 61.980 2399.750 62.120 ;
        RECT 2394.370 61.920 2394.690 61.980 ;
        RECT 2399.430 61.920 2399.750 61.980 ;
      LAYER via ;
        RECT 1772.940 1959.800 1773.200 1960.060 ;
        RECT 2394.400 1959.800 2394.660 1960.060 ;
        RECT 2394.400 61.920 2394.660 62.180 ;
        RECT 2399.460 61.920 2399.720 62.180 ;
      LAYER met2 ;
        RECT 1772.930 1963.995 1773.210 1964.365 ;
        RECT 1773.000 1960.090 1773.140 1963.995 ;
        RECT 1772.940 1959.770 1773.200 1960.090 ;
        RECT 2394.400 1959.770 2394.660 1960.090 ;
        RECT 2394.460 62.210 2394.600 1959.770 ;
        RECT 2394.400 61.890 2394.660 62.210 ;
        RECT 2399.460 61.890 2399.720 62.210 ;
        RECT 2399.520 2.400 2399.660 61.890 ;
        RECT 2399.310 -4.800 2399.870 2.400 ;
      LAYER via2 ;
        RECT 1772.930 1964.040 1773.210 1964.320 ;
      LAYER met3 ;
        RECT 1755.835 1964.330 1759.835 1964.335 ;
        RECT 1772.905 1964.330 1773.235 1964.345 ;
        RECT 1755.835 1964.030 1773.235 1964.330 ;
        RECT 1755.835 1963.735 1759.835 1964.030 ;
        RECT 1772.905 1964.015 1773.235 1964.030 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 688.765 1368.925 688.935 1393.575 ;
      LAYER mcon ;
        RECT 688.765 1393.405 688.935 1393.575 ;
      LAYER met1 ;
        RECT 688.690 1932.120 689.010 1932.180 ;
        RECT 704.330 1932.120 704.650 1932.180 ;
        RECT 688.690 1931.980 704.650 1932.120 ;
        RECT 688.690 1931.920 689.010 1931.980 ;
        RECT 704.330 1931.920 704.650 1931.980 ;
        RECT 688.690 1393.560 689.010 1393.620 ;
        RECT 688.690 1393.420 689.205 1393.560 ;
        RECT 688.690 1393.360 689.010 1393.420 ;
        RECT 688.690 1369.080 689.010 1369.140 ;
        RECT 688.495 1368.940 689.010 1369.080 ;
        RECT 688.690 1368.880 689.010 1368.940 ;
        RECT 688.690 14.860 689.010 14.920 ;
        RECT 793.570 14.860 793.890 14.920 ;
        RECT 688.690 14.720 793.890 14.860 ;
        RECT 688.690 14.660 689.010 14.720 ;
        RECT 793.570 14.660 793.890 14.720 ;
      LAYER via ;
        RECT 688.720 1931.920 688.980 1932.180 ;
        RECT 704.360 1931.920 704.620 1932.180 ;
        RECT 688.720 1393.360 688.980 1393.620 ;
        RECT 688.720 1368.880 688.980 1369.140 ;
        RECT 688.720 14.660 688.980 14.920 ;
        RECT 793.600 14.660 793.860 14.920 ;
      LAYER met2 ;
        RECT 704.350 1934.075 704.630 1934.445 ;
        RECT 704.420 1932.210 704.560 1934.075 ;
        RECT 688.720 1931.890 688.980 1932.210 ;
        RECT 704.360 1931.890 704.620 1932.210 ;
        RECT 688.780 1393.650 688.920 1931.890 ;
        RECT 688.720 1393.330 688.980 1393.650 ;
        RECT 688.720 1368.850 688.980 1369.170 ;
        RECT 688.780 14.950 688.920 1368.850 ;
        RECT 688.720 14.630 688.980 14.950 ;
        RECT 793.600 14.630 793.860 14.950 ;
        RECT 793.660 2.400 793.800 14.630 ;
        RECT 793.450 -4.800 794.010 2.400 ;
      LAYER via2 ;
        RECT 704.350 1934.120 704.630 1934.400 ;
      LAYER met3 ;
        RECT 704.325 1934.410 704.655 1934.425 ;
        RECT 715.810 1934.410 719.810 1934.415 ;
        RECT 704.325 1934.110 719.810 1934.410 ;
        RECT 704.325 1934.095 704.655 1934.110 ;
        RECT 715.810 1933.815 719.810 1934.110 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 641.310 52.940 641.630 53.000 ;
        RECT 1200.670 52.940 1200.990 53.000 ;
        RECT 641.310 52.800 1200.990 52.940 ;
        RECT 641.310 52.740 641.630 52.800 ;
        RECT 1200.670 52.740 1200.990 52.800 ;
        RECT 639.010 17.240 639.330 17.300 ;
        RECT 641.310 17.240 641.630 17.300 ;
        RECT 639.010 17.100 641.630 17.240 ;
        RECT 639.010 17.040 639.330 17.100 ;
        RECT 641.310 17.040 641.630 17.100 ;
      LAYER via ;
        RECT 641.340 52.740 641.600 53.000 ;
        RECT 1200.700 52.740 1200.960 53.000 ;
        RECT 639.040 17.040 639.300 17.300 ;
        RECT 641.340 17.040 641.600 17.300 ;
      LAYER met2 ;
        RECT 1204.420 1323.690 1204.700 1327.135 ;
        RECT 1200.760 1323.550 1204.700 1323.690 ;
        RECT 1200.760 53.030 1200.900 1323.550 ;
        RECT 1204.420 1323.135 1204.700 1323.550 ;
        RECT 641.340 52.710 641.600 53.030 ;
        RECT 1200.700 52.710 1200.960 53.030 ;
        RECT 641.400 17.330 641.540 52.710 ;
        RECT 639.040 17.010 639.300 17.330 ;
        RECT 641.340 17.010 641.600 17.330 ;
        RECT 639.100 2.400 639.240 17.010 ;
        RECT 638.890 -4.800 639.450 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1644.110 1311.280 1644.430 1311.340 ;
        RECT 1648.710 1311.280 1649.030 1311.340 ;
        RECT 1644.110 1311.140 1649.030 1311.280 ;
        RECT 1644.110 1311.080 1644.430 1311.140 ;
        RECT 1648.710 1311.080 1649.030 1311.140 ;
        RECT 1648.710 24.380 1649.030 24.440 ;
        RECT 2422.890 24.380 2423.210 24.440 ;
        RECT 1648.710 24.240 2423.210 24.380 ;
        RECT 1648.710 24.180 1649.030 24.240 ;
        RECT 2422.890 24.180 2423.210 24.240 ;
      LAYER via ;
        RECT 1644.140 1311.080 1644.400 1311.340 ;
        RECT 1648.740 1311.080 1649.000 1311.340 ;
        RECT 1648.740 24.180 1649.000 24.440 ;
        RECT 2422.920 24.180 2423.180 24.440 ;
      LAYER met2 ;
        RECT 1644.180 1323.135 1644.460 1327.135 ;
        RECT 1644.200 1311.370 1644.340 1323.135 ;
        RECT 1644.140 1311.050 1644.400 1311.370 ;
        RECT 1648.740 1311.050 1649.000 1311.370 ;
        RECT 1648.800 24.470 1648.940 1311.050 ;
        RECT 1648.740 24.150 1649.000 24.470 ;
        RECT 2422.920 24.150 2423.180 24.470 ;
        RECT 2422.980 2.400 2423.120 24.150 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1752.285 52.445 1752.455 89.335 ;
      LAYER mcon ;
        RECT 1752.285 89.165 1752.455 89.335 ;
      LAYER met1 ;
        RECT 1748.070 1311.620 1748.390 1311.680 ;
        RECT 1752.210 1311.620 1752.530 1311.680 ;
        RECT 1748.070 1311.480 1752.530 1311.620 ;
        RECT 1748.070 1311.420 1748.390 1311.480 ;
        RECT 1752.210 1311.420 1752.530 1311.480 ;
        RECT 1752.210 89.320 1752.530 89.380 ;
        RECT 1752.015 89.180 1752.530 89.320 ;
        RECT 1752.210 89.120 1752.530 89.180 ;
        RECT 1752.225 52.600 1752.515 52.645 ;
        RECT 2440.830 52.600 2441.150 52.660 ;
        RECT 1752.225 52.460 2441.150 52.600 ;
        RECT 1752.225 52.415 1752.515 52.460 ;
        RECT 2440.830 52.400 2441.150 52.460 ;
      LAYER via ;
        RECT 1748.100 1311.420 1748.360 1311.680 ;
        RECT 1752.240 1311.420 1752.500 1311.680 ;
        RECT 1752.240 89.120 1752.500 89.380 ;
        RECT 2440.860 52.400 2441.120 52.660 ;
      LAYER met2 ;
        RECT 1748.140 1323.135 1748.420 1327.135 ;
        RECT 1748.160 1311.710 1748.300 1323.135 ;
        RECT 1748.100 1311.390 1748.360 1311.710 ;
        RECT 1752.240 1311.390 1752.500 1311.710 ;
        RECT 1752.300 89.410 1752.440 1311.390 ;
        RECT 1752.240 89.090 1752.500 89.410 ;
        RECT 2440.860 52.370 2441.120 52.690 ;
        RECT 2440.920 2.400 2441.060 52.370 ;
        RECT 2440.710 -4.800 2441.270 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 848.310 59.740 848.630 59.800 ;
        RECT 2458.770 59.740 2459.090 59.800 ;
        RECT 848.310 59.600 2459.090 59.740 ;
        RECT 848.310 59.540 848.630 59.600 ;
        RECT 2458.770 59.540 2459.090 59.600 ;
      LAYER via ;
        RECT 848.340 59.540 848.600 59.800 ;
        RECT 2458.800 59.540 2459.060 59.800 ;
      LAYER met2 ;
        RECT 845.620 1323.690 845.900 1327.135 ;
        RECT 845.620 1323.550 848.540 1323.690 ;
        RECT 845.620 1323.135 845.900 1323.550 ;
        RECT 848.400 59.830 848.540 1323.550 ;
        RECT 848.340 59.510 848.600 59.830 ;
        RECT 2458.800 59.510 2459.060 59.830 ;
        RECT 2458.860 2.400 2459.000 59.510 ;
        RECT 2458.650 -4.800 2459.210 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 772.410 59.400 772.730 59.460 ;
        RECT 2476.710 59.400 2477.030 59.460 ;
        RECT 772.410 59.260 2477.030 59.400 ;
        RECT 772.410 59.200 772.730 59.260 ;
        RECT 2476.710 59.200 2477.030 59.260 ;
      LAYER via ;
        RECT 772.440 59.200 772.700 59.460 ;
        RECT 2476.740 59.200 2477.000 59.460 ;
      LAYER met2 ;
        RECT 770.180 1323.690 770.460 1327.135 ;
        RECT 770.180 1323.550 772.640 1323.690 ;
        RECT 770.180 1323.135 770.460 1323.550 ;
        RECT 772.500 59.490 772.640 1323.550 ;
        RECT 772.440 59.170 772.700 59.490 ;
        RECT 2476.740 59.170 2477.000 59.490 ;
        RECT 2476.800 2.400 2476.940 59.170 ;
        RECT 2476.590 -4.800 2477.150 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1767.850 1808.020 1768.170 1808.080 ;
        RECT 2490.970 1808.020 2491.290 1808.080 ;
        RECT 1767.850 1807.880 2491.290 1808.020 ;
        RECT 1767.850 1807.820 1768.170 1807.880 ;
        RECT 2490.970 1807.820 2491.290 1807.880 ;
      LAYER via ;
        RECT 1767.880 1807.820 1768.140 1808.080 ;
        RECT 2491.000 1807.820 2491.260 1808.080 ;
      LAYER met2 ;
        RECT 1767.870 1808.955 1768.150 1809.325 ;
        RECT 1767.940 1808.110 1768.080 1808.955 ;
        RECT 1767.880 1807.790 1768.140 1808.110 ;
        RECT 2491.000 1807.790 2491.260 1808.110 ;
        RECT 2491.060 24.210 2491.200 1807.790 ;
        RECT 2491.060 24.070 2494.880 24.210 ;
        RECT 2494.740 2.400 2494.880 24.070 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
      LAYER via2 ;
        RECT 1767.870 1809.000 1768.150 1809.280 ;
      LAYER met3 ;
        RECT 1755.835 1809.290 1759.835 1809.295 ;
        RECT 1767.845 1809.290 1768.175 1809.305 ;
        RECT 1755.835 1808.990 1768.175 1809.290 ;
        RECT 1755.835 1808.695 1759.835 1808.990 ;
        RECT 1767.845 1808.975 1768.175 1808.990 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2512.150 17.155 2512.430 17.525 ;
        RECT 2512.220 2.400 2512.360 17.155 ;
        RECT 2512.010 -4.800 2512.570 2.400 ;
      LAYER via2 ;
        RECT 2512.150 17.200 2512.430 17.480 ;
      LAYER met3 ;
        RECT 695.790 1489.690 696.170 1489.700 ;
        RECT 715.810 1489.690 719.810 1489.695 ;
        RECT 695.790 1489.390 719.810 1489.690 ;
        RECT 695.790 1489.380 696.170 1489.390 ;
        RECT 715.810 1489.095 719.810 1489.390 ;
        RECT 695.790 17.490 696.170 17.500 ;
        RECT 2512.125 17.490 2512.455 17.505 ;
        RECT 695.790 17.190 2512.455 17.490 ;
        RECT 695.790 17.180 696.170 17.190 ;
        RECT 2512.125 17.175 2512.455 17.190 ;
      LAYER via3 ;
        RECT 695.820 1489.380 696.140 1489.700 ;
        RECT 695.820 17.180 696.140 17.500 ;
      LAYER met4 ;
        RECT 695.815 1489.375 696.145 1489.705 ;
        RECT 695.830 17.505 696.130 1489.375 ;
        RECT 695.815 17.175 696.145 17.505 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1042.430 1311.280 1042.750 1311.340 ;
        RECT 1047.950 1311.280 1048.270 1311.340 ;
        RECT 1042.430 1311.140 1048.270 1311.280 ;
        RECT 1042.430 1311.080 1042.750 1311.140 ;
        RECT 1047.950 1311.080 1048.270 1311.140 ;
        RECT 1047.950 60.080 1048.270 60.140 ;
        RECT 2530.070 60.080 2530.390 60.140 ;
        RECT 1047.950 59.940 2530.390 60.080 ;
        RECT 1047.950 59.880 1048.270 59.940 ;
        RECT 2530.070 59.880 2530.390 59.940 ;
      LAYER via ;
        RECT 1042.460 1311.080 1042.720 1311.340 ;
        RECT 1047.980 1311.080 1048.240 1311.340 ;
        RECT 1047.980 59.880 1048.240 60.140 ;
        RECT 2530.100 59.880 2530.360 60.140 ;
      LAYER met2 ;
        RECT 1042.500 1323.135 1042.780 1327.135 ;
        RECT 1042.520 1311.370 1042.660 1323.135 ;
        RECT 1042.460 1311.050 1042.720 1311.370 ;
        RECT 1047.980 1311.050 1048.240 1311.370 ;
        RECT 1048.040 60.170 1048.180 1311.050 ;
        RECT 1047.980 59.850 1048.240 60.170 ;
        RECT 2530.100 59.850 2530.360 60.170 ;
        RECT 2530.160 2.400 2530.300 59.850 ;
        RECT 2529.950 -4.800 2530.510 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1691.490 17.580 1691.810 17.640 ;
        RECT 2548.010 17.580 2548.330 17.640 ;
        RECT 1691.490 17.440 2548.330 17.580 ;
        RECT 1691.490 17.380 1691.810 17.440 ;
        RECT 2548.010 17.380 2548.330 17.440 ;
      LAYER via ;
        RECT 1691.520 17.380 1691.780 17.640 ;
        RECT 2548.040 17.380 2548.300 17.640 ;
      LAYER met2 ;
        RECT 1691.510 46.395 1691.790 46.765 ;
        RECT 1691.580 17.670 1691.720 46.395 ;
        RECT 1691.520 17.350 1691.780 17.670 ;
        RECT 2548.040 17.350 2548.300 17.670 ;
        RECT 2548.100 2.400 2548.240 17.350 ;
        RECT 2547.890 -4.800 2548.450 2.400 ;
      LAYER via2 ;
        RECT 1691.510 46.440 1691.790 46.720 ;
      LAYER met3 ;
        RECT 708.670 2275.770 709.050 2275.780 ;
        RECT 715.810 2275.770 719.810 2275.775 ;
        RECT 708.670 2275.470 719.810 2275.770 ;
        RECT 708.670 2275.460 709.050 2275.470 ;
        RECT 715.810 2275.175 719.810 2275.470 ;
        RECT 708.670 46.730 709.050 46.740 ;
        RECT 1691.485 46.730 1691.815 46.745 ;
        RECT 708.670 46.430 1691.815 46.730 ;
        RECT 708.670 46.420 709.050 46.430 ;
        RECT 1691.485 46.415 1691.815 46.430 ;
      LAYER via3 ;
        RECT 708.700 2275.460 709.020 2275.780 ;
        RECT 708.700 46.420 709.020 46.740 ;
      LAYER met4 ;
        RECT 708.695 2275.455 709.025 2275.785 ;
        RECT 708.710 46.745 709.010 2275.455 ;
        RECT 708.695 46.415 709.025 46.745 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2565.970 45.035 2566.250 45.405 ;
        RECT 2566.040 2.400 2566.180 45.035 ;
        RECT 2565.830 -4.800 2566.390 2.400 ;
      LAYER via2 ;
        RECT 2565.970 45.080 2566.250 45.360 ;
      LAYER met3 ;
        RECT 710.510 2241.770 710.890 2241.780 ;
        RECT 715.810 2241.770 719.810 2241.775 ;
        RECT 710.510 2241.470 719.810 2241.770 ;
        RECT 710.510 2241.460 710.890 2241.470 ;
        RECT 715.810 2241.175 719.810 2241.470 ;
        RECT 710.510 45.370 710.890 45.380 ;
        RECT 2565.945 45.370 2566.275 45.385 ;
        RECT 710.510 45.070 2566.275 45.370 ;
        RECT 710.510 45.060 710.890 45.070 ;
        RECT 2565.945 45.055 2566.275 45.070 ;
      LAYER via3 ;
        RECT 710.540 2241.460 710.860 2241.780 ;
        RECT 710.540 45.060 710.860 45.380 ;
      LAYER met4 ;
        RECT 710.535 2241.455 710.865 2241.785 ;
        RECT 710.550 45.385 710.850 2241.455 ;
        RECT 710.535 45.055 710.865 45.385 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 760.065 14.025 760.235 18.275 ;
      LAYER mcon ;
        RECT 760.065 18.105 760.235 18.275 ;
      LAYER met1 ;
        RECT 681.790 2201.400 682.110 2201.460 ;
        RECT 685.470 2201.400 685.790 2201.460 ;
        RECT 681.790 2201.260 685.790 2201.400 ;
        RECT 681.790 2201.200 682.110 2201.260 ;
        RECT 685.470 2201.200 685.790 2201.260 ;
        RECT 758.150 18.260 758.470 18.320 ;
        RECT 760.005 18.260 760.295 18.305 ;
        RECT 758.150 18.120 760.295 18.260 ;
        RECT 758.150 18.060 758.470 18.120 ;
        RECT 760.005 18.075 760.295 18.120 ;
        RECT 760.005 14.180 760.295 14.225 ;
        RECT 2583.890 14.180 2584.210 14.240 ;
        RECT 760.005 14.040 2584.210 14.180 ;
        RECT 760.005 13.995 760.295 14.040 ;
        RECT 2583.890 13.980 2584.210 14.040 ;
      LAYER via ;
        RECT 681.820 2201.200 682.080 2201.460 ;
        RECT 685.500 2201.200 685.760 2201.460 ;
        RECT 758.180 18.060 758.440 18.320 ;
        RECT 2583.920 13.980 2584.180 14.240 ;
      LAYER met2 ;
        RECT 685.490 2207.435 685.770 2207.805 ;
        RECT 685.560 2201.490 685.700 2207.435 ;
        RECT 681.820 2201.170 682.080 2201.490 ;
        RECT 685.500 2201.170 685.760 2201.490 ;
        RECT 681.880 20.245 682.020 2201.170 ;
        RECT 681.810 19.875 682.090 20.245 ;
        RECT 758.170 19.875 758.450 20.245 ;
        RECT 758.240 18.350 758.380 19.875 ;
        RECT 758.180 18.030 758.440 18.350 ;
        RECT 2583.920 13.950 2584.180 14.270 ;
        RECT 2583.980 2.400 2584.120 13.950 ;
        RECT 2583.770 -4.800 2584.330 2.400 ;
      LAYER via2 ;
        RECT 685.490 2207.480 685.770 2207.760 ;
        RECT 681.810 19.920 682.090 20.200 ;
        RECT 758.170 19.920 758.450 20.200 ;
      LAYER met3 ;
        RECT 685.465 2207.770 685.795 2207.785 ;
        RECT 715.810 2207.770 719.810 2207.775 ;
        RECT 685.465 2207.470 719.810 2207.770 ;
        RECT 685.465 2207.455 685.795 2207.470 ;
        RECT 715.810 2207.175 719.810 2207.470 ;
        RECT 681.785 20.210 682.115 20.225 ;
        RECT 758.145 20.210 758.475 20.225 ;
        RECT 681.785 19.910 758.475 20.210 ;
        RECT 681.785 19.895 682.115 19.910 ;
        RECT 758.145 19.895 758.475 19.910 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 820.710 553.560 821.030 553.820 ;
        RECT 820.800 553.140 820.940 553.560 ;
        RECT 820.710 552.880 821.030 553.140 ;
        RECT 817.490 20.640 817.810 20.700 ;
        RECT 820.710 20.640 821.030 20.700 ;
        RECT 817.490 20.500 821.030 20.640 ;
        RECT 817.490 20.440 817.810 20.500 ;
        RECT 820.710 20.440 821.030 20.500 ;
      LAYER via ;
        RECT 820.740 553.560 821.000 553.820 ;
        RECT 820.740 552.880 821.000 553.140 ;
        RECT 817.520 20.440 817.780 20.700 ;
        RECT 820.740 20.440 821.000 20.700 ;
      LAYER met2 ;
        RECT 1700.710 2393.075 1700.990 2393.445 ;
        RECT 1700.780 2390.045 1700.920 2393.075 ;
        RECT 1664.370 2389.675 1664.650 2390.045 ;
        RECT 1700.710 2389.675 1700.990 2390.045 ;
        RECT 1664.440 2377.880 1664.580 2389.675 ;
        RECT 1664.420 2373.880 1664.700 2377.880 ;
        RECT 820.730 1320.715 821.010 1321.085 ;
        RECT 820.800 553.850 820.940 1320.715 ;
        RECT 820.740 553.530 821.000 553.850 ;
        RECT 820.740 552.850 821.000 553.170 ;
        RECT 820.800 20.730 820.940 552.850 ;
        RECT 817.520 20.410 817.780 20.730 ;
        RECT 820.740 20.410 821.000 20.730 ;
        RECT 817.580 2.400 817.720 20.410 ;
        RECT 817.370 -4.800 817.930 2.400 ;
      LAYER via2 ;
        RECT 1700.710 2393.120 1700.990 2393.400 ;
        RECT 1664.370 2389.720 1664.650 2390.000 ;
        RECT 1700.710 2389.720 1700.990 2390.000 ;
        RECT 820.730 1320.760 821.010 1321.040 ;
      LAYER met3 ;
        RECT 1700.685 2393.410 1701.015 2393.425 ;
        RECT 1773.110 2393.410 1773.490 2393.420 ;
        RECT 1700.685 2393.110 1773.490 2393.410 ;
        RECT 1700.685 2393.095 1701.015 2393.110 ;
        RECT 1773.110 2393.100 1773.490 2393.110 ;
        RECT 1664.345 2390.010 1664.675 2390.025 ;
        RECT 1700.685 2390.010 1701.015 2390.025 ;
        RECT 1664.345 2389.710 1701.015 2390.010 ;
        RECT 1664.345 2389.695 1664.675 2389.710 ;
        RECT 1700.685 2389.695 1701.015 2389.710 ;
        RECT 820.705 1321.050 821.035 1321.065 ;
        RECT 1773.110 1321.050 1773.490 1321.060 ;
        RECT 820.705 1320.750 1773.490 1321.050 ;
        RECT 820.705 1320.735 821.035 1320.750 ;
        RECT 1773.110 1320.740 1773.490 1320.750 ;
      LAYER via3 ;
        RECT 1773.140 2393.100 1773.460 2393.420 ;
        RECT 1773.140 1320.740 1773.460 1321.060 ;
      LAYER met4 ;
        RECT 1773.135 2393.095 1773.465 2393.425 ;
        RECT 1773.150 1321.065 1773.450 2393.095 ;
        RECT 1773.135 1320.735 1773.465 1321.065 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1248.050 60.420 1248.370 60.480 ;
        RECT 2601.370 60.420 2601.690 60.480 ;
        RECT 1248.050 60.280 2601.690 60.420 ;
        RECT 1248.050 60.220 1248.370 60.280 ;
        RECT 2601.370 60.220 2601.690 60.280 ;
      LAYER via ;
        RECT 1248.080 60.220 1248.340 60.480 ;
        RECT 2601.400 60.220 2601.660 60.480 ;
      LAYER met2 ;
        RECT 1244.900 1323.690 1245.180 1327.135 ;
        RECT 1244.900 1323.550 1248.280 1323.690 ;
        RECT 1244.900 1323.135 1245.180 1323.550 ;
        RECT 1248.140 60.510 1248.280 1323.550 ;
        RECT 1248.080 60.190 1248.340 60.510 ;
        RECT 2601.400 60.190 2601.660 60.510 ;
        RECT 2601.460 2.400 2601.600 60.190 ;
        RECT 2601.250 -4.800 2601.810 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2615.245 2173.705 2615.415 2221.815 ;
        RECT 2615.245 2077.145 2615.415 2125.255 ;
        RECT 2615.245 1980.245 2615.415 2028.355 ;
        RECT 2615.245 1883.685 2615.415 1931.795 ;
        RECT 2615.245 1787.125 2615.415 1835.235 ;
        RECT 2615.245 1690.565 2615.415 1738.335 ;
        RECT 2615.245 1594.005 2615.415 1642.115 ;
        RECT 2615.245 1497.445 2615.415 1545.555 ;
        RECT 2615.245 1400.885 2615.415 1448.995 ;
        RECT 2615.245 1304.325 2615.415 1352.435 ;
        RECT 2615.245 1207.425 2615.415 1255.875 ;
        RECT 2615.245 628.065 2615.415 675.835 ;
        RECT 2615.245 531.505 2615.415 579.615 ;
        RECT 2615.245 434.945 2615.415 483.055 ;
        RECT 2615.245 338.045 2615.415 386.155 ;
        RECT 2615.245 241.485 2615.415 289.595 ;
        RECT 2615.245 144.925 2615.415 193.035 ;
        RECT 2615.245 48.365 2615.415 96.475 ;
      LAYER mcon ;
        RECT 2615.245 2221.645 2615.415 2221.815 ;
        RECT 2615.245 2125.085 2615.415 2125.255 ;
        RECT 2615.245 2028.185 2615.415 2028.355 ;
        RECT 2615.245 1931.625 2615.415 1931.795 ;
        RECT 2615.245 1835.065 2615.415 1835.235 ;
        RECT 2615.245 1738.165 2615.415 1738.335 ;
        RECT 2615.245 1641.945 2615.415 1642.115 ;
        RECT 2615.245 1545.385 2615.415 1545.555 ;
        RECT 2615.245 1448.825 2615.415 1448.995 ;
        RECT 2615.245 1352.265 2615.415 1352.435 ;
        RECT 2615.245 1255.705 2615.415 1255.875 ;
        RECT 2615.245 675.665 2615.415 675.835 ;
        RECT 2615.245 579.445 2615.415 579.615 ;
        RECT 2615.245 482.885 2615.415 483.055 ;
        RECT 2615.245 385.985 2615.415 386.155 ;
        RECT 2615.245 289.425 2615.415 289.595 ;
        RECT 2615.245 192.865 2615.415 193.035 ;
        RECT 2615.245 96.305 2615.415 96.475 ;
      LAYER met1 ;
        RECT 763.210 2377.860 763.530 2377.920 ;
        RECT 896.610 2377.860 896.930 2377.920 ;
        RECT 763.210 2377.720 896.930 2377.860 ;
        RECT 763.210 2377.660 763.530 2377.720 ;
        RECT 896.610 2377.660 896.930 2377.720 ;
        RECT 2614.250 2318.360 2614.570 2318.420 ;
        RECT 2615.170 2318.360 2615.490 2318.420 ;
        RECT 2614.250 2318.220 2615.490 2318.360 ;
        RECT 2614.250 2318.160 2614.570 2318.220 ;
        RECT 2615.170 2318.160 2615.490 2318.220 ;
        RECT 2615.170 2221.800 2615.490 2221.860 ;
        RECT 2614.975 2221.660 2615.490 2221.800 ;
        RECT 2615.170 2221.600 2615.490 2221.660 ;
        RECT 2615.170 2173.860 2615.490 2173.920 ;
        RECT 2614.975 2173.720 2615.490 2173.860 ;
        RECT 2615.170 2173.660 2615.490 2173.720 ;
        RECT 2615.170 2125.240 2615.490 2125.300 ;
        RECT 2614.975 2125.100 2615.490 2125.240 ;
        RECT 2615.170 2125.040 2615.490 2125.100 ;
        RECT 2615.170 2077.300 2615.490 2077.360 ;
        RECT 2614.975 2077.160 2615.490 2077.300 ;
        RECT 2615.170 2077.100 2615.490 2077.160 ;
        RECT 2615.170 2028.340 2615.490 2028.400 ;
        RECT 2614.975 2028.200 2615.490 2028.340 ;
        RECT 2615.170 2028.140 2615.490 2028.200 ;
        RECT 2615.170 1980.400 2615.490 1980.460 ;
        RECT 2614.975 1980.260 2615.490 1980.400 ;
        RECT 2615.170 1980.200 2615.490 1980.260 ;
        RECT 2615.170 1931.780 2615.490 1931.840 ;
        RECT 2614.975 1931.640 2615.490 1931.780 ;
        RECT 2615.170 1931.580 2615.490 1931.640 ;
        RECT 2615.170 1883.840 2615.490 1883.900 ;
        RECT 2614.975 1883.700 2615.490 1883.840 ;
        RECT 2615.170 1883.640 2615.490 1883.700 ;
        RECT 2615.170 1835.220 2615.490 1835.280 ;
        RECT 2614.975 1835.080 2615.490 1835.220 ;
        RECT 2615.170 1835.020 2615.490 1835.080 ;
        RECT 2615.170 1787.280 2615.490 1787.340 ;
        RECT 2614.975 1787.140 2615.490 1787.280 ;
        RECT 2615.170 1787.080 2615.490 1787.140 ;
        RECT 2615.170 1739.820 2615.490 1740.080 ;
        RECT 2615.260 1739.060 2615.400 1739.820 ;
        RECT 2615.170 1738.800 2615.490 1739.060 ;
        RECT 2615.170 1738.320 2615.490 1738.380 ;
        RECT 2614.975 1738.180 2615.490 1738.320 ;
        RECT 2615.170 1738.120 2615.490 1738.180 ;
        RECT 2615.170 1690.720 2615.490 1690.780 ;
        RECT 2614.975 1690.580 2615.490 1690.720 ;
        RECT 2615.170 1690.520 2615.490 1690.580 ;
        RECT 2615.170 1642.100 2615.490 1642.160 ;
        RECT 2614.975 1641.960 2615.490 1642.100 ;
        RECT 2615.170 1641.900 2615.490 1641.960 ;
        RECT 2615.170 1594.160 2615.490 1594.220 ;
        RECT 2614.975 1594.020 2615.490 1594.160 ;
        RECT 2615.170 1593.960 2615.490 1594.020 ;
        RECT 2615.170 1545.540 2615.490 1545.600 ;
        RECT 2614.975 1545.400 2615.490 1545.540 ;
        RECT 2615.170 1545.340 2615.490 1545.400 ;
        RECT 2615.170 1497.600 2615.490 1497.660 ;
        RECT 2614.975 1497.460 2615.490 1497.600 ;
        RECT 2615.170 1497.400 2615.490 1497.460 ;
        RECT 2615.170 1448.980 2615.490 1449.040 ;
        RECT 2614.975 1448.840 2615.490 1448.980 ;
        RECT 2615.170 1448.780 2615.490 1448.840 ;
        RECT 2615.170 1401.040 2615.490 1401.100 ;
        RECT 2614.975 1400.900 2615.490 1401.040 ;
        RECT 2615.170 1400.840 2615.490 1400.900 ;
        RECT 2615.170 1352.420 2615.490 1352.480 ;
        RECT 2614.975 1352.280 2615.490 1352.420 ;
        RECT 2615.170 1352.220 2615.490 1352.280 ;
        RECT 2615.170 1304.480 2615.490 1304.540 ;
        RECT 2614.975 1304.340 2615.490 1304.480 ;
        RECT 2615.170 1304.280 2615.490 1304.340 ;
        RECT 2615.170 1255.860 2615.490 1255.920 ;
        RECT 2614.975 1255.720 2615.490 1255.860 ;
        RECT 2615.170 1255.660 2615.490 1255.720 ;
        RECT 2615.170 1207.580 2615.490 1207.640 ;
        RECT 2614.975 1207.440 2615.490 1207.580 ;
        RECT 2615.170 1207.380 2615.490 1207.440 ;
        RECT 2614.250 1111.020 2614.570 1111.080 ;
        RECT 2615.170 1111.020 2615.490 1111.080 ;
        RECT 2614.250 1110.880 2615.490 1111.020 ;
        RECT 2614.250 1110.820 2614.570 1110.880 ;
        RECT 2615.170 1110.820 2615.490 1110.880 ;
        RECT 2614.250 1014.460 2614.570 1014.520 ;
        RECT 2615.170 1014.460 2615.490 1014.520 ;
        RECT 2614.250 1014.320 2615.490 1014.460 ;
        RECT 2614.250 1014.260 2614.570 1014.320 ;
        RECT 2615.170 1014.260 2615.490 1014.320 ;
        RECT 2614.250 917.900 2614.570 917.960 ;
        RECT 2615.170 917.900 2615.490 917.960 ;
        RECT 2614.250 917.760 2615.490 917.900 ;
        RECT 2614.250 917.700 2614.570 917.760 ;
        RECT 2615.170 917.700 2615.490 917.760 ;
        RECT 2614.250 772.720 2614.570 772.780 ;
        RECT 2615.170 772.720 2615.490 772.780 ;
        RECT 2614.250 772.580 2615.490 772.720 ;
        RECT 2614.250 772.520 2614.570 772.580 ;
        RECT 2615.170 772.520 2615.490 772.580 ;
        RECT 2615.170 675.820 2615.490 675.880 ;
        RECT 2614.975 675.680 2615.490 675.820 ;
        RECT 2615.170 675.620 2615.490 675.680 ;
        RECT 2615.170 628.220 2615.490 628.280 ;
        RECT 2614.975 628.080 2615.490 628.220 ;
        RECT 2615.170 628.020 2615.490 628.080 ;
        RECT 2615.170 579.600 2615.490 579.660 ;
        RECT 2614.975 579.460 2615.490 579.600 ;
        RECT 2615.170 579.400 2615.490 579.460 ;
        RECT 2615.170 531.660 2615.490 531.720 ;
        RECT 2614.975 531.520 2615.490 531.660 ;
        RECT 2615.170 531.460 2615.490 531.520 ;
        RECT 2615.170 483.040 2615.490 483.100 ;
        RECT 2614.975 482.900 2615.490 483.040 ;
        RECT 2615.170 482.840 2615.490 482.900 ;
        RECT 2615.170 435.100 2615.490 435.160 ;
        RECT 2614.975 434.960 2615.490 435.100 ;
        RECT 2615.170 434.900 2615.490 434.960 ;
        RECT 2615.170 386.140 2615.490 386.200 ;
        RECT 2614.975 386.000 2615.490 386.140 ;
        RECT 2615.170 385.940 2615.490 386.000 ;
        RECT 2615.170 338.200 2615.490 338.260 ;
        RECT 2614.975 338.060 2615.490 338.200 ;
        RECT 2615.170 338.000 2615.490 338.060 ;
        RECT 2615.170 289.580 2615.490 289.640 ;
        RECT 2614.975 289.440 2615.490 289.580 ;
        RECT 2615.170 289.380 2615.490 289.440 ;
        RECT 2615.170 241.640 2615.490 241.700 ;
        RECT 2614.975 241.500 2615.490 241.640 ;
        RECT 2615.170 241.440 2615.490 241.500 ;
        RECT 2615.170 193.020 2615.490 193.080 ;
        RECT 2614.975 192.880 2615.490 193.020 ;
        RECT 2615.170 192.820 2615.490 192.880 ;
        RECT 2615.170 145.080 2615.490 145.140 ;
        RECT 2614.975 144.940 2615.490 145.080 ;
        RECT 2615.170 144.880 2615.490 144.940 ;
        RECT 2615.170 96.460 2615.490 96.520 ;
        RECT 2614.975 96.320 2615.490 96.460 ;
        RECT 2615.170 96.260 2615.490 96.320 ;
        RECT 2615.170 48.520 2615.490 48.580 ;
        RECT 2614.975 48.380 2615.490 48.520 ;
        RECT 2615.170 48.320 2615.490 48.380 ;
        RECT 2615.170 14.180 2615.490 14.240 ;
        RECT 2615.170 14.040 2619.540 14.180 ;
        RECT 2615.170 13.980 2615.490 14.040 ;
        RECT 2619.400 13.900 2619.540 14.040 ;
        RECT 2619.310 13.640 2619.630 13.900 ;
      LAYER via ;
        RECT 763.240 2377.660 763.500 2377.920 ;
        RECT 896.640 2377.660 896.900 2377.920 ;
        RECT 2614.280 2318.160 2614.540 2318.420 ;
        RECT 2615.200 2318.160 2615.460 2318.420 ;
        RECT 2615.200 2221.600 2615.460 2221.860 ;
        RECT 2615.200 2173.660 2615.460 2173.920 ;
        RECT 2615.200 2125.040 2615.460 2125.300 ;
        RECT 2615.200 2077.100 2615.460 2077.360 ;
        RECT 2615.200 2028.140 2615.460 2028.400 ;
        RECT 2615.200 1980.200 2615.460 1980.460 ;
        RECT 2615.200 1931.580 2615.460 1931.840 ;
        RECT 2615.200 1883.640 2615.460 1883.900 ;
        RECT 2615.200 1835.020 2615.460 1835.280 ;
        RECT 2615.200 1787.080 2615.460 1787.340 ;
        RECT 2615.200 1739.820 2615.460 1740.080 ;
        RECT 2615.200 1738.800 2615.460 1739.060 ;
        RECT 2615.200 1738.120 2615.460 1738.380 ;
        RECT 2615.200 1690.520 2615.460 1690.780 ;
        RECT 2615.200 1641.900 2615.460 1642.160 ;
        RECT 2615.200 1593.960 2615.460 1594.220 ;
        RECT 2615.200 1545.340 2615.460 1545.600 ;
        RECT 2615.200 1497.400 2615.460 1497.660 ;
        RECT 2615.200 1448.780 2615.460 1449.040 ;
        RECT 2615.200 1400.840 2615.460 1401.100 ;
        RECT 2615.200 1352.220 2615.460 1352.480 ;
        RECT 2615.200 1304.280 2615.460 1304.540 ;
        RECT 2615.200 1255.660 2615.460 1255.920 ;
        RECT 2615.200 1207.380 2615.460 1207.640 ;
        RECT 2614.280 1110.820 2614.540 1111.080 ;
        RECT 2615.200 1110.820 2615.460 1111.080 ;
        RECT 2614.280 1014.260 2614.540 1014.520 ;
        RECT 2615.200 1014.260 2615.460 1014.520 ;
        RECT 2614.280 917.700 2614.540 917.960 ;
        RECT 2615.200 917.700 2615.460 917.960 ;
        RECT 2614.280 772.520 2614.540 772.780 ;
        RECT 2615.200 772.520 2615.460 772.780 ;
        RECT 2615.200 675.620 2615.460 675.880 ;
        RECT 2615.200 628.020 2615.460 628.280 ;
        RECT 2615.200 579.400 2615.460 579.660 ;
        RECT 2615.200 531.460 2615.460 531.720 ;
        RECT 2615.200 482.840 2615.460 483.100 ;
        RECT 2615.200 434.900 2615.460 435.160 ;
        RECT 2615.200 385.940 2615.460 386.200 ;
        RECT 2615.200 338.000 2615.460 338.260 ;
        RECT 2615.200 289.380 2615.460 289.640 ;
        RECT 2615.200 241.440 2615.460 241.700 ;
        RECT 2615.200 192.820 2615.460 193.080 ;
        RECT 2615.200 144.880 2615.460 145.140 ;
        RECT 2615.200 96.260 2615.460 96.520 ;
        RECT 2615.200 48.320 2615.460 48.580 ;
        RECT 2615.200 13.980 2615.460 14.240 ;
        RECT 2619.340 13.640 2619.600 13.900 ;
      LAYER met2 ;
        RECT 761.900 2377.690 762.180 2377.880 ;
        RECT 763.240 2377.690 763.500 2377.950 ;
        RECT 761.900 2377.630 763.500 2377.690 ;
        RECT 896.640 2377.630 896.900 2377.950 ;
        RECT 761.900 2377.550 763.440 2377.630 ;
        RECT 761.900 2373.880 762.180 2377.550 ;
        RECT 896.700 2376.445 896.840 2377.630 ;
        RECT 2609.210 2376.755 2609.490 2377.125 ;
        RECT 896.630 2376.075 896.910 2376.445 ;
        RECT 2609.280 2366.925 2609.420 2376.755 ;
        RECT 2609.210 2366.555 2609.490 2366.925 ;
        RECT 2615.190 2366.555 2615.470 2366.925 ;
        RECT 2615.260 2318.450 2615.400 2366.555 ;
        RECT 2614.280 2318.130 2614.540 2318.450 ;
        RECT 2615.200 2318.130 2615.460 2318.450 ;
        RECT 2614.340 2270.365 2614.480 2318.130 ;
        RECT 2614.270 2269.995 2614.550 2270.365 ;
        RECT 2615.190 2269.995 2615.470 2270.365 ;
        RECT 2615.260 2221.890 2615.400 2269.995 ;
        RECT 2615.200 2221.570 2615.460 2221.890 ;
        RECT 2615.200 2173.630 2615.460 2173.950 ;
        RECT 2615.260 2125.330 2615.400 2173.630 ;
        RECT 2615.200 2125.010 2615.460 2125.330 ;
        RECT 2615.200 2077.070 2615.460 2077.390 ;
        RECT 2615.260 2028.430 2615.400 2077.070 ;
        RECT 2615.200 2028.110 2615.460 2028.430 ;
        RECT 2615.200 1980.170 2615.460 1980.490 ;
        RECT 2615.260 1931.870 2615.400 1980.170 ;
        RECT 2615.200 1931.550 2615.460 1931.870 ;
        RECT 2615.200 1883.610 2615.460 1883.930 ;
        RECT 2615.260 1835.310 2615.400 1883.610 ;
        RECT 2615.200 1834.990 2615.460 1835.310 ;
        RECT 2615.200 1787.050 2615.460 1787.370 ;
        RECT 2615.260 1740.110 2615.400 1787.050 ;
        RECT 2615.200 1739.790 2615.460 1740.110 ;
        RECT 2615.200 1738.770 2615.460 1739.090 ;
        RECT 2615.260 1738.410 2615.400 1738.770 ;
        RECT 2615.200 1738.090 2615.460 1738.410 ;
        RECT 2615.200 1690.490 2615.460 1690.810 ;
        RECT 2615.260 1642.190 2615.400 1690.490 ;
        RECT 2615.200 1641.870 2615.460 1642.190 ;
        RECT 2615.200 1593.930 2615.460 1594.250 ;
        RECT 2615.260 1545.630 2615.400 1593.930 ;
        RECT 2615.200 1545.310 2615.460 1545.630 ;
        RECT 2615.200 1497.370 2615.460 1497.690 ;
        RECT 2615.260 1449.070 2615.400 1497.370 ;
        RECT 2615.200 1448.750 2615.460 1449.070 ;
        RECT 2615.200 1400.810 2615.460 1401.130 ;
        RECT 2615.260 1352.510 2615.400 1400.810 ;
        RECT 2615.200 1352.190 2615.460 1352.510 ;
        RECT 2615.200 1304.250 2615.460 1304.570 ;
        RECT 2615.260 1255.950 2615.400 1304.250 ;
        RECT 2615.200 1255.630 2615.460 1255.950 ;
        RECT 2615.200 1207.350 2615.460 1207.670 ;
        RECT 2615.260 1159.245 2615.400 1207.350 ;
        RECT 2614.270 1158.875 2614.550 1159.245 ;
        RECT 2615.190 1158.875 2615.470 1159.245 ;
        RECT 2614.340 1111.110 2614.480 1158.875 ;
        RECT 2614.280 1110.790 2614.540 1111.110 ;
        RECT 2615.200 1110.790 2615.460 1111.110 ;
        RECT 2615.260 1062.685 2615.400 1110.790 ;
        RECT 2614.270 1062.315 2614.550 1062.685 ;
        RECT 2615.190 1062.315 2615.470 1062.685 ;
        RECT 2614.340 1014.550 2614.480 1062.315 ;
        RECT 2614.280 1014.230 2614.540 1014.550 ;
        RECT 2615.200 1014.230 2615.460 1014.550 ;
        RECT 2615.260 966.125 2615.400 1014.230 ;
        RECT 2614.270 965.755 2614.550 966.125 ;
        RECT 2615.190 965.755 2615.470 966.125 ;
        RECT 2614.340 917.990 2614.480 965.755 ;
        RECT 2614.280 917.670 2614.540 917.990 ;
        RECT 2615.200 917.670 2615.460 917.990 ;
        RECT 2615.260 869.565 2615.400 917.670 ;
        RECT 2614.270 869.195 2614.550 869.565 ;
        RECT 2615.190 869.195 2615.470 869.565 ;
        RECT 2614.340 821.285 2614.480 869.195 ;
        RECT 2614.270 820.915 2614.550 821.285 ;
        RECT 2615.190 820.915 2615.470 821.285 ;
        RECT 2615.260 772.810 2615.400 820.915 ;
        RECT 2614.280 772.490 2614.540 772.810 ;
        RECT 2615.200 772.490 2615.460 772.810 ;
        RECT 2614.340 724.725 2614.480 772.490 ;
        RECT 2614.270 724.355 2614.550 724.725 ;
        RECT 2615.190 724.355 2615.470 724.725 ;
        RECT 2615.260 675.910 2615.400 724.355 ;
        RECT 2615.200 675.590 2615.460 675.910 ;
        RECT 2615.200 627.990 2615.460 628.310 ;
        RECT 2615.260 579.690 2615.400 627.990 ;
        RECT 2615.200 579.370 2615.460 579.690 ;
        RECT 2615.200 531.430 2615.460 531.750 ;
        RECT 2615.260 483.130 2615.400 531.430 ;
        RECT 2615.200 482.810 2615.460 483.130 ;
        RECT 2615.200 434.870 2615.460 435.190 ;
        RECT 2615.260 386.230 2615.400 434.870 ;
        RECT 2615.200 385.910 2615.460 386.230 ;
        RECT 2615.200 337.970 2615.460 338.290 ;
        RECT 2615.260 289.670 2615.400 337.970 ;
        RECT 2615.200 289.350 2615.460 289.670 ;
        RECT 2615.200 241.410 2615.460 241.730 ;
        RECT 2615.260 193.110 2615.400 241.410 ;
        RECT 2615.200 192.790 2615.460 193.110 ;
        RECT 2615.200 144.850 2615.460 145.170 ;
        RECT 2615.260 96.550 2615.400 144.850 ;
        RECT 2615.200 96.230 2615.460 96.550 ;
        RECT 2615.200 48.290 2615.460 48.610 ;
        RECT 2615.260 14.270 2615.400 48.290 ;
        RECT 2615.200 13.950 2615.460 14.270 ;
        RECT 2619.340 13.610 2619.600 13.930 ;
        RECT 2619.400 2.400 2619.540 13.610 ;
        RECT 2619.190 -4.800 2619.750 2.400 ;
      LAYER via2 ;
        RECT 2609.210 2376.800 2609.490 2377.080 ;
        RECT 896.630 2376.120 896.910 2376.400 ;
        RECT 2609.210 2366.600 2609.490 2366.880 ;
        RECT 2615.190 2366.600 2615.470 2366.880 ;
        RECT 2614.270 2270.040 2614.550 2270.320 ;
        RECT 2615.190 2270.040 2615.470 2270.320 ;
        RECT 2614.270 1158.920 2614.550 1159.200 ;
        RECT 2615.190 1158.920 2615.470 1159.200 ;
        RECT 2614.270 1062.360 2614.550 1062.640 ;
        RECT 2615.190 1062.360 2615.470 1062.640 ;
        RECT 2614.270 965.800 2614.550 966.080 ;
        RECT 2615.190 965.800 2615.470 966.080 ;
        RECT 2614.270 869.240 2614.550 869.520 ;
        RECT 2615.190 869.240 2615.470 869.520 ;
        RECT 2614.270 820.960 2614.550 821.240 ;
        RECT 2615.190 820.960 2615.470 821.240 ;
        RECT 2614.270 724.400 2614.550 724.680 ;
        RECT 2615.190 724.400 2615.470 724.680 ;
      LAYER met3 ;
        RECT 2609.185 2377.090 2609.515 2377.105 ;
        RECT 930.430 2376.790 2609.515 2377.090 ;
        RECT 896.605 2376.410 896.935 2376.425 ;
        RECT 930.430 2376.410 930.730 2376.790 ;
        RECT 2609.185 2376.775 2609.515 2376.790 ;
        RECT 896.605 2376.110 930.730 2376.410 ;
        RECT 896.605 2376.095 896.935 2376.110 ;
        RECT 2609.185 2366.890 2609.515 2366.905 ;
        RECT 2615.165 2366.890 2615.495 2366.905 ;
        RECT 2609.185 2366.590 2615.495 2366.890 ;
        RECT 2609.185 2366.575 2609.515 2366.590 ;
        RECT 2615.165 2366.575 2615.495 2366.590 ;
        RECT 2614.245 2270.330 2614.575 2270.345 ;
        RECT 2615.165 2270.330 2615.495 2270.345 ;
        RECT 2614.245 2270.030 2615.495 2270.330 ;
        RECT 2614.245 2270.015 2614.575 2270.030 ;
        RECT 2615.165 2270.015 2615.495 2270.030 ;
        RECT 2614.245 1159.210 2614.575 1159.225 ;
        RECT 2615.165 1159.210 2615.495 1159.225 ;
        RECT 2614.245 1158.910 2615.495 1159.210 ;
        RECT 2614.245 1158.895 2614.575 1158.910 ;
        RECT 2615.165 1158.895 2615.495 1158.910 ;
        RECT 2614.245 1062.650 2614.575 1062.665 ;
        RECT 2615.165 1062.650 2615.495 1062.665 ;
        RECT 2614.245 1062.350 2615.495 1062.650 ;
        RECT 2614.245 1062.335 2614.575 1062.350 ;
        RECT 2615.165 1062.335 2615.495 1062.350 ;
        RECT 2614.245 966.090 2614.575 966.105 ;
        RECT 2615.165 966.090 2615.495 966.105 ;
        RECT 2614.245 965.790 2615.495 966.090 ;
        RECT 2614.245 965.775 2614.575 965.790 ;
        RECT 2615.165 965.775 2615.495 965.790 ;
        RECT 2614.245 869.530 2614.575 869.545 ;
        RECT 2615.165 869.530 2615.495 869.545 ;
        RECT 2614.245 869.230 2615.495 869.530 ;
        RECT 2614.245 869.215 2614.575 869.230 ;
        RECT 2615.165 869.215 2615.495 869.230 ;
        RECT 2614.245 821.250 2614.575 821.265 ;
        RECT 2615.165 821.250 2615.495 821.265 ;
        RECT 2614.245 820.950 2615.495 821.250 ;
        RECT 2614.245 820.935 2614.575 820.950 ;
        RECT 2615.165 820.935 2615.495 820.950 ;
        RECT 2614.245 724.690 2614.575 724.705 ;
        RECT 2615.165 724.690 2615.495 724.705 ;
        RECT 2614.245 724.390 2615.495 724.690 ;
        RECT 2614.245 724.375 2614.575 724.390 ;
        RECT 2615.165 724.375 2615.495 724.390 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1331.310 66.200 1331.630 66.260 ;
        RECT 2636.790 66.200 2637.110 66.260 ;
        RECT 1331.310 66.060 2637.110 66.200 ;
        RECT 1331.310 66.000 1331.630 66.060 ;
        RECT 2636.790 66.000 2637.110 66.060 ;
      LAYER via ;
        RECT 1331.340 66.000 1331.600 66.260 ;
        RECT 2636.820 66.000 2637.080 66.260 ;
      LAYER met2 ;
        RECT 1331.380 1323.135 1331.660 1327.135 ;
        RECT 1331.400 66.290 1331.540 1323.135 ;
        RECT 1331.340 65.970 1331.600 66.290 ;
        RECT 2636.820 65.970 2637.080 66.290 ;
        RECT 2636.880 24.210 2637.020 65.970 ;
        RECT 2636.880 24.070 2637.480 24.210 ;
        RECT 2637.340 2.400 2637.480 24.070 ;
        RECT 2637.130 -4.800 2637.690 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 717.745 1894.565 717.915 1936.895 ;
        RECT 717.285 1658.605 717.455 1694.135 ;
        RECT 718.205 1307.385 718.375 1430.295 ;
      LAYER mcon ;
        RECT 717.745 1936.725 717.915 1936.895 ;
        RECT 717.285 1693.965 717.455 1694.135 ;
        RECT 718.205 1430.125 718.375 1430.295 ;
      LAYER met1 ;
        RECT 717.670 1936.880 717.990 1936.940 ;
        RECT 717.475 1936.740 717.990 1936.880 ;
        RECT 717.670 1936.680 717.990 1936.740 ;
        RECT 717.670 1894.720 717.990 1894.780 ;
        RECT 717.475 1894.580 717.990 1894.720 ;
        RECT 717.670 1894.520 717.990 1894.580 ;
        RECT 717.210 1694.120 717.530 1694.180 ;
        RECT 717.015 1693.980 717.530 1694.120 ;
        RECT 717.210 1693.920 717.530 1693.980 ;
        RECT 717.225 1658.760 717.515 1658.805 ;
        RECT 717.225 1658.620 717.900 1658.760 ;
        RECT 717.225 1658.575 717.515 1658.620 ;
        RECT 717.760 1658.420 717.900 1658.620 ;
        RECT 717.760 1658.280 718.820 1658.420 ;
        RECT 718.680 1658.140 718.820 1658.280 ;
        RECT 718.590 1657.880 718.910 1658.140 ;
        RECT 717.210 1430.280 717.530 1430.340 ;
        RECT 718.145 1430.280 718.435 1430.325 ;
        RECT 717.210 1430.140 718.435 1430.280 ;
        RECT 717.210 1430.080 717.530 1430.140 ;
        RECT 718.145 1430.095 718.435 1430.140 ;
        RECT 718.130 1307.540 718.450 1307.600 ;
        RECT 717.935 1307.400 718.450 1307.540 ;
        RECT 718.130 1307.340 718.450 1307.400 ;
        RECT 2649.670 62.120 2649.990 62.180 ;
        RECT 2655.190 62.120 2655.510 62.180 ;
        RECT 2649.670 61.980 2655.510 62.120 ;
        RECT 2649.670 61.920 2649.990 61.980 ;
        RECT 2655.190 61.920 2655.510 61.980 ;
      LAYER via ;
        RECT 717.700 1936.680 717.960 1936.940 ;
        RECT 717.700 1894.520 717.960 1894.780 ;
        RECT 717.240 1693.920 717.500 1694.180 ;
        RECT 718.620 1657.880 718.880 1658.140 ;
        RECT 717.240 1430.080 717.500 1430.340 ;
        RECT 718.160 1307.340 718.420 1307.600 ;
        RECT 2649.700 61.920 2649.960 62.180 ;
        RECT 2655.220 61.920 2655.480 62.180 ;
      LAYER met2 ;
        RECT 717.690 1983.035 717.970 1983.405 ;
        RECT 717.760 1936.970 717.900 1983.035 ;
        RECT 717.700 1936.650 717.960 1936.970 ;
        RECT 717.700 1894.490 717.960 1894.810 ;
        RECT 717.760 1888.885 717.900 1894.490 ;
        RECT 717.690 1888.515 717.970 1888.885 ;
        RECT 717.230 1695.395 717.510 1695.765 ;
        RECT 717.300 1694.210 717.440 1695.395 ;
        RECT 717.240 1693.890 717.500 1694.210 ;
        RECT 718.620 1657.850 718.880 1658.170 ;
        RECT 718.680 1597.845 718.820 1657.850 ;
        RECT 718.610 1597.475 718.890 1597.845 ;
        RECT 718.610 1563.475 718.890 1563.845 ;
        RECT 718.680 1545.485 718.820 1563.475 ;
        RECT 718.610 1545.115 718.890 1545.485 ;
        RECT 717.230 1430.195 717.510 1430.565 ;
        RECT 717.240 1430.050 717.500 1430.195 ;
        RECT 718.160 1307.310 718.420 1307.630 ;
        RECT 718.220 1300.685 718.360 1307.310 ;
        RECT 718.150 1300.315 718.430 1300.685 ;
        RECT 2649.690 1300.315 2649.970 1300.685 ;
        RECT 2649.760 62.210 2649.900 1300.315 ;
        RECT 2649.700 61.890 2649.960 62.210 ;
        RECT 2655.220 61.890 2655.480 62.210 ;
        RECT 2655.280 2.400 2655.420 61.890 ;
        RECT 2655.070 -4.800 2655.630 2.400 ;
      LAYER via2 ;
        RECT 717.690 1983.080 717.970 1983.360 ;
        RECT 717.690 1888.560 717.970 1888.840 ;
        RECT 717.230 1695.440 717.510 1695.720 ;
        RECT 718.610 1597.520 718.890 1597.800 ;
        RECT 718.610 1563.520 718.890 1563.800 ;
        RECT 718.610 1545.160 718.890 1545.440 ;
        RECT 717.230 1430.240 717.510 1430.520 ;
        RECT 718.150 1300.360 718.430 1300.640 ;
        RECT 2649.690 1300.360 2649.970 1300.640 ;
      LAYER met3 ;
        RECT 715.810 1985.495 719.810 1986.095 ;
        RECT 717.910 1983.385 718.210 1985.495 ;
        RECT 717.665 1983.070 718.210 1983.385 ;
        RECT 717.665 1983.055 717.995 1983.070 ;
        RECT 717.665 1888.860 717.995 1888.865 ;
        RECT 717.665 1888.850 718.250 1888.860 ;
        RECT 717.440 1888.550 718.250 1888.850 ;
        RECT 717.665 1888.540 718.250 1888.550 ;
        RECT 717.665 1888.535 717.995 1888.540 ;
        RECT 717.205 1695.730 717.535 1695.745 ;
        RECT 717.870 1695.730 718.250 1695.740 ;
        RECT 717.205 1695.430 718.250 1695.730 ;
        RECT 717.205 1695.415 717.535 1695.430 ;
        RECT 717.870 1695.420 718.250 1695.430 ;
        RECT 717.870 1597.810 718.250 1597.820 ;
        RECT 718.585 1597.810 718.915 1597.825 ;
        RECT 717.870 1597.510 718.915 1597.810 ;
        RECT 717.870 1597.500 718.250 1597.510 ;
        RECT 718.585 1597.495 718.915 1597.510 ;
        RECT 717.870 1563.810 718.250 1563.820 ;
        RECT 718.585 1563.810 718.915 1563.825 ;
        RECT 717.870 1563.510 718.915 1563.810 ;
        RECT 717.870 1563.500 718.250 1563.510 ;
        RECT 718.585 1563.495 718.915 1563.510 ;
        RECT 717.870 1545.450 718.250 1545.460 ;
        RECT 718.585 1545.450 718.915 1545.465 ;
        RECT 717.870 1545.150 718.915 1545.450 ;
        RECT 717.870 1545.140 718.250 1545.150 ;
        RECT 718.585 1545.135 718.915 1545.150 ;
        RECT 717.205 1430.530 717.535 1430.545 ;
        RECT 717.870 1430.530 718.250 1430.540 ;
        RECT 717.205 1430.230 718.250 1430.530 ;
        RECT 717.205 1430.215 717.535 1430.230 ;
        RECT 717.870 1430.220 718.250 1430.230 ;
        RECT 718.125 1300.650 718.455 1300.665 ;
        RECT 2649.665 1300.650 2649.995 1300.665 ;
        RECT 718.125 1300.350 2649.995 1300.650 ;
        RECT 718.125 1300.335 718.455 1300.350 ;
        RECT 2649.665 1300.335 2649.995 1300.350 ;
      LAYER via3 ;
        RECT 717.900 1888.540 718.220 1888.860 ;
        RECT 717.900 1695.420 718.220 1695.740 ;
        RECT 717.900 1597.500 718.220 1597.820 ;
        RECT 717.900 1563.500 718.220 1563.820 ;
        RECT 717.900 1545.140 718.220 1545.460 ;
        RECT 717.900 1430.220 718.220 1430.540 ;
      LAYER met4 ;
        RECT 717.895 1888.535 718.225 1888.865 ;
        RECT 717.910 1695.745 718.210 1888.535 ;
        RECT 717.895 1695.415 718.225 1695.745 ;
        RECT 717.895 1597.495 718.225 1597.825 ;
        RECT 717.910 1563.825 718.210 1597.495 ;
        RECT 717.895 1563.495 718.225 1563.825 ;
        RECT 717.895 1545.135 718.225 1545.465 ;
        RECT 717.910 1430.545 718.210 1545.135 ;
        RECT 717.895 1430.215 718.225 1430.545 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2670.445 531.845 2670.615 579.615 ;
        RECT 2670.445 476.085 2670.615 524.195 ;
        RECT 2670.445 379.525 2670.615 427.635 ;
        RECT 2670.445 331.245 2670.615 339.235 ;
        RECT 2670.445 144.925 2670.615 210.375 ;
        RECT 2670.445 48.365 2670.615 137.955 ;
      LAYER mcon ;
        RECT 2670.445 579.445 2670.615 579.615 ;
        RECT 2670.445 524.025 2670.615 524.195 ;
        RECT 2670.445 427.465 2670.615 427.635 ;
        RECT 2670.445 339.065 2670.615 339.235 ;
        RECT 2670.445 210.205 2670.615 210.375 ;
        RECT 2670.445 137.785 2670.615 137.955 ;
      LAYER met1 ;
        RECT 2670.370 579.600 2670.690 579.660 ;
        RECT 2670.175 579.460 2670.690 579.600 ;
        RECT 2670.370 579.400 2670.690 579.460 ;
        RECT 2670.370 532.000 2670.690 532.060 ;
        RECT 2670.175 531.860 2670.690 532.000 ;
        RECT 2670.370 531.800 2670.690 531.860 ;
        RECT 2670.370 524.180 2670.690 524.240 ;
        RECT 2670.175 524.040 2670.690 524.180 ;
        RECT 2670.370 523.980 2670.690 524.040 ;
        RECT 2670.370 476.240 2670.690 476.300 ;
        RECT 2670.175 476.100 2670.690 476.240 ;
        RECT 2670.370 476.040 2670.690 476.100 ;
        RECT 2670.370 427.620 2670.690 427.680 ;
        RECT 2670.175 427.480 2670.690 427.620 ;
        RECT 2670.370 427.420 2670.690 427.480 ;
        RECT 2670.370 379.680 2670.690 379.740 ;
        RECT 2670.175 379.540 2670.690 379.680 ;
        RECT 2670.370 379.480 2670.690 379.540 ;
        RECT 2670.370 339.220 2670.690 339.280 ;
        RECT 2670.175 339.080 2670.690 339.220 ;
        RECT 2670.370 339.020 2670.690 339.080 ;
        RECT 2670.370 331.400 2670.690 331.460 ;
        RECT 2670.175 331.260 2670.690 331.400 ;
        RECT 2670.370 331.200 2670.690 331.260 ;
        RECT 2670.370 210.360 2670.690 210.420 ;
        RECT 2670.175 210.220 2670.690 210.360 ;
        RECT 2670.370 210.160 2670.690 210.220 ;
        RECT 2670.370 145.080 2670.690 145.140 ;
        RECT 2670.175 144.940 2670.690 145.080 ;
        RECT 2670.370 144.880 2670.690 144.940 ;
        RECT 2670.370 137.940 2670.690 138.000 ;
        RECT 2670.175 137.800 2670.690 137.940 ;
        RECT 2670.370 137.740 2670.690 137.800 ;
        RECT 2670.385 48.520 2670.675 48.565 ;
        RECT 2670.830 48.520 2671.150 48.580 ;
        RECT 2670.385 48.380 2671.150 48.520 ;
        RECT 2670.385 48.335 2670.675 48.380 ;
        RECT 2670.830 48.320 2671.150 48.380 ;
      LAYER via ;
        RECT 2670.400 579.400 2670.660 579.660 ;
        RECT 2670.400 531.800 2670.660 532.060 ;
        RECT 2670.400 523.980 2670.660 524.240 ;
        RECT 2670.400 476.040 2670.660 476.300 ;
        RECT 2670.400 427.420 2670.660 427.680 ;
        RECT 2670.400 379.480 2670.660 379.740 ;
        RECT 2670.400 339.020 2670.660 339.280 ;
        RECT 2670.400 331.200 2670.660 331.460 ;
        RECT 2670.400 210.160 2670.660 210.420 ;
        RECT 2670.400 144.880 2670.660 145.140 ;
        RECT 2670.400 137.740 2670.660 138.000 ;
        RECT 2670.860 48.320 2671.120 48.580 ;
      LAYER met2 ;
        RECT 1618.420 2374.290 1618.700 2377.880 ;
        RECT 1619.290 2374.290 1619.570 2374.405 ;
        RECT 1618.420 2374.150 1619.570 2374.290 ;
        RECT 1618.420 2373.880 1618.700 2374.150 ;
        RECT 1619.290 2374.035 1619.570 2374.150 ;
        RECT 2670.390 2369.955 2670.670 2370.325 ;
        RECT 2670.460 579.690 2670.600 2369.955 ;
        RECT 2670.400 579.370 2670.660 579.690 ;
        RECT 2670.400 531.770 2670.660 532.090 ;
        RECT 2670.460 524.270 2670.600 531.770 ;
        RECT 2670.400 523.950 2670.660 524.270 ;
        RECT 2670.400 476.010 2670.660 476.330 ;
        RECT 2670.460 427.710 2670.600 476.010 ;
        RECT 2670.400 427.390 2670.660 427.710 ;
        RECT 2670.400 379.450 2670.660 379.770 ;
        RECT 2670.460 339.310 2670.600 379.450 ;
        RECT 2670.400 338.990 2670.660 339.310 ;
        RECT 2670.400 331.170 2670.660 331.490 ;
        RECT 2670.460 210.450 2670.600 331.170 ;
        RECT 2670.400 210.130 2670.660 210.450 ;
        RECT 2670.400 144.850 2670.660 145.170 ;
        RECT 2670.460 138.030 2670.600 144.850 ;
        RECT 2670.400 137.710 2670.660 138.030 ;
        RECT 2670.860 48.290 2671.120 48.610 ;
        RECT 2670.920 24.890 2671.060 48.290 ;
        RECT 2670.920 24.750 2672.900 24.890 ;
        RECT 2672.760 2.400 2672.900 24.750 ;
        RECT 2672.550 -4.800 2673.110 2.400 ;
      LAYER via2 ;
        RECT 1619.290 2374.080 1619.570 2374.360 ;
        RECT 2670.390 2370.000 2670.670 2370.280 ;
      LAYER met3 ;
        RECT 1619.265 2374.380 1619.595 2374.385 ;
        RECT 1619.265 2374.370 1619.850 2374.380 ;
        RECT 1619.265 2374.070 1620.050 2374.370 ;
        RECT 1619.265 2374.060 1619.850 2374.070 ;
        RECT 1619.265 2374.055 1619.595 2374.060 ;
        RECT 1619.470 2370.290 1619.850 2370.300 ;
        RECT 2670.365 2370.290 2670.695 2370.305 ;
        RECT 1619.470 2369.990 2670.695 2370.290 ;
        RECT 1619.470 2369.980 1619.850 2369.990 ;
        RECT 2670.365 2369.975 2670.695 2369.990 ;
      LAYER via3 ;
        RECT 1619.500 2374.060 1619.820 2374.380 ;
        RECT 1619.500 2369.980 1619.820 2370.300 ;
      LAYER met4 ;
        RECT 1619.495 2374.055 1619.825 2374.385 ;
        RECT 1619.510 2370.305 1619.810 2374.055 ;
        RECT 1619.495 2369.975 1619.825 2370.305 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1771.990 2346.240 1772.310 2346.300 ;
        RECT 2684.170 2346.240 2684.490 2346.300 ;
        RECT 1771.990 2346.100 2684.490 2346.240 ;
        RECT 1771.990 2346.040 1772.310 2346.100 ;
        RECT 2684.170 2346.040 2684.490 2346.100 ;
        RECT 2684.170 9.080 2684.490 9.140 ;
        RECT 2690.610 9.080 2690.930 9.140 ;
        RECT 2684.170 8.940 2690.930 9.080 ;
        RECT 2684.170 8.880 2684.490 8.940 ;
        RECT 2690.610 8.880 2690.930 8.940 ;
      LAYER via ;
        RECT 1772.020 2346.040 1772.280 2346.300 ;
        RECT 2684.200 2346.040 2684.460 2346.300 ;
        RECT 2684.200 8.880 2684.460 9.140 ;
        RECT 2690.640 8.880 2690.900 9.140 ;
      LAYER met2 ;
        RECT 1772.010 2348.875 1772.290 2349.245 ;
        RECT 1772.080 2346.330 1772.220 2348.875 ;
        RECT 1772.020 2346.010 1772.280 2346.330 ;
        RECT 2684.200 2346.010 2684.460 2346.330 ;
        RECT 2684.260 9.170 2684.400 2346.010 ;
        RECT 2684.200 8.850 2684.460 9.170 ;
        RECT 2690.640 8.850 2690.900 9.170 ;
        RECT 2690.700 2.400 2690.840 8.850 ;
        RECT 2690.490 -4.800 2691.050 2.400 ;
      LAYER via2 ;
        RECT 1772.010 2348.920 1772.290 2349.200 ;
      LAYER met3 ;
        RECT 1755.835 2349.210 1759.835 2349.215 ;
        RECT 1771.985 2349.210 1772.315 2349.225 ;
        RECT 1755.835 2348.910 1772.315 2349.210 ;
        RECT 1755.835 2348.615 1759.835 2348.910 ;
        RECT 1771.985 2348.895 1772.315 2348.910 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1421.010 66.540 1421.330 66.600 ;
        RECT 2704.870 66.540 2705.190 66.600 ;
        RECT 1421.010 66.400 2705.190 66.540 ;
        RECT 1421.010 66.340 1421.330 66.400 ;
        RECT 2704.870 66.340 2705.190 66.400 ;
        RECT 2704.870 2.960 2705.190 3.020 ;
        RECT 2708.550 2.960 2708.870 3.020 ;
        RECT 2704.870 2.820 2708.870 2.960 ;
        RECT 2704.870 2.760 2705.190 2.820 ;
        RECT 2708.550 2.760 2708.870 2.820 ;
      LAYER via ;
        RECT 1421.040 66.340 1421.300 66.600 ;
        RECT 2704.900 66.340 2705.160 66.600 ;
        RECT 2704.900 2.760 2705.160 3.020 ;
        RECT 2708.580 2.760 2708.840 3.020 ;
      LAYER met2 ;
        RECT 1417.860 1323.690 1418.140 1327.135 ;
        RECT 1417.860 1323.550 1421.240 1323.690 ;
        RECT 1417.860 1323.135 1418.140 1323.550 ;
        RECT 1421.100 66.630 1421.240 1323.550 ;
        RECT 1421.040 66.310 1421.300 66.630 ;
        RECT 2704.900 66.310 2705.160 66.630 ;
        RECT 2704.960 3.050 2705.100 66.310 ;
        RECT 2704.900 2.730 2705.160 3.050 ;
        RECT 2708.580 2.730 2708.840 3.050 ;
        RECT 2708.640 2.400 2708.780 2.730 ;
        RECT 2708.430 -4.800 2708.990 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1772.910 1663.180 1773.230 1663.240 ;
        RECT 2342.390 1663.180 2342.710 1663.240 ;
        RECT 1772.910 1663.040 2342.710 1663.180 ;
        RECT 1772.910 1662.980 1773.230 1663.040 ;
        RECT 2342.390 1662.980 2342.710 1663.040 ;
        RECT 2342.390 18.600 2342.710 18.660 ;
        RECT 2726.490 18.600 2726.810 18.660 ;
        RECT 2342.390 18.460 2726.810 18.600 ;
        RECT 2342.390 18.400 2342.710 18.460 ;
        RECT 2726.490 18.400 2726.810 18.460 ;
      LAYER via ;
        RECT 1772.940 1662.980 1773.200 1663.240 ;
        RECT 2342.420 1662.980 2342.680 1663.240 ;
        RECT 2342.420 18.400 2342.680 18.660 ;
        RECT 2726.520 18.400 2726.780 18.660 ;
      LAYER met2 ;
        RECT 1772.930 1664.795 1773.210 1665.165 ;
        RECT 1773.000 1663.270 1773.140 1664.795 ;
        RECT 1772.940 1662.950 1773.200 1663.270 ;
        RECT 2342.420 1662.950 2342.680 1663.270 ;
        RECT 2342.480 18.690 2342.620 1662.950 ;
        RECT 2342.420 18.370 2342.680 18.690 ;
        RECT 2726.520 18.370 2726.780 18.690 ;
        RECT 2726.580 2.400 2726.720 18.370 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
      LAYER via2 ;
        RECT 1772.930 1664.840 1773.210 1665.120 ;
      LAYER met3 ;
        RECT 1755.835 1665.130 1759.835 1665.135 ;
        RECT 1772.905 1665.130 1773.235 1665.145 ;
        RECT 1755.835 1664.830 1773.235 1665.130 ;
        RECT 1755.835 1664.535 1759.835 1664.830 ;
        RECT 1772.905 1664.815 1773.235 1664.830 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1772.910 1801.220 1773.230 1801.280 ;
        RECT 2356.190 1801.220 2356.510 1801.280 ;
        RECT 1772.910 1801.080 2356.510 1801.220 ;
        RECT 1772.910 1801.020 1773.230 1801.080 ;
        RECT 2356.190 1801.020 2356.510 1801.080 ;
        RECT 2356.190 18.260 2356.510 18.320 ;
        RECT 2744.430 18.260 2744.750 18.320 ;
        RECT 2356.190 18.120 2744.750 18.260 ;
        RECT 2356.190 18.060 2356.510 18.120 ;
        RECT 2744.430 18.060 2744.750 18.120 ;
      LAYER via ;
        RECT 1772.940 1801.020 1773.200 1801.280 ;
        RECT 2356.220 1801.020 2356.480 1801.280 ;
        RECT 2356.220 18.060 2356.480 18.320 ;
        RECT 2744.460 18.060 2744.720 18.320 ;
      LAYER met2 ;
        RECT 1772.940 1801.165 1773.200 1801.310 ;
        RECT 1772.930 1800.795 1773.210 1801.165 ;
        RECT 2356.220 1800.990 2356.480 1801.310 ;
        RECT 2356.280 18.350 2356.420 1800.990 ;
        RECT 2356.220 18.030 2356.480 18.350 ;
        RECT 2744.460 18.030 2744.720 18.350 ;
        RECT 2744.520 2.400 2744.660 18.030 ;
        RECT 2744.310 -4.800 2744.870 2.400 ;
      LAYER via2 ;
        RECT 1772.930 1800.840 1773.210 1801.120 ;
      LAYER met3 ;
        RECT 1755.835 1801.130 1759.835 1801.135 ;
        RECT 1772.905 1801.130 1773.235 1801.145 ;
        RECT 1755.835 1800.830 1773.235 1801.130 ;
        RECT 1755.835 1800.535 1759.835 1800.830 ;
        RECT 1772.905 1800.815 1773.235 1800.830 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2760.090 886.195 2760.370 886.565 ;
        RECT 2760.160 17.410 2760.300 886.195 ;
        RECT 2760.160 17.270 2762.140 17.410 ;
        RECT 2762.000 2.400 2762.140 17.270 ;
        RECT 2761.790 -4.800 2762.350 2.400 ;
      LAYER via2 ;
        RECT 2760.090 886.240 2760.370 886.520 ;
      LAYER met3 ;
        RECT 704.070 1412.170 704.450 1412.180 ;
        RECT 715.810 1412.170 719.810 1412.175 ;
        RECT 704.070 1411.870 719.810 1412.170 ;
        RECT 704.070 1411.860 704.450 1411.870 ;
        RECT 715.810 1411.575 719.810 1411.870 ;
        RECT 704.070 886.530 704.450 886.540 ;
        RECT 2760.065 886.530 2760.395 886.545 ;
        RECT 704.070 886.230 2760.395 886.530 ;
        RECT 704.070 886.220 704.450 886.230 ;
        RECT 2760.065 886.215 2760.395 886.230 ;
      LAYER via3 ;
        RECT 704.100 1411.860 704.420 1412.180 ;
        RECT 704.100 886.220 704.420 886.540 ;
      LAYER met4 ;
        RECT 704.095 1411.855 704.425 1412.185 ;
        RECT 704.110 886.545 704.410 1411.855 ;
        RECT 704.095 886.215 704.425 886.545 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 704.405 1310.785 704.575 1362.295 ;
        RECT 759.605 13.685 759.775 15.215 ;
      LAYER mcon ;
        RECT 704.405 1362.125 704.575 1362.295 ;
        RECT 759.605 15.045 759.775 15.215 ;
      LAYER met1 ;
        RECT 704.345 1362.280 704.635 1362.325 ;
        RECT 707.090 1362.280 707.410 1362.340 ;
        RECT 704.345 1362.140 707.410 1362.280 ;
        RECT 704.345 1362.095 704.635 1362.140 ;
        RECT 707.090 1362.080 707.410 1362.140 ;
        RECT 704.345 1310.940 704.635 1310.985 ;
        RECT 727.790 1310.940 728.110 1311.000 ;
        RECT 704.345 1310.800 728.110 1310.940 ;
        RECT 704.345 1310.755 704.635 1310.800 ;
        RECT 727.790 1310.740 728.110 1310.800 ;
        RECT 759.545 15.200 759.835 15.245 ;
        RECT 786.670 15.200 786.990 15.260 ;
        RECT 759.545 15.060 786.990 15.200 ;
        RECT 759.545 15.015 759.835 15.060 ;
        RECT 786.670 15.000 786.990 15.060 ;
        RECT 800.470 14.860 800.790 14.920 ;
        RECT 835.430 14.860 835.750 14.920 ;
        RECT 800.470 14.720 835.750 14.860 ;
        RECT 800.470 14.660 800.790 14.720 ;
        RECT 835.430 14.660 835.750 14.720 ;
        RECT 727.790 14.180 728.110 14.240 ;
        RECT 727.790 14.040 741.820 14.180 ;
        RECT 727.790 13.980 728.110 14.040 ;
        RECT 741.680 13.840 741.820 14.040 ;
        RECT 759.545 13.840 759.835 13.885 ;
        RECT 741.680 13.700 759.835 13.840 ;
        RECT 759.545 13.655 759.835 13.700 ;
      LAYER via ;
        RECT 707.120 1362.080 707.380 1362.340 ;
        RECT 727.820 1310.740 728.080 1311.000 ;
        RECT 786.700 15.000 786.960 15.260 ;
        RECT 800.500 14.660 800.760 14.920 ;
        RECT 835.460 14.660 835.720 14.920 ;
        RECT 727.820 13.980 728.080 14.240 ;
      LAYER met2 ;
        RECT 707.110 2061.915 707.390 2062.285 ;
        RECT 707.180 1362.370 707.320 2061.915 ;
        RECT 707.120 1362.050 707.380 1362.370 ;
        RECT 727.820 1310.710 728.080 1311.030 ;
        RECT 727.880 14.270 728.020 1310.710 ;
        RECT 786.700 14.970 786.960 15.290 ;
        RECT 727.820 13.950 728.080 14.270 ;
        RECT 786.760 14.125 786.900 14.970 ;
        RECT 800.500 14.630 800.760 14.950 ;
        RECT 835.460 14.630 835.720 14.950 ;
        RECT 800.560 14.125 800.700 14.630 ;
        RECT 786.690 13.755 786.970 14.125 ;
        RECT 800.490 13.755 800.770 14.125 ;
        RECT 835.520 2.400 835.660 14.630 ;
        RECT 835.310 -4.800 835.870 2.400 ;
      LAYER via2 ;
        RECT 707.110 2061.960 707.390 2062.240 ;
        RECT 786.690 13.800 786.970 14.080 ;
        RECT 800.490 13.800 800.770 14.080 ;
      LAYER met3 ;
        RECT 707.085 2062.250 707.415 2062.265 ;
        RECT 715.810 2062.250 719.810 2062.255 ;
        RECT 707.085 2061.950 719.810 2062.250 ;
        RECT 707.085 2061.935 707.415 2061.950 ;
        RECT 715.810 2061.655 719.810 2061.950 ;
        RECT 786.665 14.090 786.995 14.105 ;
        RECT 800.465 14.090 800.795 14.105 ;
        RECT 786.665 13.790 800.795 14.090 ;
        RECT 786.665 13.775 786.995 13.790 ;
        RECT 800.465 13.775 800.795 13.790 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2773.870 18.260 2774.190 18.320 ;
        RECT 2779.850 18.260 2780.170 18.320 ;
        RECT 2773.870 18.120 2780.170 18.260 ;
        RECT 2773.870 18.060 2774.190 18.120 ;
        RECT 2779.850 18.060 2780.170 18.120 ;
      LAYER via ;
        RECT 2773.900 18.060 2774.160 18.320 ;
        RECT 2779.880 18.060 2780.140 18.320 ;
      LAYER met2 ;
        RECT 1145.490 2380.155 1145.770 2380.525 ;
        RECT 1197.470 2380.155 1197.750 2380.525 ;
        RECT 1306.950 2380.155 1307.230 2380.525 ;
        RECT 1126.220 2374.290 1126.500 2377.880 ;
        RECT 1145.560 2374.405 1145.700 2380.155 ;
        RECT 1197.540 2374.405 1197.680 2380.155 ;
        RECT 1307.020 2374.405 1307.160 2380.155 ;
        RECT 1127.550 2374.290 1127.830 2374.405 ;
        RECT 1126.220 2374.150 1127.830 2374.290 ;
        RECT 1126.220 2373.880 1126.500 2374.150 ;
        RECT 1127.550 2374.035 1127.830 2374.150 ;
        RECT 1145.490 2374.035 1145.770 2374.405 ;
        RECT 1197.470 2374.035 1197.750 2374.405 ;
        RECT 1306.950 2374.035 1307.230 2374.405 ;
        RECT 2773.890 2374.035 2774.170 2374.405 ;
        RECT 2773.960 18.350 2774.100 2374.035 ;
        RECT 2773.900 18.030 2774.160 18.350 ;
        RECT 2779.880 18.030 2780.140 18.350 ;
        RECT 2779.940 2.400 2780.080 18.030 ;
        RECT 2779.730 -4.800 2780.290 2.400 ;
      LAYER via2 ;
        RECT 1145.490 2380.200 1145.770 2380.480 ;
        RECT 1197.470 2380.200 1197.750 2380.480 ;
        RECT 1306.950 2380.200 1307.230 2380.480 ;
        RECT 1127.550 2374.080 1127.830 2374.360 ;
        RECT 1145.490 2374.080 1145.770 2374.360 ;
        RECT 1197.470 2374.080 1197.750 2374.360 ;
        RECT 1306.950 2374.080 1307.230 2374.360 ;
        RECT 2773.890 2374.080 2774.170 2374.360 ;
      LAYER met3 ;
        RECT 1145.465 2380.490 1145.795 2380.505 ;
        RECT 1197.445 2380.490 1197.775 2380.505 ;
        RECT 1145.465 2380.190 1197.775 2380.490 ;
        RECT 1145.465 2380.175 1145.795 2380.190 ;
        RECT 1197.445 2380.175 1197.775 2380.190 ;
        RECT 1242.270 2380.490 1242.650 2380.500 ;
        RECT 1306.925 2380.490 1307.255 2380.505 ;
        RECT 1242.270 2380.190 1307.255 2380.490 ;
        RECT 1242.270 2380.180 1242.650 2380.190 ;
        RECT 1306.925 2380.175 1307.255 2380.190 ;
        RECT 1127.525 2374.370 1127.855 2374.385 ;
        RECT 1145.465 2374.370 1145.795 2374.385 ;
        RECT 1127.525 2374.070 1145.795 2374.370 ;
        RECT 1127.525 2374.055 1127.855 2374.070 ;
        RECT 1145.465 2374.055 1145.795 2374.070 ;
        RECT 1197.445 2374.370 1197.775 2374.385 ;
        RECT 1242.270 2374.370 1242.650 2374.380 ;
        RECT 1197.445 2374.070 1242.650 2374.370 ;
        RECT 1197.445 2374.055 1197.775 2374.070 ;
        RECT 1242.270 2374.060 1242.650 2374.070 ;
        RECT 1306.925 2374.370 1307.255 2374.385 ;
        RECT 2773.865 2374.370 2774.195 2374.385 ;
        RECT 1306.925 2374.070 1618.890 2374.370 ;
        RECT 1306.925 2374.055 1307.255 2374.070 ;
        RECT 1618.590 2373.690 1618.890 2374.070 ;
        RECT 1620.430 2374.070 1740.330 2374.370 ;
        RECT 1620.430 2373.690 1620.730 2374.070 ;
        RECT 1618.590 2373.390 1620.730 2373.690 ;
        RECT 1740.030 2373.690 1740.330 2374.070 ;
        RECT 1750.150 2374.070 2774.195 2374.370 ;
        RECT 1750.150 2373.690 1750.450 2374.070 ;
        RECT 2773.865 2374.055 2774.195 2374.070 ;
        RECT 1740.030 2373.390 1750.450 2373.690 ;
      LAYER via3 ;
        RECT 1242.300 2380.180 1242.620 2380.500 ;
        RECT 1242.300 2374.060 1242.620 2374.380 ;
      LAYER met4 ;
        RECT 1242.295 2380.175 1242.625 2380.505 ;
        RECT 1242.310 2374.385 1242.610 2380.175 ;
        RECT 1242.295 2374.055 1242.625 2374.385 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 884.650 2375.140 884.970 2375.200 ;
        RECT 931.570 2375.140 931.890 2375.200 ;
        RECT 884.650 2375.000 931.890 2375.140 ;
        RECT 884.650 2374.940 884.970 2375.000 ;
        RECT 931.570 2374.940 931.890 2375.000 ;
      LAYER via ;
        RECT 884.680 2374.940 884.940 2375.200 ;
        RECT 931.600 2374.940 931.860 2375.200 ;
      LAYER met2 ;
        RECT 883.340 2374.970 883.620 2377.880 ;
        RECT 931.590 2376.075 931.870 2376.445 ;
        RECT 2794.590 2376.075 2794.870 2376.445 ;
        RECT 931.660 2375.230 931.800 2376.075 ;
        RECT 884.680 2374.970 884.940 2375.230 ;
        RECT 883.340 2374.910 884.940 2374.970 ;
        RECT 931.600 2374.910 931.860 2375.230 ;
        RECT 883.340 2374.830 884.880 2374.910 ;
        RECT 883.340 2373.880 883.620 2374.830 ;
        RECT 2794.660 17.410 2794.800 2376.075 ;
        RECT 2794.660 17.270 2798.020 17.410 ;
        RECT 2797.880 2.400 2798.020 17.270 ;
        RECT 2797.670 -4.800 2798.230 2.400 ;
      LAYER via2 ;
        RECT 931.590 2376.120 931.870 2376.400 ;
        RECT 2794.590 2376.120 2794.870 2376.400 ;
      LAYER met3 ;
        RECT 931.565 2376.410 931.895 2376.425 ;
        RECT 2794.565 2376.410 2794.895 2376.425 ;
        RECT 931.565 2376.110 2794.895 2376.410 ;
        RECT 931.565 2376.095 931.895 2376.110 ;
        RECT 2794.565 2376.095 2794.895 2376.110 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 717.745 1543.005 717.915 1589.415 ;
        RECT 718.665 1339.005 718.835 1373.855 ;
      LAYER mcon ;
        RECT 717.745 1589.245 717.915 1589.415 ;
        RECT 718.665 1373.685 718.835 1373.855 ;
      LAYER met1 ;
        RECT 717.685 1589.400 717.975 1589.445 ;
        RECT 718.590 1589.400 718.910 1589.460 ;
        RECT 717.685 1589.260 718.910 1589.400 ;
        RECT 717.685 1589.215 717.975 1589.260 ;
        RECT 718.590 1589.200 718.910 1589.260 ;
        RECT 717.685 1543.160 717.975 1543.205 ;
        RECT 718.590 1543.160 718.910 1543.220 ;
        RECT 717.685 1543.020 718.910 1543.160 ;
        RECT 717.685 1542.975 717.975 1543.020 ;
        RECT 718.590 1542.960 718.910 1543.020 ;
        RECT 717.210 1373.840 717.530 1373.900 ;
        RECT 718.605 1373.840 718.895 1373.885 ;
        RECT 717.210 1373.700 718.895 1373.840 ;
        RECT 717.210 1373.640 717.530 1373.700 ;
        RECT 718.605 1373.655 718.895 1373.700 ;
        RECT 718.605 1339.160 718.895 1339.205 ;
        RECT 719.970 1339.160 720.290 1339.220 ;
        RECT 718.605 1339.020 720.290 1339.160 ;
        RECT 718.605 1338.975 718.895 1339.020 ;
        RECT 719.970 1338.960 720.290 1339.020 ;
      LAYER via ;
        RECT 718.620 1589.200 718.880 1589.460 ;
        RECT 718.620 1542.960 718.880 1543.220 ;
        RECT 717.240 1373.640 717.500 1373.900 ;
        RECT 720.000 1338.960 720.260 1339.220 ;
      LAYER met2 ;
        RECT 718.610 1589.315 718.890 1589.685 ;
        RECT 718.620 1589.170 718.880 1589.315 ;
        RECT 718.620 1542.930 718.880 1543.250 ;
        RECT 718.680 1542.085 718.820 1542.930 ;
        RECT 718.610 1541.715 718.890 1542.085 ;
        RECT 717.230 1373.755 717.510 1374.125 ;
        RECT 717.240 1373.610 717.500 1373.755 ;
        RECT 720.000 1338.930 720.260 1339.250 ;
        RECT 720.060 1326.525 720.200 1338.930 ;
        RECT 719.990 1326.155 720.270 1326.525 ;
        RECT 724.130 1283.995 724.410 1284.365 ;
        RECT 724.200 1249.685 724.340 1283.995 ;
        RECT 724.130 1249.315 724.410 1249.685 ;
        RECT 723.210 1139.155 723.490 1139.525 ;
        RECT 723.280 1090.565 723.420 1139.155 ;
        RECT 723.210 1090.195 723.490 1090.565 ;
        RECT 723.670 1042.595 723.950 1042.965 ;
        RECT 723.740 1007.605 723.880 1042.595 ;
        RECT 723.670 1007.235 723.950 1007.605 ;
        RECT 723.670 848.115 723.950 848.485 ;
        RECT 723.740 773.005 723.880 848.115 ;
        RECT 723.670 772.635 723.950 773.005 ;
        RECT 723.670 750.875 723.950 751.245 ;
        RECT 723.740 676.445 723.880 750.875 ;
        RECT 723.670 676.075 723.950 676.445 ;
        RECT 723.210 529.875 723.490 530.245 ;
        RECT 723.280 494.885 723.420 529.875 ;
        RECT 723.210 494.515 723.490 494.885 ;
        RECT 723.670 467.995 723.950 468.365 ;
        RECT 723.740 421.445 723.880 467.995 ;
        RECT 723.670 421.075 723.950 421.445 ;
        RECT 723.670 269.435 723.950 269.805 ;
        RECT 723.740 235.125 723.880 269.435 ;
        RECT 723.670 234.755 723.950 235.125 ;
        RECT 723.670 221.835 723.950 222.205 ;
        RECT 723.740 194.325 723.880 221.835 ;
        RECT 723.670 193.955 723.950 194.325 ;
        RECT 723.210 144.315 723.490 144.685 ;
        RECT 723.280 97.085 723.420 144.315 ;
        RECT 723.210 96.715 723.490 97.085 ;
        RECT 723.670 95.355 723.950 95.725 ;
        RECT 723.740 76.005 723.880 95.355 ;
        RECT 723.670 75.635 723.950 76.005 ;
        RECT 724.590 62.035 724.870 62.405 ;
        RECT 724.660 44.725 724.800 62.035 ;
        RECT 724.590 44.355 724.870 44.725 ;
        RECT 2815.750 44.355 2816.030 44.725 ;
        RECT 2815.820 2.400 2815.960 44.355 ;
        RECT 2815.610 -4.800 2816.170 2.400 ;
      LAYER via2 ;
        RECT 718.610 1589.360 718.890 1589.640 ;
        RECT 718.610 1541.760 718.890 1542.040 ;
        RECT 717.230 1373.800 717.510 1374.080 ;
        RECT 719.990 1326.200 720.270 1326.480 ;
        RECT 724.130 1284.040 724.410 1284.320 ;
        RECT 724.130 1249.360 724.410 1249.640 ;
        RECT 723.210 1139.200 723.490 1139.480 ;
        RECT 723.210 1090.240 723.490 1090.520 ;
        RECT 723.670 1042.640 723.950 1042.920 ;
        RECT 723.670 1007.280 723.950 1007.560 ;
        RECT 723.670 848.160 723.950 848.440 ;
        RECT 723.670 772.680 723.950 772.960 ;
        RECT 723.670 750.920 723.950 751.200 ;
        RECT 723.670 676.120 723.950 676.400 ;
        RECT 723.210 529.920 723.490 530.200 ;
        RECT 723.210 494.560 723.490 494.840 ;
        RECT 723.670 468.040 723.950 468.320 ;
        RECT 723.670 421.120 723.950 421.400 ;
        RECT 723.670 269.480 723.950 269.760 ;
        RECT 723.670 234.800 723.950 235.080 ;
        RECT 723.670 221.880 723.950 222.160 ;
        RECT 723.670 194.000 723.950 194.280 ;
        RECT 723.210 144.360 723.490 144.640 ;
        RECT 723.210 96.760 723.490 97.040 ;
        RECT 723.670 95.400 723.950 95.680 ;
        RECT 723.670 75.680 723.950 75.960 ;
        RECT 724.590 62.080 724.870 62.360 ;
        RECT 724.590 44.400 724.870 44.680 ;
        RECT 2815.750 44.400 2816.030 44.680 ;
      LAYER met3 ;
        RECT 715.810 1616.935 719.810 1617.535 ;
        RECT 718.830 1614.820 719.130 1616.935 ;
        RECT 718.790 1614.500 719.170 1614.820 ;
        RECT 718.585 1589.660 718.915 1589.665 ;
        RECT 718.585 1589.650 719.170 1589.660 ;
        RECT 718.360 1589.350 719.170 1589.650 ;
        RECT 718.585 1589.340 719.170 1589.350 ;
        RECT 718.585 1589.335 718.915 1589.340 ;
        RECT 718.585 1542.060 718.915 1542.065 ;
        RECT 718.585 1542.050 719.170 1542.060 ;
        RECT 718.360 1541.750 719.170 1542.050 ;
        RECT 718.585 1541.740 719.170 1541.750 ;
        RECT 718.585 1541.735 718.915 1541.740 ;
        RECT 717.205 1374.090 717.535 1374.105 ;
        RECT 718.790 1374.090 719.170 1374.100 ;
        RECT 717.205 1373.790 719.170 1374.090 ;
        RECT 717.205 1373.775 717.535 1373.790 ;
        RECT 718.790 1373.780 719.170 1373.790 ;
        RECT 719.965 1326.490 720.295 1326.505 ;
        RECT 723.390 1326.490 723.770 1326.500 ;
        RECT 719.965 1326.190 723.770 1326.490 ;
        RECT 719.965 1326.175 720.295 1326.190 ;
        RECT 723.390 1326.180 723.770 1326.190 ;
        RECT 724.105 1284.340 724.435 1284.345 ;
        RECT 724.105 1284.330 724.690 1284.340 ;
        RECT 723.880 1284.030 724.690 1284.330 ;
        RECT 724.105 1284.020 724.690 1284.030 ;
        RECT 724.105 1284.015 724.435 1284.020 ;
        RECT 724.105 1249.660 724.435 1249.665 ;
        RECT 724.105 1249.650 724.690 1249.660 ;
        RECT 724.105 1249.350 724.890 1249.650 ;
        RECT 724.105 1249.340 724.690 1249.350 ;
        RECT 724.105 1249.335 724.435 1249.340 ;
        RECT 723.390 1248.970 723.770 1248.980 ;
        RECT 725.230 1248.970 725.610 1248.980 ;
        RECT 723.390 1248.670 725.610 1248.970 ;
        RECT 723.390 1248.660 723.770 1248.670 ;
        RECT 725.230 1248.660 725.610 1248.670 ;
        RECT 723.390 1187.090 723.770 1187.100 ;
        RECT 725.230 1187.090 725.610 1187.100 ;
        RECT 723.390 1186.790 725.610 1187.090 ;
        RECT 723.390 1186.780 723.770 1186.790 ;
        RECT 725.230 1186.780 725.610 1186.790 ;
        RECT 723.185 1139.500 723.515 1139.505 ;
        RECT 723.185 1139.490 723.770 1139.500 ;
        RECT 722.960 1139.190 723.770 1139.490 ;
        RECT 723.185 1139.180 723.770 1139.190 ;
        RECT 723.185 1139.175 723.515 1139.180 ;
        RECT 723.185 1090.540 723.515 1090.545 ;
        RECT 723.185 1090.530 723.770 1090.540 ;
        RECT 723.185 1090.230 723.970 1090.530 ;
        RECT 723.185 1090.220 723.770 1090.230 ;
        RECT 723.185 1090.215 723.515 1090.220 ;
        RECT 723.645 1042.940 723.975 1042.945 ;
        RECT 723.390 1042.930 723.975 1042.940 ;
        RECT 723.190 1042.630 723.975 1042.930 ;
        RECT 723.390 1042.620 723.975 1042.630 ;
        RECT 723.645 1042.615 723.975 1042.620 ;
        RECT 723.645 1007.570 723.975 1007.585 ;
        RECT 724.310 1007.570 724.690 1007.580 ;
        RECT 723.645 1007.270 724.690 1007.570 ;
        RECT 723.645 1007.255 723.975 1007.270 ;
        RECT 724.310 1007.260 724.690 1007.270 ;
        RECT 724.310 994.650 724.690 994.660 ;
        RECT 723.430 994.350 724.690 994.650 ;
        RECT 723.430 993.300 723.730 994.350 ;
        RECT 724.310 994.340 724.690 994.350 ;
        RECT 723.390 992.980 723.770 993.300 ;
        RECT 723.645 848.450 723.975 848.465 ;
        RECT 724.310 848.450 724.690 848.460 ;
        RECT 723.645 848.150 724.690 848.450 ;
        RECT 723.645 848.135 723.975 848.150 ;
        RECT 724.310 848.140 724.690 848.150 ;
        RECT 723.645 772.980 723.975 772.985 ;
        RECT 723.390 772.970 723.975 772.980 ;
        RECT 723.190 772.670 723.975 772.970 ;
        RECT 723.390 772.660 723.975 772.670 ;
        RECT 723.645 772.655 723.975 772.660 ;
        RECT 723.645 751.220 723.975 751.225 ;
        RECT 723.390 751.210 723.975 751.220 ;
        RECT 723.390 750.910 724.200 751.210 ;
        RECT 723.390 750.900 723.975 750.910 ;
        RECT 723.645 750.895 723.975 750.900 ;
        RECT 723.645 676.420 723.975 676.425 ;
        RECT 723.390 676.410 723.975 676.420 ;
        RECT 723.190 676.110 723.975 676.410 ;
        RECT 723.390 676.100 723.975 676.110 ;
        RECT 723.645 676.095 723.975 676.100 ;
        RECT 724.310 608.410 724.690 608.420 ;
        RECT 723.430 608.110 724.690 608.410 ;
        RECT 723.430 607.740 723.730 608.110 ;
        RECT 724.310 608.100 724.690 608.110 ;
        RECT 723.390 607.420 723.770 607.740 ;
        RECT 723.390 531.090 723.770 531.410 ;
        RECT 723.430 530.225 723.730 531.090 ;
        RECT 723.185 529.910 723.730 530.225 ;
        RECT 723.185 529.895 723.515 529.910 ;
        RECT 723.185 494.860 723.515 494.865 ;
        RECT 723.185 494.850 723.770 494.860 ;
        RECT 722.960 494.550 723.770 494.850 ;
        RECT 723.185 494.540 723.770 494.550 ;
        RECT 723.185 494.535 723.515 494.540 ;
        RECT 723.390 468.700 723.770 469.020 ;
        RECT 723.430 468.345 723.730 468.700 ;
        RECT 723.430 468.030 723.975 468.345 ;
        RECT 723.645 468.015 723.975 468.030 ;
        RECT 723.645 421.410 723.975 421.425 ;
        RECT 724.310 421.410 724.690 421.420 ;
        RECT 723.645 421.110 724.690 421.410 ;
        RECT 723.645 421.095 723.975 421.110 ;
        RECT 724.310 421.100 724.690 421.110 ;
        RECT 725.230 318.730 725.610 318.740 ;
        RECT 723.430 318.430 725.610 318.730 ;
        RECT 723.430 318.060 723.730 318.430 ;
        RECT 725.230 318.420 725.610 318.430 ;
        RECT 723.390 317.740 723.770 318.060 ;
        RECT 723.645 269.780 723.975 269.785 ;
        RECT 723.390 269.770 723.975 269.780 ;
        RECT 723.190 269.470 723.975 269.770 ;
        RECT 723.390 269.460 723.975 269.470 ;
        RECT 723.645 269.455 723.975 269.460 ;
        RECT 723.645 235.090 723.975 235.105 ;
        RECT 725.230 235.090 725.610 235.100 ;
        RECT 723.645 234.790 725.610 235.090 ;
        RECT 723.645 234.775 723.975 234.790 ;
        RECT 725.230 234.780 725.610 234.790 ;
        RECT 723.645 222.170 723.975 222.185 ;
        RECT 725.230 222.170 725.610 222.180 ;
        RECT 723.645 221.870 725.610 222.170 ;
        RECT 723.645 221.855 723.975 221.870 ;
        RECT 725.230 221.860 725.610 221.870 ;
        RECT 723.645 194.290 723.975 194.305 ;
        RECT 723.430 193.975 723.975 194.290 ;
        RECT 723.430 193.620 723.730 193.975 ;
        RECT 723.390 193.300 723.770 193.620 ;
        RECT 723.185 144.660 723.515 144.665 ;
        RECT 723.185 144.650 723.770 144.660 ;
        RECT 722.960 144.350 723.770 144.650 ;
        RECT 723.185 144.340 723.770 144.350 ;
        RECT 723.185 144.335 723.515 144.340 ;
        RECT 723.185 97.060 723.515 97.065 ;
        RECT 723.185 97.050 723.770 97.060 ;
        RECT 722.960 96.750 723.770 97.050 ;
        RECT 723.185 96.740 723.770 96.750 ;
        RECT 723.185 96.735 723.515 96.740 ;
        RECT 723.645 95.700 723.975 95.705 ;
        RECT 723.390 95.690 723.975 95.700 ;
        RECT 723.190 95.390 723.975 95.690 ;
        RECT 723.390 95.380 723.975 95.390 ;
        RECT 723.645 95.375 723.975 95.380 ;
        RECT 723.645 75.980 723.975 75.985 ;
        RECT 723.390 75.970 723.975 75.980 ;
        RECT 723.390 75.670 724.200 75.970 ;
        RECT 723.390 75.660 723.975 75.670 ;
        RECT 723.645 75.655 723.975 75.660 ;
        RECT 724.565 62.380 724.895 62.385 ;
        RECT 724.310 62.370 724.895 62.380 ;
        RECT 724.310 62.070 725.120 62.370 ;
        RECT 724.310 62.060 724.895 62.070 ;
        RECT 724.565 62.055 724.895 62.060 ;
        RECT 724.565 44.690 724.895 44.705 ;
        RECT 2815.725 44.690 2816.055 44.705 ;
        RECT 724.565 44.390 2816.055 44.690 ;
        RECT 724.565 44.375 724.895 44.390 ;
        RECT 2815.725 44.375 2816.055 44.390 ;
      LAYER via3 ;
        RECT 718.820 1614.500 719.140 1614.820 ;
        RECT 718.820 1589.340 719.140 1589.660 ;
        RECT 718.820 1541.740 719.140 1542.060 ;
        RECT 718.820 1373.780 719.140 1374.100 ;
        RECT 723.420 1326.180 723.740 1326.500 ;
        RECT 724.340 1284.020 724.660 1284.340 ;
        RECT 724.340 1249.340 724.660 1249.660 ;
        RECT 723.420 1248.660 723.740 1248.980 ;
        RECT 725.260 1248.660 725.580 1248.980 ;
        RECT 723.420 1186.780 723.740 1187.100 ;
        RECT 725.260 1186.780 725.580 1187.100 ;
        RECT 723.420 1139.180 723.740 1139.500 ;
        RECT 723.420 1090.220 723.740 1090.540 ;
        RECT 723.420 1042.620 723.740 1042.940 ;
        RECT 724.340 1007.260 724.660 1007.580 ;
        RECT 724.340 994.340 724.660 994.660 ;
        RECT 723.420 992.980 723.740 993.300 ;
        RECT 724.340 848.140 724.660 848.460 ;
        RECT 723.420 772.660 723.740 772.980 ;
        RECT 723.420 750.900 723.740 751.220 ;
        RECT 723.420 676.100 723.740 676.420 ;
        RECT 724.340 608.100 724.660 608.420 ;
        RECT 723.420 607.420 723.740 607.740 ;
        RECT 723.420 531.090 723.740 531.410 ;
        RECT 723.420 494.540 723.740 494.860 ;
        RECT 723.420 468.700 723.740 469.020 ;
        RECT 724.340 421.100 724.660 421.420 ;
        RECT 725.260 318.420 725.580 318.740 ;
        RECT 723.420 317.740 723.740 318.060 ;
        RECT 723.420 269.460 723.740 269.780 ;
        RECT 725.260 234.780 725.580 235.100 ;
        RECT 725.260 221.860 725.580 222.180 ;
        RECT 723.420 193.300 723.740 193.620 ;
        RECT 723.420 144.340 723.740 144.660 ;
        RECT 723.420 96.740 723.740 97.060 ;
        RECT 723.420 95.380 723.740 95.700 ;
        RECT 723.420 75.660 723.740 75.980 ;
        RECT 724.340 62.060 724.660 62.380 ;
      LAYER met4 ;
        RECT 718.815 1614.495 719.145 1614.825 ;
        RECT 718.830 1589.665 719.130 1614.495 ;
        RECT 718.815 1589.335 719.145 1589.665 ;
        RECT 718.815 1542.050 719.145 1542.065 ;
        RECT 718.815 1541.750 726.490 1542.050 ;
        RECT 718.815 1541.735 719.145 1541.750 ;
        RECT 726.190 1494.890 726.490 1541.750 ;
        RECT 720.230 1493.710 721.410 1494.890 ;
        RECT 725.750 1493.710 726.930 1494.890 ;
        RECT 720.670 1489.690 720.970 1493.710 ;
        RECT 720.670 1489.390 721.890 1489.690 ;
        RECT 721.590 1480.850 721.890 1489.390 ;
        RECT 721.590 1480.550 724.650 1480.850 ;
        RECT 724.350 1419.650 724.650 1480.550 ;
        RECT 722.510 1419.350 724.650 1419.650 ;
        RECT 722.510 1389.050 722.810 1419.350 ;
        RECT 720.670 1388.750 722.810 1389.050 ;
        RECT 720.670 1378.850 720.970 1388.750 ;
        RECT 718.830 1378.550 720.970 1378.850 ;
        RECT 718.830 1374.105 719.130 1378.550 ;
        RECT 718.815 1373.775 719.145 1374.105 ;
        RECT 723.415 1326.175 723.745 1326.505 ;
        RECT 723.430 1321.050 723.730 1326.175 ;
        RECT 723.430 1320.750 724.650 1321.050 ;
        RECT 724.350 1284.345 724.650 1320.750 ;
        RECT 724.335 1284.015 724.665 1284.345 ;
        RECT 724.335 1249.650 724.665 1249.665 ;
        RECT 723.430 1249.350 724.665 1249.650 ;
        RECT 723.430 1248.985 723.730 1249.350 ;
        RECT 724.335 1249.335 724.665 1249.350 ;
        RECT 723.415 1248.655 723.745 1248.985 ;
        RECT 725.255 1248.655 725.585 1248.985 ;
        RECT 725.270 1187.105 725.570 1248.655 ;
        RECT 723.415 1186.775 723.745 1187.105 ;
        RECT 725.255 1186.775 725.585 1187.105 ;
        RECT 723.430 1139.505 723.730 1186.775 ;
        RECT 723.415 1139.175 723.745 1139.505 ;
        RECT 723.415 1090.215 723.745 1090.545 ;
        RECT 723.430 1042.945 723.730 1090.215 ;
        RECT 723.415 1042.615 723.745 1042.945 ;
        RECT 724.335 1007.255 724.665 1007.585 ;
        RECT 724.350 994.665 724.650 1007.255 ;
        RECT 724.335 994.335 724.665 994.665 ;
        RECT 723.415 992.975 723.745 993.305 ;
        RECT 723.430 848.450 723.730 992.975 ;
        RECT 724.335 848.450 724.665 848.465 ;
        RECT 723.430 848.150 724.665 848.450 ;
        RECT 724.335 848.135 724.665 848.150 ;
        RECT 723.415 772.655 723.745 772.985 ;
        RECT 723.430 751.225 723.730 772.655 ;
        RECT 723.415 750.895 723.745 751.225 ;
        RECT 723.415 676.095 723.745 676.425 ;
        RECT 723.430 654.650 723.730 676.095 ;
        RECT 723.430 654.350 724.650 654.650 ;
        RECT 724.350 608.425 724.650 654.350 ;
        RECT 724.335 608.095 724.665 608.425 ;
        RECT 723.415 607.415 723.745 607.745 ;
        RECT 723.430 531.415 723.730 607.415 ;
        RECT 723.415 531.085 723.745 531.415 ;
        RECT 723.415 494.535 723.745 494.865 ;
        RECT 723.430 469.025 723.730 494.535 ;
        RECT 723.415 468.695 723.745 469.025 ;
        RECT 724.335 421.095 724.665 421.425 ;
        RECT 724.350 420.050 724.650 421.095 ;
        RECT 723.430 419.750 724.650 420.050 ;
        RECT 723.430 365.650 723.730 419.750 ;
        RECT 723.430 365.350 725.570 365.650 ;
        RECT 725.270 318.745 725.570 365.350 ;
        RECT 725.255 318.415 725.585 318.745 ;
        RECT 723.415 317.735 723.745 318.065 ;
        RECT 723.430 269.785 723.730 317.735 ;
        RECT 723.415 269.455 723.745 269.785 ;
        RECT 725.255 234.775 725.585 235.105 ;
        RECT 725.270 222.185 725.570 234.775 ;
        RECT 725.255 221.855 725.585 222.185 ;
        RECT 723.415 193.295 723.745 193.625 ;
        RECT 723.430 144.665 723.730 193.295 ;
        RECT 723.415 144.335 723.745 144.665 ;
        RECT 723.415 96.735 723.745 97.065 ;
        RECT 723.430 95.705 723.730 96.735 ;
        RECT 723.415 95.375 723.745 95.705 ;
        RECT 723.415 75.970 723.745 75.985 ;
        RECT 723.415 75.670 724.650 75.970 ;
        RECT 723.415 75.655 723.745 75.670 ;
        RECT 724.350 62.385 724.650 75.670 ;
        RECT 724.335 62.055 724.665 62.385 ;
      LAYER met5 ;
        RECT 720.020 1493.500 727.140 1495.100 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1048.410 59.060 1048.730 59.120 ;
        RECT 2829.070 59.060 2829.390 59.120 ;
        RECT 1048.410 58.920 2829.390 59.060 ;
        RECT 1048.410 58.860 1048.730 58.920 ;
        RECT 2829.070 58.860 2829.390 58.920 ;
      LAYER via ;
        RECT 1048.440 58.860 1048.700 59.120 ;
        RECT 2829.100 58.860 2829.360 59.120 ;
      LAYER met2 ;
        RECT 1048.020 1323.690 1048.300 1327.135 ;
        RECT 1048.020 1323.550 1048.640 1323.690 ;
        RECT 1048.020 1323.135 1048.300 1323.550 ;
        RECT 1048.500 59.150 1048.640 1323.550 ;
        RECT 1048.440 58.830 1048.700 59.150 ;
        RECT 2829.100 58.830 2829.360 59.150 ;
        RECT 2829.160 17.410 2829.300 58.830 ;
        RECT 2829.160 17.270 2833.900 17.410 ;
        RECT 2833.760 2.400 2833.900 17.270 ;
        RECT 2833.550 -4.800 2834.110 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1427.060 2375.650 1427.340 2377.880 ;
        RECT 1427.930 2375.650 1428.210 2375.765 ;
        RECT 1427.060 2375.510 1428.210 2375.650 ;
        RECT 1427.060 2373.880 1427.340 2375.510 ;
        RECT 1427.930 2375.395 1428.210 2375.510 ;
        RECT 2849.790 2375.395 2850.070 2375.765 ;
        RECT 2849.860 17.410 2850.000 2375.395 ;
        RECT 2849.860 17.270 2851.380 17.410 ;
        RECT 2851.240 2.400 2851.380 17.270 ;
        RECT 2851.030 -4.800 2851.590 2.400 ;
      LAYER via2 ;
        RECT 1427.930 2375.440 1428.210 2375.720 ;
        RECT 2849.790 2375.440 2850.070 2375.720 ;
      LAYER met3 ;
        RECT 1427.905 2375.730 1428.235 2375.745 ;
        RECT 2849.765 2375.730 2850.095 2375.745 ;
        RECT 1427.905 2375.430 2850.095 2375.730 ;
        RECT 1427.905 2375.415 1428.235 2375.430 ;
        RECT 2849.765 2375.415 2850.095 2375.430 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1772.910 1497.600 1773.230 1497.660 ;
        RECT 2128.490 1497.600 2128.810 1497.660 ;
        RECT 1772.910 1497.460 2128.810 1497.600 ;
        RECT 1772.910 1497.400 1773.230 1497.460 ;
        RECT 2128.490 1497.400 2128.810 1497.460 ;
        RECT 2128.490 17.240 2128.810 17.300 ;
        RECT 2869.090 17.240 2869.410 17.300 ;
        RECT 2128.490 17.100 2869.410 17.240 ;
        RECT 2128.490 17.040 2128.810 17.100 ;
        RECT 2869.090 17.040 2869.410 17.100 ;
      LAYER via ;
        RECT 1772.940 1497.400 1773.200 1497.660 ;
        RECT 2128.520 1497.400 2128.780 1497.660 ;
        RECT 2128.520 17.040 2128.780 17.300 ;
        RECT 2869.120 17.040 2869.380 17.300 ;
      LAYER met2 ;
        RECT 1772.930 1501.595 1773.210 1501.965 ;
        RECT 1773.000 1497.690 1773.140 1501.595 ;
        RECT 1772.940 1497.370 1773.200 1497.690 ;
        RECT 2128.520 1497.370 2128.780 1497.690 ;
        RECT 2128.580 17.330 2128.720 1497.370 ;
        RECT 2128.520 17.010 2128.780 17.330 ;
        RECT 2869.120 17.010 2869.380 17.330 ;
        RECT 2869.180 2.400 2869.320 17.010 ;
        RECT 2868.970 -4.800 2869.530 2.400 ;
      LAYER via2 ;
        RECT 1772.930 1501.640 1773.210 1501.920 ;
      LAYER met3 ;
        RECT 1755.835 1501.930 1759.835 1501.935 ;
        RECT 1772.905 1501.930 1773.235 1501.945 ;
        RECT 1755.835 1501.630 1773.235 1501.930 ;
        RECT 1755.835 1501.335 1759.835 1501.630 ;
        RECT 1772.905 1501.615 1773.235 1501.630 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1221.830 1311.280 1222.150 1311.340 ;
        RECT 1227.810 1311.280 1228.130 1311.340 ;
        RECT 1221.830 1311.140 1228.130 1311.280 ;
        RECT 1221.830 1311.080 1222.150 1311.140 ;
        RECT 1227.810 1311.080 1228.130 1311.140 ;
        RECT 1227.810 65.520 1228.130 65.580 ;
        RECT 2884.270 65.520 2884.590 65.580 ;
        RECT 1227.810 65.380 2884.590 65.520 ;
        RECT 1227.810 65.320 1228.130 65.380 ;
        RECT 2884.270 65.320 2884.590 65.380 ;
        RECT 2884.270 2.960 2884.590 3.020 ;
        RECT 2887.030 2.960 2887.350 3.020 ;
        RECT 2884.270 2.820 2887.350 2.960 ;
        RECT 2884.270 2.760 2884.590 2.820 ;
        RECT 2887.030 2.760 2887.350 2.820 ;
      LAYER via ;
        RECT 1221.860 1311.080 1222.120 1311.340 ;
        RECT 1227.840 1311.080 1228.100 1311.340 ;
        RECT 1227.840 65.320 1228.100 65.580 ;
        RECT 2884.300 65.320 2884.560 65.580 ;
        RECT 2884.300 2.760 2884.560 3.020 ;
        RECT 2887.060 2.760 2887.320 3.020 ;
      LAYER met2 ;
        RECT 1221.900 1323.135 1222.180 1327.135 ;
        RECT 1221.920 1311.370 1222.060 1323.135 ;
        RECT 1221.860 1311.050 1222.120 1311.370 ;
        RECT 1227.840 1311.050 1228.100 1311.370 ;
        RECT 1227.900 65.610 1228.040 1311.050 ;
        RECT 1227.840 65.290 1228.100 65.610 ;
        RECT 2884.300 65.290 2884.560 65.610 ;
        RECT 2884.360 3.050 2884.500 65.290 ;
        RECT 2884.300 2.730 2884.560 3.050 ;
        RECT 2887.060 2.730 2887.320 3.050 ;
        RECT 2887.120 2.400 2887.260 2.730 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1579.250 65.860 1579.570 65.920 ;
        RECT 2904.970 65.860 2905.290 65.920 ;
        RECT 1579.250 65.720 2905.290 65.860 ;
        RECT 1579.250 65.660 1579.570 65.720 ;
        RECT 2904.970 65.660 2905.290 65.720 ;
      LAYER via ;
        RECT 1579.280 65.660 1579.540 65.920 ;
        RECT 2905.000 65.660 2905.260 65.920 ;
      LAYER met2 ;
        RECT 1579.780 1323.690 1580.060 1327.135 ;
        RECT 1579.340 1323.550 1580.060 1323.690 ;
        RECT 1579.340 65.950 1579.480 1323.550 ;
        RECT 1579.780 1323.135 1580.060 1323.550 ;
        RECT 1579.280 65.630 1579.540 65.950 ;
        RECT 2905.000 65.630 2905.260 65.950 ;
        RECT 2905.060 2.400 2905.200 65.630 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 813.810 20.980 814.130 21.040 ;
        RECT 852.910 20.980 853.230 21.040 ;
        RECT 813.810 20.840 853.230 20.980 ;
        RECT 813.810 20.780 814.130 20.840 ;
        RECT 852.910 20.780 853.230 20.840 ;
      LAYER via ;
        RECT 813.840 20.780 814.100 21.040 ;
        RECT 852.940 20.780 853.200 21.040 ;
      LAYER met2 ;
        RECT 810.660 1323.690 810.940 1327.135 ;
        RECT 810.660 1323.550 814.040 1323.690 ;
        RECT 810.660 1323.135 810.940 1323.550 ;
        RECT 813.900 21.070 814.040 1323.550 ;
        RECT 813.840 20.750 814.100 21.070 ;
        RECT 852.940 20.750 853.200 21.070 ;
        RECT 853.000 2.400 853.140 20.750 ;
        RECT 852.790 -4.800 853.350 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 759.145 1325.745 759.315 1327.955 ;
        RECT 806.525 1325.745 806.695 1327.955 ;
      LAYER mcon ;
        RECT 759.145 1327.785 759.315 1327.955 ;
        RECT 806.525 1327.785 806.695 1327.955 ;
      LAYER met1 ;
        RECT 698.350 2390.440 698.670 2390.500 ;
        RECT 1317.510 2390.440 1317.830 2390.500 ;
        RECT 698.350 2390.300 1317.830 2390.440 ;
        RECT 698.350 2390.240 698.670 2390.300 ;
        RECT 1317.510 2390.240 1317.830 2390.300 ;
        RECT 698.350 1327.940 698.670 1328.000 ;
        RECT 759.085 1327.940 759.375 1327.985 ;
        RECT 698.350 1327.800 759.375 1327.940 ;
        RECT 698.350 1327.740 698.670 1327.800 ;
        RECT 759.085 1327.755 759.375 1327.800 ;
        RECT 806.465 1327.940 806.755 1327.985 ;
        RECT 806.465 1327.800 869.700 1327.940 ;
        RECT 806.465 1327.755 806.755 1327.800 ;
        RECT 869.560 1326.640 869.700 1327.800 ;
        RECT 869.470 1326.380 869.790 1326.640 ;
        RECT 759.085 1325.900 759.375 1325.945 ;
        RECT 806.465 1325.900 806.755 1325.945 ;
        RECT 759.085 1325.760 806.755 1325.900 ;
        RECT 759.085 1325.715 759.375 1325.760 ;
        RECT 806.465 1325.715 806.755 1325.760 ;
      LAYER via ;
        RECT 698.380 2390.240 698.640 2390.500 ;
        RECT 1317.540 2390.240 1317.800 2390.500 ;
        RECT 698.380 1327.740 698.640 1328.000 ;
        RECT 869.500 1326.380 869.760 1326.640 ;
      LAYER met2 ;
        RECT 698.380 2390.210 698.640 2390.530 ;
        RECT 1317.540 2390.210 1317.800 2390.530 ;
        RECT 698.440 1393.845 698.580 2390.210 ;
        RECT 1317.600 2377.880 1317.740 2390.210 ;
        RECT 1317.580 2373.880 1317.860 2377.880 ;
        RECT 698.370 1393.475 698.650 1393.845 ;
        RECT 698.370 1392.115 698.650 1392.485 ;
        RECT 698.440 1328.030 698.580 1392.115 ;
        RECT 698.380 1327.710 698.640 1328.030 ;
        RECT 869.500 1326.350 869.760 1326.670 ;
        RECT 869.560 24.210 869.700 1326.350 ;
        RECT 869.560 24.070 871.080 24.210 ;
        RECT 870.940 2.400 871.080 24.070 ;
        RECT 870.730 -4.800 871.290 2.400 ;
      LAYER via2 ;
        RECT 698.370 1393.520 698.650 1393.800 ;
        RECT 698.370 1392.160 698.650 1392.440 ;
      LAYER met3 ;
        RECT 698.345 1393.810 698.675 1393.825 ;
        RECT 698.345 1393.495 698.890 1393.810 ;
        RECT 698.590 1392.465 698.890 1393.495 ;
        RECT 698.345 1392.150 698.890 1392.465 ;
        RECT 698.345 1392.135 698.675 1392.150 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 747.645 2374.305 748.735 2374.475 ;
        RECT 862.645 2374.305 862.815 2375.155 ;
        RECT 884.265 2374.475 884.435 2375.155 ;
        RECT 884.265 2374.305 884.895 2374.475 ;
        RECT 930.725 2374.305 930.895 2377.535 ;
        RECT 1000.185 2374.305 1000.355 2377.535 ;
        RECT 1013.525 2374.305 1014.615 2374.475 ;
        RECT 1062.745 2374.305 1062.915 2377.195 ;
        RECT 1186.485 2374.305 1186.655 2377.195 ;
        RECT 1193.845 2374.305 1194.015 2377.535 ;
        RECT 1241.685 2374.305 1241.855 2377.535 ;
        RECT 1242.145 2374.305 1242.315 2376.855 ;
        RECT 1289.985 2374.305 1290.155 2376.855 ;
        RECT 1317.125 2374.305 1318.215 2374.475 ;
        RECT 1345.185 2374.305 1345.355 2376.855 ;
        RECT 1386.585 2374.305 1386.755 2376.855 ;
        RECT 883.805 1326.425 883.975 1331.355 ;
      LAYER mcon ;
        RECT 930.725 2377.365 930.895 2377.535 ;
        RECT 862.645 2374.985 862.815 2375.155 ;
        RECT 748.565 2374.305 748.735 2374.475 ;
        RECT 884.265 2374.985 884.435 2375.155 ;
        RECT 884.725 2374.305 884.895 2374.475 ;
        RECT 1000.185 2377.365 1000.355 2377.535 ;
        RECT 1193.845 2377.365 1194.015 2377.535 ;
        RECT 1062.745 2377.025 1062.915 2377.195 ;
        RECT 1014.445 2374.305 1014.615 2374.475 ;
        RECT 1186.485 2377.025 1186.655 2377.195 ;
        RECT 1241.685 2377.365 1241.855 2377.535 ;
        RECT 1242.145 2376.685 1242.315 2376.855 ;
        RECT 1289.985 2376.685 1290.155 2376.855 ;
        RECT 1345.185 2376.685 1345.355 2376.855 ;
        RECT 1318.045 2374.305 1318.215 2374.475 ;
        RECT 1386.585 2376.685 1386.755 2376.855 ;
        RECT 883.805 1331.185 883.975 1331.355 ;
      LAYER met1 ;
        RECT 930.665 2377.520 930.955 2377.565 ;
        RECT 1000.125 2377.520 1000.415 2377.565 ;
        RECT 930.665 2377.380 1000.415 2377.520 ;
        RECT 930.665 2377.335 930.955 2377.380 ;
        RECT 1000.125 2377.335 1000.415 2377.380 ;
        RECT 1193.785 2377.520 1194.075 2377.565 ;
        RECT 1241.625 2377.520 1241.915 2377.565 ;
        RECT 1193.785 2377.380 1241.915 2377.520 ;
        RECT 1193.785 2377.335 1194.075 2377.380 ;
        RECT 1241.625 2377.335 1241.915 2377.380 ;
        RECT 1062.685 2377.180 1062.975 2377.225 ;
        RECT 1186.425 2377.180 1186.715 2377.225 ;
        RECT 1062.685 2377.040 1186.715 2377.180 ;
        RECT 1062.685 2376.995 1062.975 2377.040 ;
        RECT 1186.425 2376.995 1186.715 2377.040 ;
        RECT 1242.085 2376.840 1242.375 2376.885 ;
        RECT 1289.925 2376.840 1290.215 2376.885 ;
        RECT 1242.085 2376.700 1290.215 2376.840 ;
        RECT 1242.085 2376.655 1242.375 2376.700 ;
        RECT 1289.925 2376.655 1290.215 2376.700 ;
        RECT 1345.125 2376.840 1345.415 2376.885 ;
        RECT 1386.525 2376.840 1386.815 2376.885 ;
        RECT 1345.125 2376.700 1386.815 2376.840 ;
        RECT 1345.125 2376.655 1345.415 2376.700 ;
        RECT 1386.525 2376.655 1386.815 2376.700 ;
        RECT 862.585 2375.140 862.875 2375.185 ;
        RECT 884.205 2375.140 884.495 2375.185 ;
        RECT 862.585 2375.000 884.495 2375.140 ;
        RECT 862.585 2374.955 862.875 2375.000 ;
        RECT 884.205 2374.955 884.495 2375.000 ;
        RECT 687.310 2374.460 687.630 2374.520 ;
        RECT 747.585 2374.460 747.875 2374.505 ;
        RECT 687.310 2374.320 747.875 2374.460 ;
        RECT 687.310 2374.260 687.630 2374.320 ;
        RECT 747.585 2374.275 747.875 2374.320 ;
        RECT 748.505 2374.275 748.795 2374.505 ;
        RECT 862.585 2374.460 862.875 2374.505 ;
        RECT 820.800 2374.320 862.875 2374.460 ;
        RECT 748.580 2374.120 748.720 2374.275 ;
        RECT 820.800 2374.120 820.940 2374.320 ;
        RECT 862.585 2374.275 862.875 2374.320 ;
        RECT 884.665 2374.275 884.955 2374.505 ;
        RECT 930.665 2374.275 930.955 2374.505 ;
        RECT 1000.125 2374.275 1000.415 2374.505 ;
        RECT 1013.465 2374.275 1013.755 2374.505 ;
        RECT 1014.385 2374.460 1014.675 2374.505 ;
        RECT 1062.685 2374.460 1062.975 2374.505 ;
        RECT 1014.385 2374.320 1062.975 2374.460 ;
        RECT 1014.385 2374.275 1014.675 2374.320 ;
        RECT 1062.685 2374.275 1062.975 2374.320 ;
        RECT 1186.425 2374.275 1186.715 2374.505 ;
        RECT 1193.785 2374.275 1194.075 2374.505 ;
        RECT 1241.625 2374.460 1241.915 2374.505 ;
        RECT 1242.085 2374.460 1242.375 2374.505 ;
        RECT 1241.625 2374.320 1242.375 2374.460 ;
        RECT 1241.625 2374.275 1241.915 2374.320 ;
        RECT 1242.085 2374.275 1242.375 2374.320 ;
        RECT 1289.925 2374.275 1290.215 2374.505 ;
        RECT 1317.065 2374.275 1317.355 2374.505 ;
        RECT 1317.985 2374.275 1318.275 2374.505 ;
        RECT 1345.125 2374.275 1345.415 2374.505 ;
        RECT 1386.525 2374.275 1386.815 2374.505 ;
        RECT 748.580 2373.980 820.940 2374.120 ;
        RECT 884.740 2374.120 884.880 2374.275 ;
        RECT 930.740 2374.120 930.880 2374.275 ;
        RECT 884.740 2373.980 930.880 2374.120 ;
        RECT 1000.200 2374.120 1000.340 2374.275 ;
        RECT 1013.540 2374.120 1013.680 2374.275 ;
        RECT 1000.200 2373.980 1013.680 2374.120 ;
        RECT 1186.500 2374.120 1186.640 2374.275 ;
        RECT 1193.860 2374.120 1194.000 2374.275 ;
        RECT 1186.500 2373.980 1194.000 2374.120 ;
        RECT 1290.000 2374.120 1290.140 2374.275 ;
        RECT 1317.140 2374.120 1317.280 2374.275 ;
        RECT 1290.000 2373.980 1317.280 2374.120 ;
        RECT 1318.060 2374.120 1318.200 2374.275 ;
        RECT 1345.200 2374.120 1345.340 2374.275 ;
        RECT 1318.060 2373.980 1345.340 2374.120 ;
        RECT 1386.600 2374.120 1386.740 2374.275 ;
        RECT 1401.690 2374.260 1402.010 2374.520 ;
        RECT 1401.780 2374.120 1401.920 2374.260 ;
        RECT 1386.600 2373.980 1401.920 2374.120 ;
        RECT 687.310 1331.340 687.630 1331.400 ;
        RECT 883.745 1331.340 884.035 1331.385 ;
        RECT 687.310 1331.200 884.035 1331.340 ;
        RECT 687.310 1331.140 687.630 1331.200 ;
        RECT 883.745 1331.155 884.035 1331.200 ;
        RECT 883.730 1326.580 884.050 1326.640 ;
        RECT 883.535 1326.440 884.050 1326.580 ;
        RECT 883.730 1326.380 884.050 1326.440 ;
        RECT 883.730 20.640 884.050 20.700 ;
        RECT 888.790 20.640 889.110 20.700 ;
        RECT 883.730 20.500 889.110 20.640 ;
        RECT 883.730 20.440 884.050 20.500 ;
        RECT 888.790 20.440 889.110 20.500 ;
      LAYER via ;
        RECT 687.340 2374.260 687.600 2374.520 ;
        RECT 1401.720 2374.260 1401.980 2374.520 ;
        RECT 687.340 1331.140 687.600 1331.400 ;
        RECT 883.760 1326.380 884.020 1326.640 ;
        RECT 883.760 20.440 884.020 20.700 ;
        RECT 888.820 20.440 889.080 20.700 ;
      LAYER met2 ;
        RECT 687.340 2374.230 687.600 2374.550 ;
        RECT 1401.720 2374.290 1401.980 2374.550 ;
        RECT 1404.060 2374.290 1404.340 2377.880 ;
        RECT 1401.720 2374.230 1404.340 2374.290 ;
        RECT 687.400 1393.845 687.540 2374.230 ;
        RECT 1401.780 2374.150 1404.340 2374.230 ;
        RECT 1404.060 2373.880 1404.340 2374.150 ;
        RECT 687.330 1393.475 687.610 1393.845 ;
        RECT 687.330 1392.115 687.610 1392.485 ;
        RECT 687.400 1331.430 687.540 1392.115 ;
        RECT 687.340 1331.110 687.600 1331.430 ;
        RECT 883.760 1326.350 884.020 1326.670 ;
        RECT 883.820 20.730 883.960 1326.350 ;
        RECT 883.760 20.410 884.020 20.730 ;
        RECT 888.820 20.410 889.080 20.730 ;
        RECT 888.880 2.400 889.020 20.410 ;
        RECT 888.670 -4.800 889.230 2.400 ;
      LAYER via2 ;
        RECT 687.330 1393.520 687.610 1393.800 ;
        RECT 687.330 1392.160 687.610 1392.440 ;
      LAYER met3 ;
        RECT 687.305 1393.810 687.635 1393.825 ;
        RECT 687.305 1393.495 687.850 1393.810 ;
        RECT 687.550 1392.465 687.850 1393.495 ;
        RECT 687.305 1392.150 687.850 1392.465 ;
        RECT 687.305 1392.135 687.635 1392.150 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1111.965 1256.045 1112.135 1304.155 ;
        RECT 1111.965 786.505 1112.135 821.015 ;
        RECT 1111.965 689.605 1112.135 724.455 ;
        RECT 1111.965 579.785 1112.135 593.895 ;
        RECT 1111.965 496.485 1112.135 531.335 ;
        RECT 1111.965 386.325 1112.135 400.775 ;
        RECT 1111.965 338.045 1112.135 352.495 ;
      LAYER mcon ;
        RECT 1111.965 1303.985 1112.135 1304.155 ;
        RECT 1111.965 820.845 1112.135 821.015 ;
        RECT 1111.965 724.285 1112.135 724.455 ;
        RECT 1111.965 593.725 1112.135 593.895 ;
        RECT 1111.965 531.165 1112.135 531.335 ;
        RECT 1111.965 400.605 1112.135 400.775 ;
        RECT 1111.965 352.325 1112.135 352.495 ;
      LAYER met1 ;
        RECT 1111.890 1304.140 1112.210 1304.200 ;
        RECT 1111.695 1304.000 1112.210 1304.140 ;
        RECT 1111.890 1303.940 1112.210 1304.000 ;
        RECT 1111.905 1256.200 1112.195 1256.245 ;
        RECT 1112.350 1256.200 1112.670 1256.260 ;
        RECT 1111.905 1256.060 1112.670 1256.200 ;
        RECT 1111.905 1256.015 1112.195 1256.060 ;
        RECT 1112.350 1256.000 1112.670 1256.060 ;
        RECT 1111.430 1221.520 1111.750 1221.580 ;
        RECT 1112.350 1221.520 1112.670 1221.580 ;
        RECT 1111.430 1221.380 1112.670 1221.520 ;
        RECT 1111.430 1221.320 1111.750 1221.380 ;
        RECT 1112.350 1221.320 1112.670 1221.380 ;
        RECT 1111.430 1124.960 1111.750 1125.020 ;
        RECT 1112.350 1124.960 1112.670 1125.020 ;
        RECT 1111.430 1124.820 1112.670 1124.960 ;
        RECT 1111.430 1124.760 1111.750 1124.820 ;
        RECT 1112.350 1124.760 1112.670 1124.820 ;
        RECT 1111.430 1028.400 1111.750 1028.460 ;
        RECT 1112.350 1028.400 1112.670 1028.460 ;
        RECT 1111.430 1028.260 1112.670 1028.400 ;
        RECT 1111.430 1028.200 1111.750 1028.260 ;
        RECT 1112.350 1028.200 1112.670 1028.260 ;
        RECT 1111.430 931.840 1111.750 931.900 ;
        RECT 1112.350 931.840 1112.670 931.900 ;
        RECT 1111.430 931.700 1112.670 931.840 ;
        RECT 1111.430 931.640 1111.750 931.700 ;
        RECT 1112.350 931.640 1112.670 931.700 ;
        RECT 1110.970 869.620 1111.290 869.680 ;
        RECT 1112.350 869.620 1112.670 869.680 ;
        RECT 1110.970 869.480 1112.670 869.620 ;
        RECT 1110.970 869.420 1111.290 869.480 ;
        RECT 1112.350 869.420 1112.670 869.480 ;
        RECT 1111.430 835.280 1111.750 835.340 ;
        RECT 1112.350 835.280 1112.670 835.340 ;
        RECT 1111.430 835.140 1112.670 835.280 ;
        RECT 1111.430 835.080 1111.750 835.140 ;
        RECT 1112.350 835.080 1112.670 835.140 ;
        RECT 1111.890 821.000 1112.210 821.060 ;
        RECT 1111.695 820.860 1112.210 821.000 ;
        RECT 1111.890 820.800 1112.210 820.860 ;
        RECT 1111.890 786.660 1112.210 786.720 ;
        RECT 1111.695 786.520 1112.210 786.660 ;
        RECT 1111.890 786.460 1112.210 786.520 ;
        RECT 1111.430 738.380 1111.750 738.440 ;
        RECT 1112.350 738.380 1112.670 738.440 ;
        RECT 1111.430 738.240 1112.670 738.380 ;
        RECT 1111.430 738.180 1111.750 738.240 ;
        RECT 1112.350 738.180 1112.670 738.240 ;
        RECT 1111.890 724.440 1112.210 724.500 ;
        RECT 1111.695 724.300 1112.210 724.440 ;
        RECT 1111.890 724.240 1112.210 724.300 ;
        RECT 1111.890 689.760 1112.210 689.820 ;
        RECT 1111.695 689.620 1112.210 689.760 ;
        RECT 1111.890 689.560 1112.210 689.620 ;
        RECT 1111.430 641.820 1111.750 641.880 ;
        RECT 1112.350 641.820 1112.670 641.880 ;
        RECT 1111.430 641.680 1112.670 641.820 ;
        RECT 1111.430 641.620 1111.750 641.680 ;
        RECT 1112.350 641.620 1112.670 641.680 ;
        RECT 1111.905 593.880 1112.195 593.925 ;
        RECT 1112.350 593.880 1112.670 593.940 ;
        RECT 1111.905 593.740 1112.670 593.880 ;
        RECT 1111.905 593.695 1112.195 593.740 ;
        RECT 1112.350 593.680 1112.670 593.740 ;
        RECT 1111.890 579.940 1112.210 580.000 ;
        RECT 1111.695 579.800 1112.210 579.940 ;
        RECT 1111.890 579.740 1112.210 579.800 ;
        RECT 1111.890 531.320 1112.210 531.380 ;
        RECT 1111.695 531.180 1112.210 531.320 ;
        RECT 1111.890 531.120 1112.210 531.180 ;
        RECT 1111.890 496.640 1112.210 496.700 ;
        RECT 1111.695 496.500 1112.210 496.640 ;
        RECT 1111.890 496.440 1112.210 496.500 ;
        RECT 1111.430 448.700 1111.750 448.760 ;
        RECT 1112.350 448.700 1112.670 448.760 ;
        RECT 1111.430 448.560 1112.670 448.700 ;
        RECT 1111.430 448.500 1111.750 448.560 ;
        RECT 1112.350 448.500 1112.670 448.560 ;
        RECT 1111.905 400.760 1112.195 400.805 ;
        RECT 1112.350 400.760 1112.670 400.820 ;
        RECT 1111.905 400.620 1112.670 400.760 ;
        RECT 1111.905 400.575 1112.195 400.620 ;
        RECT 1112.350 400.560 1112.670 400.620 ;
        RECT 1111.890 386.480 1112.210 386.540 ;
        RECT 1111.695 386.340 1112.210 386.480 ;
        RECT 1111.890 386.280 1112.210 386.340 ;
        RECT 1111.890 352.480 1112.210 352.540 ;
        RECT 1111.695 352.340 1112.210 352.480 ;
        RECT 1111.890 352.280 1112.210 352.340 ;
        RECT 1111.890 338.200 1112.210 338.260 ;
        RECT 1111.695 338.060 1112.210 338.200 ;
        RECT 1111.890 338.000 1112.210 338.060 ;
        RECT 1111.890 241.640 1112.210 241.700 ;
        RECT 1112.350 241.640 1112.670 241.700 ;
        RECT 1111.890 241.500 1112.670 241.640 ;
        RECT 1111.890 241.440 1112.210 241.500 ;
        RECT 1112.350 241.440 1112.670 241.500 ;
        RECT 906.730 61.100 907.050 61.160 ;
        RECT 1111.430 61.100 1111.750 61.160 ;
        RECT 906.730 60.960 1111.750 61.100 ;
        RECT 906.730 60.900 907.050 60.960 ;
        RECT 1111.430 60.900 1111.750 60.960 ;
      LAYER via ;
        RECT 1111.920 1303.940 1112.180 1304.200 ;
        RECT 1112.380 1256.000 1112.640 1256.260 ;
        RECT 1111.460 1221.320 1111.720 1221.580 ;
        RECT 1112.380 1221.320 1112.640 1221.580 ;
        RECT 1111.460 1124.760 1111.720 1125.020 ;
        RECT 1112.380 1124.760 1112.640 1125.020 ;
        RECT 1111.460 1028.200 1111.720 1028.460 ;
        RECT 1112.380 1028.200 1112.640 1028.460 ;
        RECT 1111.460 931.640 1111.720 931.900 ;
        RECT 1112.380 931.640 1112.640 931.900 ;
        RECT 1111.000 869.420 1111.260 869.680 ;
        RECT 1112.380 869.420 1112.640 869.680 ;
        RECT 1111.460 835.080 1111.720 835.340 ;
        RECT 1112.380 835.080 1112.640 835.340 ;
        RECT 1111.920 820.800 1112.180 821.060 ;
        RECT 1111.920 786.460 1112.180 786.720 ;
        RECT 1111.460 738.180 1111.720 738.440 ;
        RECT 1112.380 738.180 1112.640 738.440 ;
        RECT 1111.920 724.240 1112.180 724.500 ;
        RECT 1111.920 689.560 1112.180 689.820 ;
        RECT 1111.460 641.620 1111.720 641.880 ;
        RECT 1112.380 641.620 1112.640 641.880 ;
        RECT 1112.380 593.680 1112.640 593.940 ;
        RECT 1111.920 579.740 1112.180 580.000 ;
        RECT 1111.920 531.120 1112.180 531.380 ;
        RECT 1111.920 496.440 1112.180 496.700 ;
        RECT 1111.460 448.500 1111.720 448.760 ;
        RECT 1112.380 448.500 1112.640 448.760 ;
        RECT 1112.380 400.560 1112.640 400.820 ;
        RECT 1111.920 386.280 1112.180 386.540 ;
        RECT 1111.920 352.280 1112.180 352.540 ;
        RECT 1111.920 338.000 1112.180 338.260 ;
        RECT 1111.920 241.440 1112.180 241.700 ;
        RECT 1112.380 241.440 1112.640 241.700 ;
        RECT 906.760 60.900 907.020 61.160 ;
        RECT 1111.460 60.900 1111.720 61.160 ;
      LAYER met2 ;
        RECT 1117.020 1323.690 1117.300 1327.135 ;
        RECT 1112.900 1323.550 1117.300 1323.690 ;
        RECT 1112.900 1320.970 1113.040 1323.550 ;
        RECT 1117.020 1323.135 1117.300 1323.550 ;
        RECT 1111.980 1320.830 1113.040 1320.970 ;
        RECT 1111.980 1304.230 1112.120 1320.830 ;
        RECT 1111.920 1303.910 1112.180 1304.230 ;
        RECT 1112.380 1255.970 1112.640 1256.290 ;
        RECT 1112.440 1221.610 1112.580 1255.970 ;
        RECT 1111.460 1221.290 1111.720 1221.610 ;
        RECT 1112.380 1221.290 1112.640 1221.610 ;
        RECT 1111.520 1221.010 1111.660 1221.290 ;
        RECT 1111.520 1220.870 1112.120 1221.010 ;
        RECT 1111.980 1173.410 1112.120 1220.870 ;
        RECT 1111.980 1173.270 1112.580 1173.410 ;
        RECT 1112.440 1125.050 1112.580 1173.270 ;
        RECT 1111.460 1124.730 1111.720 1125.050 ;
        RECT 1112.380 1124.730 1112.640 1125.050 ;
        RECT 1111.520 1124.450 1111.660 1124.730 ;
        RECT 1111.520 1124.310 1112.120 1124.450 ;
        RECT 1111.980 1076.850 1112.120 1124.310 ;
        RECT 1111.980 1076.710 1112.580 1076.850 ;
        RECT 1112.440 1028.490 1112.580 1076.710 ;
        RECT 1111.460 1028.170 1111.720 1028.490 ;
        RECT 1112.380 1028.170 1112.640 1028.490 ;
        RECT 1111.520 1027.890 1111.660 1028.170 ;
        RECT 1111.520 1027.750 1112.120 1027.890 ;
        RECT 1111.980 980.290 1112.120 1027.750 ;
        RECT 1111.980 980.150 1112.580 980.290 ;
        RECT 1112.440 931.930 1112.580 980.150 ;
        RECT 1111.460 931.610 1111.720 931.930 ;
        RECT 1112.380 931.610 1112.640 931.930 ;
        RECT 1111.520 931.330 1111.660 931.610 ;
        RECT 1111.520 931.190 1112.120 931.330 ;
        RECT 1111.980 917.845 1112.120 931.190 ;
        RECT 1110.990 917.475 1111.270 917.845 ;
        RECT 1111.910 917.475 1112.190 917.845 ;
        RECT 1111.060 869.710 1111.200 917.475 ;
        RECT 1111.000 869.390 1111.260 869.710 ;
        RECT 1112.380 869.390 1112.640 869.710 ;
        RECT 1112.440 835.370 1112.580 869.390 ;
        RECT 1111.460 835.050 1111.720 835.370 ;
        RECT 1112.380 835.050 1112.640 835.370 ;
        RECT 1111.520 834.770 1111.660 835.050 ;
        RECT 1111.520 834.630 1112.120 834.770 ;
        RECT 1111.980 821.090 1112.120 834.630 ;
        RECT 1111.920 820.770 1112.180 821.090 ;
        RECT 1111.920 786.430 1112.180 786.750 ;
        RECT 1111.980 772.890 1112.120 786.430 ;
        RECT 1111.980 772.750 1112.580 772.890 ;
        RECT 1112.440 738.470 1112.580 772.750 ;
        RECT 1111.460 738.210 1111.720 738.470 ;
        RECT 1111.460 738.150 1112.120 738.210 ;
        RECT 1112.380 738.150 1112.640 738.470 ;
        RECT 1111.520 738.070 1112.120 738.150 ;
        RECT 1111.980 724.530 1112.120 738.070 ;
        RECT 1111.920 724.210 1112.180 724.530 ;
        RECT 1111.920 689.530 1112.180 689.850 ;
        RECT 1111.980 676.330 1112.120 689.530 ;
        RECT 1111.980 676.190 1112.580 676.330 ;
        RECT 1112.440 641.910 1112.580 676.190 ;
        RECT 1111.460 641.650 1111.720 641.910 ;
        RECT 1112.380 641.650 1112.640 641.910 ;
        RECT 1111.460 641.590 1112.640 641.650 ;
        RECT 1111.520 641.510 1112.580 641.590 ;
        RECT 1112.440 593.970 1112.580 641.510 ;
        RECT 1112.380 593.650 1112.640 593.970 ;
        RECT 1111.920 579.710 1112.180 580.030 ;
        RECT 1111.980 545.770 1112.120 579.710 ;
        RECT 1111.520 545.630 1112.120 545.770 ;
        RECT 1111.520 545.090 1111.660 545.630 ;
        RECT 1111.520 544.950 1112.120 545.090 ;
        RECT 1111.980 531.410 1112.120 544.950 ;
        RECT 1111.920 531.090 1112.180 531.410 ;
        RECT 1111.920 496.410 1112.180 496.730 ;
        RECT 1111.980 483.210 1112.120 496.410 ;
        RECT 1111.980 483.070 1112.580 483.210 ;
        RECT 1112.440 448.790 1112.580 483.070 ;
        RECT 1111.460 448.530 1111.720 448.790 ;
        RECT 1112.380 448.530 1112.640 448.790 ;
        RECT 1111.460 448.470 1112.640 448.530 ;
        RECT 1111.520 448.390 1112.580 448.470 ;
        RECT 1112.440 400.850 1112.580 448.390 ;
        RECT 1112.380 400.530 1112.640 400.850 ;
        RECT 1111.920 386.250 1112.180 386.570 ;
        RECT 1111.980 352.570 1112.120 386.250 ;
        RECT 1111.920 352.250 1112.180 352.570 ;
        RECT 1111.920 337.970 1112.180 338.290 ;
        RECT 1111.980 303.690 1112.120 337.970 ;
        RECT 1111.980 303.550 1112.580 303.690 ;
        RECT 1112.440 241.730 1112.580 303.550 ;
        RECT 1111.920 241.410 1112.180 241.730 ;
        RECT 1112.380 241.410 1112.640 241.730 ;
        RECT 1111.980 207.130 1112.120 241.410 ;
        RECT 1111.980 206.990 1112.580 207.130 ;
        RECT 1112.440 158.850 1112.580 206.990 ;
        RECT 1111.520 158.710 1112.580 158.850 ;
        RECT 1111.520 158.170 1111.660 158.710 ;
        RECT 1111.520 158.030 1112.120 158.170 ;
        RECT 1111.980 62.290 1112.120 158.030 ;
        RECT 1111.520 62.150 1112.120 62.290 ;
        RECT 1111.520 61.190 1111.660 62.150 ;
        RECT 906.760 60.870 907.020 61.190 ;
        RECT 1111.460 60.870 1111.720 61.190 ;
        RECT 906.820 2.400 906.960 60.870 ;
        RECT 906.610 -4.800 907.170 2.400 ;
      LAYER via2 ;
        RECT 1110.990 917.520 1111.270 917.800 ;
        RECT 1111.910 917.520 1112.190 917.800 ;
      LAYER met3 ;
        RECT 1110.965 917.810 1111.295 917.825 ;
        RECT 1111.885 917.810 1112.215 917.825 ;
        RECT 1110.965 917.510 1112.215 917.810 ;
        RECT 1110.965 917.495 1111.295 917.510 ;
        RECT 1111.885 917.495 1112.215 917.510 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 924.210 67.900 924.530 67.960 ;
        RECT 1656.070 67.900 1656.390 67.960 ;
        RECT 924.210 67.760 1656.390 67.900 ;
        RECT 924.210 67.700 924.530 67.760 ;
        RECT 1656.070 67.700 1656.390 67.760 ;
      LAYER via ;
        RECT 924.240 67.700 924.500 67.960 ;
        RECT 1656.100 67.700 1656.360 67.960 ;
      LAYER met2 ;
        RECT 1660.740 1323.690 1661.020 1327.135 ;
        RECT 1656.160 1323.550 1661.020 1323.690 ;
        RECT 1656.160 67.990 1656.300 1323.550 ;
        RECT 1660.740 1323.135 1661.020 1323.550 ;
        RECT 924.240 67.670 924.500 67.990 ;
        RECT 1656.100 67.670 1656.360 67.990 ;
        RECT 924.300 2.400 924.440 67.670 ;
        RECT 924.090 -4.800 924.650 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 759.145 2393.685 759.315 2394.535 ;
        RECT 855.745 2388.925 855.915 2393.855 ;
        RECT 903.585 2388.925 903.755 2393.855 ;
        RECT 952.345 2393.685 952.975 2393.855 ;
        RECT 952.805 2392.325 952.975 2393.685 ;
        RECT 939.005 1326.425 939.175 1331.015 ;
      LAYER mcon ;
        RECT 759.145 2394.365 759.315 2394.535 ;
        RECT 855.745 2393.685 855.915 2393.855 ;
        RECT 903.585 2393.685 903.755 2393.855 ;
        RECT 939.005 1330.845 939.175 1331.015 ;
      LAYER met1 ;
        RECT 759.085 2394.520 759.375 2394.565 ;
        RECT 759.085 2394.380 787.360 2394.520 ;
        RECT 759.085 2394.335 759.375 2394.380 ;
        RECT 697.430 2393.840 697.750 2393.900 ;
        RECT 759.085 2393.840 759.375 2393.885 ;
        RECT 697.430 2393.700 759.375 2393.840 ;
        RECT 787.220 2393.840 787.360 2394.380 ;
        RECT 855.685 2393.840 855.975 2393.885 ;
        RECT 787.220 2393.700 855.975 2393.840 ;
        RECT 697.430 2393.640 697.750 2393.700 ;
        RECT 759.085 2393.655 759.375 2393.700 ;
        RECT 855.685 2393.655 855.975 2393.700 ;
        RECT 903.525 2393.840 903.815 2393.885 ;
        RECT 952.285 2393.840 952.575 2393.885 ;
        RECT 903.525 2393.700 952.575 2393.840 ;
        RECT 903.525 2393.655 903.815 2393.700 ;
        RECT 952.285 2393.655 952.575 2393.700 ;
        RECT 952.745 2392.480 953.035 2392.525 ;
        RECT 1010.230 2392.480 1010.550 2392.540 ;
        RECT 952.745 2392.340 1010.550 2392.480 ;
        RECT 952.745 2392.295 953.035 2392.340 ;
        RECT 1010.230 2392.280 1010.550 2392.340 ;
        RECT 855.685 2389.080 855.975 2389.125 ;
        RECT 903.525 2389.080 903.815 2389.125 ;
        RECT 855.685 2388.940 903.815 2389.080 ;
        RECT 855.685 2388.895 855.975 2388.940 ;
        RECT 903.525 2388.895 903.815 2388.940 ;
        RECT 697.430 1331.000 697.750 1331.060 ;
        RECT 938.945 1331.000 939.235 1331.045 ;
        RECT 697.430 1330.860 939.235 1331.000 ;
        RECT 697.430 1330.800 697.750 1330.860 ;
        RECT 938.945 1330.815 939.235 1330.860 ;
        RECT 938.930 1326.580 939.250 1326.640 ;
        RECT 938.735 1326.440 939.250 1326.580 ;
        RECT 938.930 1326.380 939.250 1326.440 ;
        RECT 938.930 20.640 939.250 20.700 ;
        RECT 942.150 20.640 942.470 20.700 ;
        RECT 938.930 20.500 942.470 20.640 ;
        RECT 938.930 20.440 939.250 20.500 ;
        RECT 942.150 20.440 942.470 20.500 ;
      LAYER via ;
        RECT 697.460 2393.640 697.720 2393.900 ;
        RECT 1010.260 2392.280 1010.520 2392.540 ;
        RECT 697.460 1330.800 697.720 1331.060 ;
        RECT 938.960 1326.380 939.220 1326.640 ;
        RECT 938.960 20.440 939.220 20.700 ;
        RECT 942.180 20.440 942.440 20.700 ;
      LAYER met2 ;
        RECT 697.460 2393.610 697.720 2393.930 ;
        RECT 697.520 1393.845 697.660 2393.610 ;
        RECT 1010.260 2392.250 1010.520 2392.570 ;
        RECT 1010.320 2377.880 1010.460 2392.250 ;
        RECT 1010.300 2373.880 1010.580 2377.880 ;
        RECT 697.450 1393.475 697.730 1393.845 ;
        RECT 697.450 1390.755 697.730 1391.125 ;
        RECT 697.520 1331.090 697.660 1390.755 ;
        RECT 697.460 1330.770 697.720 1331.090 ;
        RECT 938.960 1326.350 939.220 1326.670 ;
        RECT 939.020 20.730 939.160 1326.350 ;
        RECT 938.960 20.410 939.220 20.730 ;
        RECT 942.180 20.410 942.440 20.730 ;
        RECT 942.240 2.400 942.380 20.410 ;
        RECT 942.030 -4.800 942.590 2.400 ;
      LAYER via2 ;
        RECT 697.450 1393.520 697.730 1393.800 ;
        RECT 697.450 1390.800 697.730 1391.080 ;
      LAYER met3 ;
        RECT 697.425 1393.810 697.755 1393.825 ;
        RECT 697.425 1393.495 697.970 1393.810 ;
        RECT 697.670 1391.105 697.970 1393.495 ;
        RECT 697.425 1390.790 697.970 1391.105 ;
        RECT 697.425 1390.775 697.755 1390.790 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 965.610 65.860 965.930 65.920 ;
        RECT 1455.970 65.860 1456.290 65.920 ;
        RECT 965.610 65.720 1456.290 65.860 ;
        RECT 965.610 65.660 965.930 65.720 ;
        RECT 1455.970 65.660 1456.290 65.720 ;
        RECT 960.090 20.640 960.410 20.700 ;
        RECT 965.610 20.640 965.930 20.700 ;
        RECT 960.090 20.500 965.930 20.640 ;
        RECT 960.090 20.440 960.410 20.500 ;
        RECT 965.610 20.440 965.930 20.500 ;
      LAYER via ;
        RECT 965.640 65.660 965.900 65.920 ;
        RECT 1456.000 65.660 1456.260 65.920 ;
        RECT 960.120 20.440 960.380 20.700 ;
        RECT 965.640 20.440 965.900 20.700 ;
      LAYER met2 ;
        RECT 1458.340 1323.690 1458.620 1327.135 ;
        RECT 1456.060 1323.550 1458.620 1323.690 ;
        RECT 1456.060 65.950 1456.200 1323.550 ;
        RECT 1458.340 1323.135 1458.620 1323.550 ;
        RECT 965.640 65.630 965.900 65.950 ;
        RECT 1456.000 65.630 1456.260 65.950 ;
        RECT 965.700 20.730 965.840 65.630 ;
        RECT 960.120 20.410 960.380 20.730 ;
        RECT 965.640 20.410 965.900 20.730 ;
        RECT 960.180 2.400 960.320 20.410 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 979.410 1301.420 979.730 1301.480 ;
        RECT 1770.150 1301.420 1770.470 1301.480 ;
        RECT 979.410 1301.280 1770.470 1301.420 ;
        RECT 979.410 1301.220 979.730 1301.280 ;
        RECT 1770.150 1301.220 1770.470 1301.280 ;
      LAYER via ;
        RECT 979.440 1301.220 979.700 1301.480 ;
        RECT 1770.180 1301.220 1770.440 1301.480 ;
      LAYER met2 ;
        RECT 1770.170 2117.675 1770.450 2118.045 ;
        RECT 1770.240 1301.510 1770.380 2117.675 ;
        RECT 979.440 1301.190 979.700 1301.510 ;
        RECT 1770.180 1301.190 1770.440 1301.510 ;
        RECT 979.500 7.210 979.640 1301.190 ;
        RECT 978.120 7.070 979.640 7.210 ;
        RECT 978.120 2.400 978.260 7.070 ;
        RECT 977.910 -4.800 978.470 2.400 ;
      LAYER via2 ;
        RECT 1770.170 2117.720 1770.450 2118.000 ;
      LAYER met3 ;
        RECT 1755.835 2118.010 1759.835 2118.015 ;
        RECT 1770.145 2118.010 1770.475 2118.025 ;
        RECT 1755.835 2117.710 1770.475 2118.010 ;
        RECT 1755.835 2117.415 1759.835 2117.710 ;
        RECT 1770.145 2117.695 1770.475 2117.710 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 662.010 2376.840 662.330 2376.900 ;
        RECT 1241.610 2376.840 1241.930 2376.900 ;
        RECT 662.010 2376.700 1241.930 2376.840 ;
        RECT 662.010 2376.640 662.330 2376.700 ;
        RECT 1241.610 2376.640 1241.930 2376.700 ;
        RECT 656.950 17.240 657.270 17.300 ;
        RECT 662.010 17.240 662.330 17.300 ;
        RECT 656.950 17.100 662.330 17.240 ;
        RECT 656.950 17.040 657.270 17.100 ;
        RECT 662.010 17.040 662.330 17.100 ;
      LAYER via ;
        RECT 662.040 2376.640 662.300 2376.900 ;
        RECT 1241.640 2376.640 1241.900 2376.900 ;
        RECT 656.980 17.040 657.240 17.300 ;
        RECT 662.040 17.040 662.300 17.300 ;
      LAYER met2 ;
        RECT 1242.140 2377.010 1242.420 2377.880 ;
        RECT 1241.700 2376.930 1242.420 2377.010 ;
        RECT 662.040 2376.610 662.300 2376.930 ;
        RECT 1241.640 2376.870 1242.420 2376.930 ;
        RECT 1241.640 2376.610 1241.900 2376.870 ;
        RECT 662.100 17.330 662.240 2376.610 ;
        RECT 1242.140 2373.880 1242.420 2376.870 ;
        RECT 656.980 17.010 657.240 17.330 ;
        RECT 662.040 17.010 662.300 17.330 ;
        RECT 657.040 2.400 657.180 17.010 ;
        RECT 656.830 -4.800 657.390 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 995.970 20.640 996.290 20.700 ;
        RECT 1000.110 20.640 1000.430 20.700 ;
        RECT 995.970 20.500 1000.430 20.640 ;
        RECT 995.970 20.440 996.290 20.500 ;
        RECT 1000.110 20.440 1000.430 20.500 ;
      LAYER via ;
        RECT 996.000 20.440 996.260 20.700 ;
        RECT 1000.140 20.440 1000.400 20.700 ;
      LAYER met2 ;
        RECT 1000.130 889.595 1000.410 889.965 ;
        RECT 1000.200 20.730 1000.340 889.595 ;
        RECT 996.000 20.410 996.260 20.730 ;
        RECT 1000.140 20.410 1000.400 20.730 ;
        RECT 996.060 2.400 996.200 20.410 ;
        RECT 995.850 -4.800 996.410 2.400 ;
      LAYER via2 ;
        RECT 1000.130 889.640 1000.410 889.920 ;
      LAYER met3 ;
        RECT 1755.835 2220.010 1759.835 2220.015 ;
        RECT 1769.430 2220.010 1769.810 2220.020 ;
        RECT 1755.835 2219.710 1769.810 2220.010 ;
        RECT 1755.835 2219.415 1759.835 2219.710 ;
        RECT 1769.430 2219.700 1769.810 2219.710 ;
        RECT 1000.105 889.930 1000.435 889.945 ;
        RECT 1769.430 889.930 1769.810 889.940 ;
        RECT 1000.105 889.630 1769.810 889.930 ;
        RECT 1000.105 889.615 1000.435 889.630 ;
        RECT 1769.430 889.620 1769.810 889.630 ;
      LAYER via3 ;
        RECT 1769.460 2219.700 1769.780 2220.020 ;
        RECT 1769.460 889.620 1769.780 889.940 ;
      LAYER met4 ;
        RECT 1769.455 2219.695 1769.785 2220.025 ;
        RECT 1769.470 889.945 1769.770 2219.695 ;
        RECT 1769.455 889.615 1769.785 889.945 ;
    END
  END la_data_out[20]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 719.125 1307.385 719.295 1340.195 ;
      LAYER mcon ;
        RECT 719.125 1340.025 719.295 1340.195 ;
      LAYER met1 ;
        RECT 719.050 1340.180 719.370 1340.240 ;
        RECT 718.855 1340.040 719.370 1340.180 ;
        RECT 719.050 1339.980 719.370 1340.040 ;
        RECT 719.050 1307.540 719.370 1307.600 ;
        RECT 718.855 1307.400 719.370 1307.540 ;
        RECT 719.050 1307.340 719.370 1307.400 ;
        RECT 719.050 887.300 719.370 887.360 ;
        RECT 1028.170 887.300 1028.490 887.360 ;
        RECT 719.050 887.160 1028.490 887.300 ;
        RECT 719.050 887.100 719.370 887.160 ;
        RECT 1028.170 887.100 1028.490 887.160 ;
        RECT 1028.170 2.960 1028.490 3.020 ;
        RECT 1031.390 2.960 1031.710 3.020 ;
        RECT 1028.170 2.820 1031.710 2.960 ;
        RECT 1028.170 2.760 1028.490 2.820 ;
        RECT 1031.390 2.760 1031.710 2.820 ;
      LAYER via ;
        RECT 719.080 1339.980 719.340 1340.240 ;
        RECT 719.080 1307.340 719.340 1307.600 ;
        RECT 719.080 887.100 719.340 887.360 ;
        RECT 1028.200 887.100 1028.460 887.360 ;
        RECT 1028.200 2.760 1028.460 3.020 ;
        RECT 1031.420 2.760 1031.680 3.020 ;
      LAYER met2 ;
        RECT 719.070 2023.835 719.350 2024.205 ;
        RECT 719.140 1340.270 719.280 2023.835 ;
        RECT 719.080 1339.950 719.340 1340.270 ;
        RECT 719.080 1307.310 719.340 1307.630 ;
        RECT 719.140 887.390 719.280 1307.310 ;
        RECT 719.080 887.070 719.340 887.390 ;
        RECT 1028.200 887.070 1028.460 887.390 ;
        RECT 1028.260 3.050 1028.400 887.070 ;
        RECT 1028.200 2.730 1028.460 3.050 ;
        RECT 1031.420 2.730 1031.680 3.050 ;
        RECT 1031.480 2.400 1031.620 2.730 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
      LAYER via2 ;
        RECT 719.070 2023.880 719.350 2024.160 ;
      LAYER met3 ;
        RECT 715.810 2027.655 719.810 2028.255 ;
        RECT 717.910 2024.170 718.210 2027.655 ;
        RECT 719.045 2024.170 719.375 2024.185 ;
        RECT 717.910 2023.870 719.375 2024.170 ;
        RECT 719.045 2023.855 719.375 2023.870 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1049.330 47.160 1049.650 47.220 ;
        RECT 1771.990 47.160 1772.310 47.220 ;
        RECT 1049.330 47.020 1772.310 47.160 ;
        RECT 1049.330 46.960 1049.650 47.020 ;
        RECT 1771.990 46.960 1772.310 47.020 ;
      LAYER via ;
        RECT 1049.360 46.960 1049.620 47.220 ;
        RECT 1772.020 46.960 1772.280 47.220 ;
      LAYER met2 ;
        RECT 1772.010 1621.275 1772.290 1621.645 ;
        RECT 1772.080 47.250 1772.220 1621.275 ;
        RECT 1049.360 46.930 1049.620 47.250 ;
        RECT 1772.020 46.930 1772.280 47.250 ;
        RECT 1049.420 2.400 1049.560 46.930 ;
        RECT 1049.210 -4.800 1049.770 2.400 ;
      LAYER via2 ;
        RECT 1772.010 1621.320 1772.290 1621.600 ;
      LAYER met3 ;
        RECT 1755.835 1621.610 1759.835 1621.615 ;
        RECT 1771.985 1621.610 1772.315 1621.625 ;
        RECT 1755.835 1621.310 1772.315 1621.610 ;
        RECT 1755.835 1621.015 1759.835 1621.310 ;
        RECT 1771.985 1621.295 1772.315 1621.310 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 759.145 13.345 759.315 14.195 ;
        RECT 793.645 13.345 793.815 18.275 ;
      LAYER mcon ;
        RECT 793.645 18.105 793.815 18.275 ;
        RECT 759.145 14.025 759.315 14.195 ;
      LAYER met1 ;
        RECT 707.090 1308.900 707.410 1308.960 ;
        RECT 742.050 1308.900 742.370 1308.960 ;
        RECT 707.090 1308.760 742.370 1308.900 ;
        RECT 707.090 1308.700 707.410 1308.760 ;
        RECT 742.050 1308.700 742.370 1308.760 ;
        RECT 793.585 18.260 793.875 18.305 ;
        RECT 1067.270 18.260 1067.590 18.320 ;
        RECT 793.585 18.120 1067.590 18.260 ;
        RECT 793.585 18.075 793.875 18.120 ;
        RECT 1067.270 18.060 1067.590 18.120 ;
        RECT 742.050 14.180 742.370 14.240 ;
        RECT 759.085 14.180 759.375 14.225 ;
        RECT 742.050 14.040 759.375 14.180 ;
        RECT 742.050 13.980 742.370 14.040 ;
        RECT 759.085 13.995 759.375 14.040 ;
        RECT 759.085 13.500 759.375 13.545 ;
        RECT 793.585 13.500 793.875 13.545 ;
        RECT 759.085 13.360 793.875 13.500 ;
        RECT 759.085 13.315 759.375 13.360 ;
        RECT 793.585 13.315 793.875 13.360 ;
      LAYER via ;
        RECT 707.120 1308.700 707.380 1308.960 ;
        RECT 742.080 1308.700 742.340 1308.960 ;
        RECT 1067.300 18.060 1067.560 18.320 ;
        RECT 742.080 13.980 742.340 14.240 ;
      LAYER met2 ;
        RECT 706.190 1822.555 706.470 1822.925 ;
        RECT 706.260 1355.650 706.400 1822.555 ;
        RECT 706.260 1355.510 707.320 1355.650 ;
        RECT 707.180 1308.990 707.320 1355.510 ;
        RECT 707.120 1308.670 707.380 1308.990 ;
        RECT 742.080 1308.670 742.340 1308.990 ;
        RECT 742.140 14.270 742.280 1308.670 ;
        RECT 1067.300 18.030 1067.560 18.350 ;
        RECT 742.080 13.950 742.340 14.270 ;
        RECT 1067.360 2.400 1067.500 18.030 ;
        RECT 1067.150 -4.800 1067.710 2.400 ;
      LAYER via2 ;
        RECT 706.190 1822.600 706.470 1822.880 ;
      LAYER met3 ;
        RECT 706.165 1822.890 706.495 1822.905 ;
        RECT 715.810 1822.890 719.810 1822.895 ;
        RECT 706.165 1822.590 719.810 1822.890 ;
        RECT 706.165 1822.575 706.495 1822.590 ;
        RECT 715.810 1822.295 719.810 1822.590 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1085.210 20.640 1085.530 20.700 ;
        RECT 1089.810 20.640 1090.130 20.700 ;
        RECT 1085.210 20.500 1090.130 20.640 ;
        RECT 1085.210 20.440 1085.530 20.500 ;
        RECT 1089.810 20.440 1090.130 20.500 ;
      LAYER via ;
        RECT 1085.240 20.440 1085.500 20.700 ;
        RECT 1089.840 20.440 1090.100 20.700 ;
      LAYER met2 ;
        RECT 1089.830 885.515 1090.110 885.885 ;
        RECT 1089.900 20.730 1090.040 885.515 ;
        RECT 1085.240 20.410 1085.500 20.730 ;
        RECT 1089.840 20.410 1090.100 20.730 ;
        RECT 1085.300 2.400 1085.440 20.410 ;
        RECT 1085.090 -4.800 1085.650 2.400 ;
      LAYER via2 ;
        RECT 1089.830 885.560 1090.110 885.840 ;
      LAYER met3 ;
        RECT 1755.835 2263.530 1759.835 2263.535 ;
        RECT 1768.510 2263.530 1768.890 2263.540 ;
        RECT 1755.835 2263.230 1768.890 2263.530 ;
        RECT 1755.835 2262.935 1759.835 2263.230 ;
        RECT 1768.510 2263.220 1768.890 2263.230 ;
        RECT 1089.805 885.850 1090.135 885.865 ;
        RECT 1768.510 885.850 1768.890 885.860 ;
        RECT 1089.805 885.550 1768.890 885.850 ;
        RECT 1089.805 885.535 1090.135 885.550 ;
        RECT 1768.510 885.540 1768.890 885.550 ;
      LAYER via3 ;
        RECT 1768.540 2263.220 1768.860 2263.540 ;
        RECT 1768.540 885.540 1768.860 885.860 ;
      LAYER met4 ;
        RECT 1768.535 2263.215 1768.865 2263.545 ;
        RECT 1768.550 885.865 1768.850 2263.215 ;
        RECT 1768.535 885.535 1768.865 885.865 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1102.690 53.960 1103.010 54.020 ;
        RECT 1766.930 53.960 1767.250 54.020 ;
        RECT 1102.690 53.820 1767.250 53.960 ;
        RECT 1102.690 53.760 1103.010 53.820 ;
        RECT 1766.930 53.760 1767.250 53.820 ;
      LAYER via ;
        RECT 1102.720 53.760 1102.980 54.020 ;
        RECT 1766.960 53.760 1767.220 54.020 ;
      LAYER met2 ;
        RECT 1766.950 1920.475 1767.230 1920.845 ;
        RECT 1767.020 54.050 1767.160 1920.475 ;
        RECT 1102.720 53.730 1102.980 54.050 ;
        RECT 1766.960 53.730 1767.220 54.050 ;
        RECT 1102.780 2.400 1102.920 53.730 ;
        RECT 1102.570 -4.800 1103.130 2.400 ;
      LAYER via2 ;
        RECT 1766.950 1920.520 1767.230 1920.800 ;
      LAYER met3 ;
        RECT 1755.835 1920.810 1759.835 1920.815 ;
        RECT 1766.925 1920.810 1767.255 1920.825 ;
        RECT 1755.835 1920.510 1767.255 1920.810 ;
        RECT 1755.835 1920.215 1759.835 1920.510 ;
        RECT 1766.925 1920.495 1767.255 1920.510 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 718.665 1301.605 718.835 1328.975 ;
        RECT 1117.945 1207.425 1118.115 1255.875 ;
        RECT 1117.945 241.485 1118.115 289.595 ;
        RECT 1117.945 144.925 1118.115 193.035 ;
        RECT 1117.945 48.365 1118.115 96.475 ;
      LAYER mcon ;
        RECT 718.665 1328.805 718.835 1328.975 ;
        RECT 1117.945 1255.705 1118.115 1255.875 ;
        RECT 1117.945 289.425 1118.115 289.595 ;
        RECT 1117.945 192.865 1118.115 193.035 ;
        RECT 1117.945 96.305 1118.115 96.475 ;
      LAYER met1 ;
        RECT 718.590 1328.960 718.910 1329.020 ;
        RECT 718.395 1328.820 718.910 1328.960 ;
        RECT 718.590 1328.760 718.910 1328.820 ;
        RECT 718.605 1301.760 718.895 1301.805 ;
        RECT 1117.870 1301.760 1118.190 1301.820 ;
        RECT 718.605 1301.620 1118.190 1301.760 ;
        RECT 718.605 1301.575 718.895 1301.620 ;
        RECT 1117.870 1301.560 1118.190 1301.620 ;
        RECT 1117.870 1255.860 1118.190 1255.920 ;
        RECT 1117.675 1255.720 1118.190 1255.860 ;
        RECT 1117.870 1255.660 1118.190 1255.720 ;
        RECT 1117.870 1207.580 1118.190 1207.640 ;
        RECT 1117.675 1207.440 1118.190 1207.580 ;
        RECT 1117.870 1207.380 1118.190 1207.440 ;
        RECT 1117.870 1111.020 1118.190 1111.080 ;
        RECT 1118.790 1111.020 1119.110 1111.080 ;
        RECT 1117.870 1110.880 1119.110 1111.020 ;
        RECT 1117.870 1110.820 1118.190 1110.880 ;
        RECT 1118.790 1110.820 1119.110 1110.880 ;
        RECT 1117.870 1014.460 1118.190 1014.520 ;
        RECT 1118.790 1014.460 1119.110 1014.520 ;
        RECT 1117.870 1014.320 1119.110 1014.460 ;
        RECT 1117.870 1014.260 1118.190 1014.320 ;
        RECT 1118.790 1014.260 1119.110 1014.320 ;
        RECT 1117.870 917.900 1118.190 917.960 ;
        RECT 1118.790 917.900 1119.110 917.960 ;
        RECT 1117.870 917.760 1119.110 917.900 ;
        RECT 1117.870 917.700 1118.190 917.760 ;
        RECT 1118.790 917.700 1119.110 917.760 ;
        RECT 1117.870 772.720 1118.190 772.780 ;
        RECT 1118.790 772.720 1119.110 772.780 ;
        RECT 1117.870 772.580 1119.110 772.720 ;
        RECT 1117.870 772.520 1118.190 772.580 ;
        RECT 1118.790 772.520 1119.110 772.580 ;
        RECT 1117.870 676.160 1118.190 676.220 ;
        RECT 1118.790 676.160 1119.110 676.220 ;
        RECT 1117.870 676.020 1119.110 676.160 ;
        RECT 1117.870 675.960 1118.190 676.020 ;
        RECT 1118.790 675.960 1119.110 676.020 ;
        RECT 1117.870 579.600 1118.190 579.660 ;
        RECT 1118.790 579.600 1119.110 579.660 ;
        RECT 1117.870 579.460 1119.110 579.600 ;
        RECT 1117.870 579.400 1118.190 579.460 ;
        RECT 1118.790 579.400 1119.110 579.460 ;
        RECT 1117.870 483.040 1118.190 483.100 ;
        RECT 1118.790 483.040 1119.110 483.100 ;
        RECT 1117.870 482.900 1119.110 483.040 ;
        RECT 1117.870 482.840 1118.190 482.900 ;
        RECT 1118.790 482.840 1119.110 482.900 ;
        RECT 1117.870 289.580 1118.190 289.640 ;
        RECT 1117.675 289.440 1118.190 289.580 ;
        RECT 1117.870 289.380 1118.190 289.440 ;
        RECT 1117.870 241.640 1118.190 241.700 ;
        RECT 1117.675 241.500 1118.190 241.640 ;
        RECT 1117.870 241.440 1118.190 241.500 ;
        RECT 1117.870 193.020 1118.190 193.080 ;
        RECT 1117.675 192.880 1118.190 193.020 ;
        RECT 1117.870 192.820 1118.190 192.880 ;
        RECT 1117.870 145.080 1118.190 145.140 ;
        RECT 1117.675 144.940 1118.190 145.080 ;
        RECT 1117.870 144.880 1118.190 144.940 ;
        RECT 1117.870 96.460 1118.190 96.520 ;
        RECT 1117.675 96.320 1118.190 96.460 ;
        RECT 1117.870 96.260 1118.190 96.320 ;
        RECT 1117.870 48.520 1118.190 48.580 ;
        RECT 1117.675 48.380 1118.190 48.520 ;
        RECT 1117.870 48.320 1118.190 48.380 ;
        RECT 1117.410 2.960 1117.730 3.020 ;
        RECT 1120.630 2.960 1120.950 3.020 ;
        RECT 1117.410 2.820 1120.950 2.960 ;
        RECT 1117.410 2.760 1117.730 2.820 ;
        RECT 1120.630 2.760 1120.950 2.820 ;
      LAYER via ;
        RECT 718.620 1328.760 718.880 1329.020 ;
        RECT 1117.900 1301.560 1118.160 1301.820 ;
        RECT 1117.900 1255.660 1118.160 1255.920 ;
        RECT 1117.900 1207.380 1118.160 1207.640 ;
        RECT 1117.900 1110.820 1118.160 1111.080 ;
        RECT 1118.820 1110.820 1119.080 1111.080 ;
        RECT 1117.900 1014.260 1118.160 1014.520 ;
        RECT 1118.820 1014.260 1119.080 1014.520 ;
        RECT 1117.900 917.700 1118.160 917.960 ;
        RECT 1118.820 917.700 1119.080 917.960 ;
        RECT 1117.900 772.520 1118.160 772.780 ;
        RECT 1118.820 772.520 1119.080 772.780 ;
        RECT 1117.900 675.960 1118.160 676.220 ;
        RECT 1118.820 675.960 1119.080 676.220 ;
        RECT 1117.900 579.400 1118.160 579.660 ;
        RECT 1118.820 579.400 1119.080 579.660 ;
        RECT 1117.900 482.840 1118.160 483.100 ;
        RECT 1118.820 482.840 1119.080 483.100 ;
        RECT 1117.900 289.380 1118.160 289.640 ;
        RECT 1117.900 241.440 1118.160 241.700 ;
        RECT 1117.900 192.820 1118.160 193.080 ;
        RECT 1117.900 144.880 1118.160 145.140 ;
        RECT 1117.900 96.260 1118.160 96.520 ;
        RECT 1117.900 48.320 1118.160 48.580 ;
        RECT 1117.440 2.760 1117.700 3.020 ;
        RECT 1120.660 2.760 1120.920 3.020 ;
      LAYER met2 ;
        RECT 718.150 2033.355 718.430 2033.725 ;
        RECT 718.220 1355.650 718.360 2033.355 ;
        RECT 718.220 1355.510 718.820 1355.650 ;
        RECT 718.680 1329.050 718.820 1355.510 ;
        RECT 718.620 1328.730 718.880 1329.050 ;
        RECT 1117.900 1301.530 1118.160 1301.850 ;
        RECT 1117.960 1255.950 1118.100 1301.530 ;
        RECT 1117.900 1255.630 1118.160 1255.950 ;
        RECT 1117.900 1207.350 1118.160 1207.670 ;
        RECT 1117.960 1159.245 1118.100 1207.350 ;
        RECT 1117.890 1158.875 1118.170 1159.245 ;
        RECT 1118.810 1158.875 1119.090 1159.245 ;
        RECT 1118.880 1111.110 1119.020 1158.875 ;
        RECT 1117.900 1110.790 1118.160 1111.110 ;
        RECT 1118.820 1110.790 1119.080 1111.110 ;
        RECT 1117.960 1062.685 1118.100 1110.790 ;
        RECT 1117.890 1062.315 1118.170 1062.685 ;
        RECT 1118.810 1062.315 1119.090 1062.685 ;
        RECT 1118.880 1014.550 1119.020 1062.315 ;
        RECT 1117.900 1014.230 1118.160 1014.550 ;
        RECT 1118.820 1014.230 1119.080 1014.550 ;
        RECT 1117.960 966.125 1118.100 1014.230 ;
        RECT 1117.890 965.755 1118.170 966.125 ;
        RECT 1118.810 965.755 1119.090 966.125 ;
        RECT 1118.880 917.990 1119.020 965.755 ;
        RECT 1117.900 917.670 1118.160 917.990 ;
        RECT 1118.820 917.670 1119.080 917.990 ;
        RECT 1117.960 869.565 1118.100 917.670 ;
        RECT 1117.890 869.195 1118.170 869.565 ;
        RECT 1118.810 869.195 1119.090 869.565 ;
        RECT 1118.880 821.285 1119.020 869.195 ;
        RECT 1117.890 820.915 1118.170 821.285 ;
        RECT 1118.810 820.915 1119.090 821.285 ;
        RECT 1117.960 772.810 1118.100 820.915 ;
        RECT 1117.900 772.490 1118.160 772.810 ;
        RECT 1118.820 772.490 1119.080 772.810 ;
        RECT 1118.880 724.725 1119.020 772.490 ;
        RECT 1117.890 724.355 1118.170 724.725 ;
        RECT 1118.810 724.355 1119.090 724.725 ;
        RECT 1117.960 676.250 1118.100 724.355 ;
        RECT 1117.900 675.930 1118.160 676.250 ;
        RECT 1118.820 675.930 1119.080 676.250 ;
        RECT 1118.880 628.165 1119.020 675.930 ;
        RECT 1117.890 627.795 1118.170 628.165 ;
        RECT 1118.810 627.795 1119.090 628.165 ;
        RECT 1117.960 579.690 1118.100 627.795 ;
        RECT 1117.900 579.370 1118.160 579.690 ;
        RECT 1118.820 579.370 1119.080 579.690 ;
        RECT 1118.880 531.605 1119.020 579.370 ;
        RECT 1117.890 531.235 1118.170 531.605 ;
        RECT 1118.810 531.235 1119.090 531.605 ;
        RECT 1117.960 483.130 1118.100 531.235 ;
        RECT 1117.900 482.810 1118.160 483.130 ;
        RECT 1118.820 482.810 1119.080 483.130 ;
        RECT 1118.880 435.045 1119.020 482.810 ;
        RECT 1117.890 434.675 1118.170 435.045 ;
        RECT 1118.810 434.675 1119.090 435.045 ;
        RECT 1117.960 289.670 1118.100 434.675 ;
        RECT 1117.900 289.350 1118.160 289.670 ;
        RECT 1117.900 241.410 1118.160 241.730 ;
        RECT 1117.960 193.110 1118.100 241.410 ;
        RECT 1117.900 192.790 1118.160 193.110 ;
        RECT 1117.900 144.850 1118.160 145.170 ;
        RECT 1117.960 96.550 1118.100 144.850 ;
        RECT 1117.900 96.230 1118.160 96.550 ;
        RECT 1117.900 48.290 1118.160 48.610 ;
        RECT 1117.960 14.690 1118.100 48.290 ;
        RECT 1117.500 14.550 1118.100 14.690 ;
        RECT 1117.500 3.050 1117.640 14.550 ;
        RECT 1117.440 2.730 1117.700 3.050 ;
        RECT 1120.660 2.730 1120.920 3.050 ;
        RECT 1120.720 2.400 1120.860 2.730 ;
        RECT 1120.510 -4.800 1121.070 2.400 ;
      LAYER via2 ;
        RECT 718.150 2033.400 718.430 2033.680 ;
        RECT 1117.890 1158.920 1118.170 1159.200 ;
        RECT 1118.810 1158.920 1119.090 1159.200 ;
        RECT 1117.890 1062.360 1118.170 1062.640 ;
        RECT 1118.810 1062.360 1119.090 1062.640 ;
        RECT 1117.890 965.800 1118.170 966.080 ;
        RECT 1118.810 965.800 1119.090 966.080 ;
        RECT 1117.890 869.240 1118.170 869.520 ;
        RECT 1118.810 869.240 1119.090 869.520 ;
        RECT 1117.890 820.960 1118.170 821.240 ;
        RECT 1118.810 820.960 1119.090 821.240 ;
        RECT 1117.890 724.400 1118.170 724.680 ;
        RECT 1118.810 724.400 1119.090 724.680 ;
        RECT 1117.890 627.840 1118.170 628.120 ;
        RECT 1118.810 627.840 1119.090 628.120 ;
        RECT 1117.890 531.280 1118.170 531.560 ;
        RECT 1118.810 531.280 1119.090 531.560 ;
        RECT 1117.890 434.720 1118.170 435.000 ;
        RECT 1118.810 434.720 1119.090 435.000 ;
      LAYER met3 ;
        RECT 715.810 2035.815 719.810 2036.415 ;
        RECT 717.910 2033.705 718.210 2035.815 ;
        RECT 717.910 2033.390 718.455 2033.705 ;
        RECT 718.125 2033.375 718.455 2033.390 ;
        RECT 1117.865 1159.210 1118.195 1159.225 ;
        RECT 1118.785 1159.210 1119.115 1159.225 ;
        RECT 1117.865 1158.910 1119.115 1159.210 ;
        RECT 1117.865 1158.895 1118.195 1158.910 ;
        RECT 1118.785 1158.895 1119.115 1158.910 ;
        RECT 1117.865 1062.650 1118.195 1062.665 ;
        RECT 1118.785 1062.650 1119.115 1062.665 ;
        RECT 1117.865 1062.350 1119.115 1062.650 ;
        RECT 1117.865 1062.335 1118.195 1062.350 ;
        RECT 1118.785 1062.335 1119.115 1062.350 ;
        RECT 1117.865 966.090 1118.195 966.105 ;
        RECT 1118.785 966.090 1119.115 966.105 ;
        RECT 1117.865 965.790 1119.115 966.090 ;
        RECT 1117.865 965.775 1118.195 965.790 ;
        RECT 1118.785 965.775 1119.115 965.790 ;
        RECT 1117.865 869.530 1118.195 869.545 ;
        RECT 1118.785 869.530 1119.115 869.545 ;
        RECT 1117.865 869.230 1119.115 869.530 ;
        RECT 1117.865 869.215 1118.195 869.230 ;
        RECT 1118.785 869.215 1119.115 869.230 ;
        RECT 1117.865 821.250 1118.195 821.265 ;
        RECT 1118.785 821.250 1119.115 821.265 ;
        RECT 1117.865 820.950 1119.115 821.250 ;
        RECT 1117.865 820.935 1118.195 820.950 ;
        RECT 1118.785 820.935 1119.115 820.950 ;
        RECT 1117.865 724.690 1118.195 724.705 ;
        RECT 1118.785 724.690 1119.115 724.705 ;
        RECT 1117.865 724.390 1119.115 724.690 ;
        RECT 1117.865 724.375 1118.195 724.390 ;
        RECT 1118.785 724.375 1119.115 724.390 ;
        RECT 1117.865 628.130 1118.195 628.145 ;
        RECT 1118.785 628.130 1119.115 628.145 ;
        RECT 1117.865 627.830 1119.115 628.130 ;
        RECT 1117.865 627.815 1118.195 627.830 ;
        RECT 1118.785 627.815 1119.115 627.830 ;
        RECT 1117.865 531.570 1118.195 531.585 ;
        RECT 1118.785 531.570 1119.115 531.585 ;
        RECT 1117.865 531.270 1119.115 531.570 ;
        RECT 1117.865 531.255 1118.195 531.270 ;
        RECT 1118.785 531.255 1119.115 531.270 ;
        RECT 1117.865 435.010 1118.195 435.025 ;
        RECT 1118.785 435.010 1119.115 435.025 ;
        RECT 1117.865 434.710 1119.115 435.010 ;
        RECT 1117.865 434.695 1118.195 434.710 ;
        RECT 1118.785 434.695 1119.115 434.710 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1145.010 1309.580 1145.330 1309.640 ;
        RECT 1768.770 1309.580 1769.090 1309.640 ;
        RECT 1145.010 1309.440 1769.090 1309.580 ;
        RECT 1145.010 1309.380 1145.330 1309.440 ;
        RECT 1768.770 1309.380 1769.090 1309.440 ;
        RECT 1138.570 16.220 1138.890 16.280 ;
        RECT 1145.010 16.220 1145.330 16.280 ;
        RECT 1138.570 16.080 1145.330 16.220 ;
        RECT 1138.570 16.020 1138.890 16.080 ;
        RECT 1145.010 16.020 1145.330 16.080 ;
      LAYER via ;
        RECT 1145.040 1309.380 1145.300 1309.640 ;
        RECT 1768.800 1309.380 1769.060 1309.640 ;
        RECT 1138.600 16.020 1138.860 16.280 ;
        RECT 1145.040 16.020 1145.300 16.280 ;
      LAYER met2 ;
        RECT 1768.790 1706.955 1769.070 1707.325 ;
        RECT 1768.860 1309.670 1769.000 1706.955 ;
        RECT 1145.040 1309.350 1145.300 1309.670 ;
        RECT 1768.800 1309.350 1769.060 1309.670 ;
        RECT 1145.100 16.310 1145.240 1309.350 ;
        RECT 1138.600 15.990 1138.860 16.310 ;
        RECT 1145.040 15.990 1145.300 16.310 ;
        RECT 1138.660 2.400 1138.800 15.990 ;
        RECT 1138.450 -4.800 1139.010 2.400 ;
      LAYER via2 ;
        RECT 1768.790 1707.000 1769.070 1707.280 ;
      LAYER met3 ;
        RECT 1755.835 1707.290 1759.835 1707.295 ;
        RECT 1768.765 1707.290 1769.095 1707.305 ;
        RECT 1755.835 1706.990 1769.095 1707.290 ;
        RECT 1755.835 1706.695 1759.835 1706.990 ;
        RECT 1768.765 1706.975 1769.095 1706.990 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 891.550 1311.620 891.870 1311.680 ;
        RECT 896.150 1311.620 896.470 1311.680 ;
        RECT 891.550 1311.480 896.470 1311.620 ;
        RECT 891.550 1311.420 891.870 1311.480 ;
        RECT 896.150 1311.420 896.470 1311.480 ;
        RECT 896.150 65.520 896.470 65.580 ;
        RECT 1152.370 65.520 1152.690 65.580 ;
        RECT 896.150 65.380 1152.690 65.520 ;
        RECT 896.150 65.320 896.470 65.380 ;
        RECT 1152.370 65.320 1152.690 65.380 ;
        RECT 1152.370 2.960 1152.690 3.020 ;
        RECT 1156.510 2.960 1156.830 3.020 ;
        RECT 1152.370 2.820 1156.830 2.960 ;
        RECT 1152.370 2.760 1152.690 2.820 ;
        RECT 1156.510 2.760 1156.830 2.820 ;
      LAYER via ;
        RECT 891.580 1311.420 891.840 1311.680 ;
        RECT 896.180 1311.420 896.440 1311.680 ;
        RECT 896.180 65.320 896.440 65.580 ;
        RECT 1152.400 65.320 1152.660 65.580 ;
        RECT 1152.400 2.760 1152.660 3.020 ;
        RECT 1156.540 2.760 1156.800 3.020 ;
      LAYER met2 ;
        RECT 891.620 1323.135 891.900 1327.135 ;
        RECT 891.640 1311.710 891.780 1323.135 ;
        RECT 891.580 1311.390 891.840 1311.710 ;
        RECT 896.180 1311.390 896.440 1311.710 ;
        RECT 896.240 65.610 896.380 1311.390 ;
        RECT 896.180 65.290 896.440 65.610 ;
        RECT 1152.400 65.290 1152.660 65.610 ;
        RECT 1152.460 3.050 1152.600 65.290 ;
        RECT 1152.400 2.730 1152.660 3.050 ;
        RECT 1156.540 2.730 1156.800 3.050 ;
        RECT 1156.600 2.400 1156.740 2.730 ;
        RECT 1156.390 -4.800 1156.950 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 675.810 52.260 676.130 52.320 ;
        RECT 1767.850 52.260 1768.170 52.320 ;
        RECT 675.810 52.120 1768.170 52.260 ;
        RECT 675.810 52.060 676.130 52.120 ;
        RECT 1767.850 52.060 1768.170 52.120 ;
      LAYER via ;
        RECT 675.840 52.060 676.100 52.320 ;
        RECT 1767.880 52.060 1768.140 52.320 ;
      LAYER met2 ;
        RECT 1767.870 1698.795 1768.150 1699.165 ;
        RECT 1767.940 52.350 1768.080 1698.795 ;
        RECT 675.840 52.030 676.100 52.350 ;
        RECT 1767.880 52.030 1768.140 52.350 ;
        RECT 675.900 3.130 676.040 52.030 ;
        RECT 674.520 2.990 676.040 3.130 ;
        RECT 674.520 2.400 674.660 2.990 ;
        RECT 674.310 -4.800 674.870 2.400 ;
      LAYER via2 ;
        RECT 1767.870 1698.840 1768.150 1699.120 ;
      LAYER met3 ;
        RECT 1755.835 1699.130 1759.835 1699.135 ;
        RECT 1767.845 1699.130 1768.175 1699.145 ;
        RECT 1755.835 1698.830 1768.175 1699.130 ;
        RECT 1755.835 1698.535 1759.835 1698.830 ;
        RECT 1767.845 1698.815 1768.175 1698.830 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1173.605 1326.425 1173.775 1329.995 ;
      LAYER mcon ;
        RECT 1173.605 1329.825 1173.775 1329.995 ;
      LAYER met1 ;
        RECT 716.290 1329.980 716.610 1330.040 ;
        RECT 1173.545 1329.980 1173.835 1330.025 ;
        RECT 716.290 1329.840 1173.835 1329.980 ;
        RECT 716.290 1329.780 716.610 1329.840 ;
        RECT 1173.545 1329.795 1173.835 1329.840 ;
        RECT 1173.530 1326.580 1173.850 1326.640 ;
        RECT 1173.335 1326.440 1173.850 1326.580 ;
        RECT 1173.530 1326.380 1173.850 1326.440 ;
      LAYER via ;
        RECT 716.320 1329.780 716.580 1330.040 ;
        RECT 1173.560 1326.380 1173.820 1326.640 ;
      LAYER met2 ;
        RECT 716.310 2042.875 716.590 2043.245 ;
        RECT 716.380 1330.070 716.520 2042.875 ;
        RECT 716.320 1329.750 716.580 1330.070 ;
        RECT 1173.560 1326.350 1173.820 1326.670 ;
        RECT 1173.620 3.130 1173.760 1326.350 ;
        RECT 1173.620 2.990 1174.220 3.130 ;
        RECT 1174.080 2.400 1174.220 2.990 ;
        RECT 1173.870 -4.800 1174.430 2.400 ;
      LAYER via2 ;
        RECT 716.310 2042.920 716.590 2043.200 ;
      LAYER met3 ;
        RECT 715.810 2045.335 719.810 2045.935 ;
        RECT 716.070 2043.225 716.370 2045.335 ;
        RECT 716.070 2042.910 716.615 2043.225 ;
        RECT 716.285 2042.895 716.615 2042.910 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 729.245 1324.045 729.415 1332.375 ;
      LAYER mcon ;
        RECT 729.245 1332.205 729.415 1332.375 ;
      LAYER met1 ;
        RECT 719.050 1332.360 719.370 1332.420 ;
        RECT 729.185 1332.360 729.475 1332.405 ;
        RECT 719.050 1332.220 729.475 1332.360 ;
        RECT 719.050 1332.160 719.370 1332.220 ;
        RECT 729.185 1332.175 729.475 1332.220 ;
        RECT 729.170 1324.200 729.490 1324.260 ;
        RECT 728.975 1324.060 729.490 1324.200 ;
        RECT 729.170 1324.000 729.490 1324.060 ;
      LAYER via ;
        RECT 719.080 1332.160 719.340 1332.420 ;
        RECT 729.200 1324.000 729.460 1324.260 ;
      LAYER met2 ;
        RECT 719.070 1332.275 719.350 1332.645 ;
        RECT 719.080 1332.130 719.340 1332.275 ;
        RECT 729.200 1323.970 729.460 1324.290 ;
        RECT 729.260 1323.805 729.400 1323.970 ;
        RECT 729.190 1323.435 729.470 1323.805 ;
        RECT 1191.950 31.435 1192.230 31.805 ;
        RECT 1192.020 2.400 1192.160 31.435 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
      LAYER via2 ;
        RECT 719.070 1332.320 719.350 1332.600 ;
        RECT 729.190 1323.480 729.470 1323.760 ;
        RECT 1191.950 31.480 1192.230 31.760 ;
      LAYER met3 ;
        RECT 715.810 1335.415 719.810 1336.015 ;
        RECT 718.830 1332.625 719.130 1335.415 ;
        RECT 718.830 1332.310 719.375 1332.625 ;
        RECT 719.045 1332.295 719.375 1332.310 ;
        RECT 729.165 1323.770 729.495 1323.785 ;
        RECT 729.830 1323.770 730.210 1323.780 ;
        RECT 729.165 1323.470 730.210 1323.770 ;
        RECT 729.165 1323.455 729.495 1323.470 ;
        RECT 729.830 1323.460 730.210 1323.470 ;
        RECT 729.830 31.770 730.210 31.780 ;
        RECT 1191.925 31.770 1192.255 31.785 ;
        RECT 729.830 31.470 1192.255 31.770 ;
        RECT 729.830 31.460 730.210 31.470 ;
        RECT 1191.925 31.455 1192.255 31.470 ;
      LAYER via3 ;
        RECT 729.860 1323.460 730.180 1323.780 ;
        RECT 729.860 31.460 730.180 31.780 ;
      LAYER met4 ;
        RECT 729.855 1323.455 730.185 1323.785 ;
        RECT 729.870 31.785 730.170 1323.455 ;
        RECT 729.855 31.455 730.185 31.785 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1211.325 1326.425 1211.495 1333.055 ;
      LAYER mcon ;
        RECT 1211.325 1332.885 1211.495 1333.055 ;
      LAYER met1 ;
        RECT 1754.510 1488.420 1754.830 1488.480 ;
        RECT 1765.090 1488.420 1765.410 1488.480 ;
        RECT 1754.510 1488.280 1765.410 1488.420 ;
        RECT 1754.510 1488.220 1754.830 1488.280 ;
        RECT 1765.090 1488.220 1765.410 1488.280 ;
        RECT 1211.265 1333.040 1211.555 1333.085 ;
        RECT 1752.210 1333.040 1752.530 1333.100 ;
        RECT 1211.265 1332.900 1752.530 1333.040 ;
        RECT 1211.265 1332.855 1211.555 1332.900 ;
        RECT 1752.210 1332.840 1752.530 1332.900 ;
        RECT 1211.250 1326.580 1211.570 1326.640 ;
        RECT 1211.055 1326.440 1211.570 1326.580 ;
        RECT 1211.250 1326.380 1211.570 1326.440 ;
      LAYER via ;
        RECT 1754.540 1488.220 1754.800 1488.480 ;
        RECT 1765.120 1488.220 1765.380 1488.480 ;
        RECT 1752.240 1332.840 1752.500 1333.100 ;
        RECT 1211.280 1326.380 1211.540 1326.640 ;
      LAYER met2 ;
        RECT 1490.490 2379.475 1490.770 2379.845 ;
        RECT 1490.560 2377.880 1490.700 2379.475 ;
        RECT 1490.540 2373.880 1490.820 2377.880 ;
        RECT 1765.110 1498.875 1765.390 1499.245 ;
        RECT 1765.180 1488.510 1765.320 1498.875 ;
        RECT 1754.540 1488.250 1754.800 1488.510 ;
        RECT 1753.220 1488.190 1754.800 1488.250 ;
        RECT 1765.120 1488.190 1765.380 1488.510 ;
        RECT 1753.220 1488.110 1754.740 1488.190 ;
        RECT 1753.220 1487.740 1753.360 1488.110 ;
        RECT 1752.300 1487.600 1753.360 1487.740 ;
        RECT 1752.300 1333.130 1752.440 1487.600 ;
        RECT 1752.240 1332.810 1752.500 1333.130 ;
        RECT 1211.280 1326.525 1211.540 1326.670 ;
        RECT 1211.270 1326.155 1211.550 1326.525 ;
        RECT 1209.890 14.435 1210.170 14.805 ;
        RECT 1209.960 2.400 1210.100 14.435 ;
        RECT 1209.750 -4.800 1210.310 2.400 ;
      LAYER via2 ;
        RECT 1490.490 2379.520 1490.770 2379.800 ;
        RECT 1765.110 1498.920 1765.390 1499.200 ;
        RECT 1211.270 1326.200 1211.550 1326.480 ;
        RECT 1209.890 14.480 1210.170 14.760 ;
      LAYER met3 ;
        RECT 1490.465 2379.810 1490.795 2379.825 ;
        RECT 1764.830 2379.810 1765.210 2379.820 ;
        RECT 1490.465 2379.510 1765.210 2379.810 ;
        RECT 1490.465 2379.495 1490.795 2379.510 ;
        RECT 1764.830 2379.500 1765.210 2379.510 ;
        RECT 1765.085 1499.220 1765.415 1499.225 ;
        RECT 1764.830 1499.210 1765.415 1499.220 ;
        RECT 1764.830 1498.910 1765.640 1499.210 ;
        RECT 1764.830 1498.900 1765.415 1498.910 ;
        RECT 1765.085 1498.895 1765.415 1498.900 ;
        RECT 1210.070 1326.490 1210.450 1326.500 ;
        RECT 1211.245 1326.490 1211.575 1326.505 ;
        RECT 1210.070 1326.190 1211.575 1326.490 ;
        RECT 1210.070 1326.180 1210.450 1326.190 ;
        RECT 1211.245 1326.175 1211.575 1326.190 ;
        RECT 1209.865 14.780 1210.195 14.785 ;
        RECT 1209.865 14.770 1210.450 14.780 ;
        RECT 1209.640 14.470 1210.450 14.770 ;
        RECT 1209.865 14.460 1210.450 14.470 ;
        RECT 1209.865 14.455 1210.195 14.460 ;
      LAYER via3 ;
        RECT 1764.860 2379.500 1765.180 2379.820 ;
        RECT 1764.860 1498.900 1765.180 1499.220 ;
        RECT 1210.100 1326.180 1210.420 1326.500 ;
        RECT 1210.100 14.460 1210.420 14.780 ;
      LAYER met4 ;
        RECT 1764.855 2379.495 1765.185 2379.825 ;
        RECT 1764.870 1499.225 1765.170 2379.495 ;
        RECT 1764.855 1498.895 1765.185 1499.225 ;
        RECT 1210.095 1326.175 1210.425 1326.505 ;
        RECT 1210.110 14.785 1210.410 1326.175 ;
        RECT 1210.095 14.455 1210.425 14.785 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1227.885 2.805 1228.055 14.535 ;
      LAYER mcon ;
        RECT 1227.885 14.365 1228.055 14.535 ;
      LAYER met1 ;
        RECT 1227.350 68.580 1227.670 68.640 ;
        RECT 1725.530 68.580 1725.850 68.640 ;
        RECT 1227.350 68.440 1725.850 68.580 ;
        RECT 1227.350 68.380 1227.670 68.440 ;
        RECT 1725.530 68.380 1725.850 68.440 ;
        RECT 1227.810 14.520 1228.130 14.580 ;
        RECT 1227.615 14.380 1228.130 14.520 ;
        RECT 1227.810 14.320 1228.130 14.380 ;
        RECT 1227.810 2.960 1228.130 3.020 ;
        RECT 1227.615 2.820 1228.130 2.960 ;
        RECT 1227.810 2.760 1228.130 2.820 ;
      LAYER via ;
        RECT 1227.380 68.380 1227.640 68.640 ;
        RECT 1725.560 68.380 1725.820 68.640 ;
        RECT 1227.840 14.320 1228.100 14.580 ;
        RECT 1227.840 2.760 1228.100 3.020 ;
      LAYER met2 ;
        RECT 1730.660 1323.690 1730.940 1327.135 ;
        RECT 1725.620 1323.550 1730.940 1323.690 ;
        RECT 1725.620 68.670 1725.760 1323.550 ;
        RECT 1730.660 1323.135 1730.940 1323.550 ;
        RECT 1227.380 68.350 1227.640 68.670 ;
        RECT 1725.560 68.350 1725.820 68.670 ;
        RECT 1227.440 34.410 1227.580 68.350 ;
        RECT 1227.440 34.270 1228.040 34.410 ;
        RECT 1227.900 14.610 1228.040 34.270 ;
        RECT 1227.840 14.290 1228.100 14.610 ;
        RECT 1227.840 2.730 1228.100 3.050 ;
        RECT 1227.900 2.400 1228.040 2.730 ;
        RECT 1227.690 -4.800 1228.250 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1758.190 1524.460 1758.510 1524.520 ;
        RECT 1759.110 1524.460 1759.430 1524.520 ;
        RECT 1758.190 1524.320 1759.430 1524.460 ;
        RECT 1758.190 1524.260 1758.510 1524.320 ;
        RECT 1759.110 1524.260 1759.430 1524.320 ;
        RECT 1248.510 1301.760 1248.830 1301.820 ;
        RECT 1757.730 1301.760 1758.050 1301.820 ;
        RECT 1248.510 1301.620 1758.050 1301.760 ;
        RECT 1248.510 1301.560 1248.830 1301.620 ;
        RECT 1757.730 1301.560 1758.050 1301.620 ;
        RECT 1245.750 16.560 1246.070 16.620 ;
        RECT 1248.510 16.560 1248.830 16.620 ;
        RECT 1245.750 16.420 1248.830 16.560 ;
        RECT 1245.750 16.360 1246.070 16.420 ;
        RECT 1248.510 16.360 1248.830 16.420 ;
      LAYER via ;
        RECT 1758.220 1524.260 1758.480 1524.520 ;
        RECT 1759.140 1524.260 1759.400 1524.520 ;
        RECT 1248.540 1301.560 1248.800 1301.820 ;
        RECT 1757.760 1301.560 1758.020 1301.820 ;
        RECT 1245.780 16.360 1246.040 16.620 ;
        RECT 1248.540 16.360 1248.800 16.620 ;
      LAYER met2 ;
        RECT 1759.130 1551.915 1759.410 1552.285 ;
        RECT 1759.200 1524.550 1759.340 1551.915 ;
        RECT 1758.220 1524.230 1758.480 1524.550 ;
        RECT 1759.140 1524.230 1759.400 1524.550 ;
        RECT 1758.280 1342.050 1758.420 1524.230 ;
        RECT 1757.820 1341.910 1758.420 1342.050 ;
        RECT 1757.820 1301.850 1757.960 1341.910 ;
        RECT 1248.540 1301.530 1248.800 1301.850 ;
        RECT 1757.760 1301.530 1758.020 1301.850 ;
        RECT 1248.600 16.650 1248.740 1301.530 ;
        RECT 1245.780 16.330 1246.040 16.650 ;
        RECT 1248.540 16.330 1248.800 16.650 ;
        RECT 1245.840 2.400 1245.980 16.330 ;
        RECT 1245.630 -4.800 1246.190 2.400 ;
      LAYER via2 ;
        RECT 1759.130 1551.960 1759.410 1552.240 ;
      LAYER met3 ;
        RECT 1755.835 1553.015 1759.835 1553.615 ;
        RECT 1759.350 1552.265 1759.650 1553.015 ;
        RECT 1759.105 1551.950 1759.650 1552.265 ;
        RECT 1759.105 1551.935 1759.435 1551.950 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1768.310 1421.100 1768.630 1421.160 ;
        RECT 1772.910 1421.100 1773.230 1421.160 ;
        RECT 1768.310 1420.960 1773.230 1421.100 ;
        RECT 1768.310 1420.900 1768.630 1420.960 ;
        RECT 1772.910 1420.900 1773.230 1420.960 ;
        RECT 1263.230 54.300 1263.550 54.360 ;
        RECT 1772.910 54.300 1773.230 54.360 ;
        RECT 1263.230 54.160 1773.230 54.300 ;
        RECT 1263.230 54.100 1263.550 54.160 ;
        RECT 1772.910 54.100 1773.230 54.160 ;
      LAYER via ;
        RECT 1768.340 1420.900 1768.600 1421.160 ;
        RECT 1772.940 1420.900 1773.200 1421.160 ;
        RECT 1263.260 54.100 1263.520 54.360 ;
        RECT 1772.940 54.100 1773.200 54.360 ;
      LAYER met2 ;
        RECT 1768.330 1433.595 1768.610 1433.965 ;
        RECT 1768.400 1421.190 1768.540 1433.595 ;
        RECT 1768.340 1420.870 1768.600 1421.190 ;
        RECT 1772.940 1420.870 1773.200 1421.190 ;
        RECT 1773.000 54.390 1773.140 1420.870 ;
        RECT 1263.260 54.070 1263.520 54.390 ;
        RECT 1772.940 54.070 1773.200 54.390 ;
        RECT 1263.320 2.400 1263.460 54.070 ;
        RECT 1263.110 -4.800 1263.670 2.400 ;
      LAYER via2 ;
        RECT 1768.330 1433.640 1768.610 1433.920 ;
      LAYER met3 ;
        RECT 1755.835 1433.930 1759.835 1433.935 ;
        RECT 1768.305 1433.930 1768.635 1433.945 ;
        RECT 1755.835 1433.630 1768.635 1433.930 ;
        RECT 1755.835 1433.335 1759.835 1433.630 ;
        RECT 1768.305 1433.615 1768.635 1433.630 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1241.610 45.800 1241.930 45.860 ;
        RECT 1281.170 45.800 1281.490 45.860 ;
        RECT 1241.610 45.660 1281.490 45.800 ;
        RECT 1241.610 45.600 1241.930 45.660 ;
        RECT 1281.170 45.600 1281.490 45.660 ;
      LAYER via ;
        RECT 1241.640 45.600 1241.900 45.860 ;
        RECT 1281.200 45.600 1281.460 45.860 ;
      LAYER met2 ;
        RECT 1238.460 1323.690 1238.740 1327.135 ;
        RECT 1238.460 1323.550 1241.840 1323.690 ;
        RECT 1238.460 1323.135 1238.740 1323.550 ;
        RECT 1241.700 45.890 1241.840 1323.550 ;
        RECT 1241.640 45.570 1241.900 45.890 ;
        RECT 1281.200 45.570 1281.460 45.890 ;
        RECT 1281.260 2.400 1281.400 45.570 ;
        RECT 1281.050 -4.800 1281.610 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1756.885 1341.385 1757.055 1372.495 ;
      LAYER mcon ;
        RECT 1756.885 1372.325 1757.055 1372.495 ;
      LAYER met1 ;
        RECT 1756.810 1372.480 1757.130 1372.540 ;
        RECT 1756.810 1372.340 1757.325 1372.480 ;
        RECT 1756.810 1372.280 1757.130 1372.340 ;
        RECT 1756.825 1341.540 1757.115 1341.585 ;
        RECT 1758.190 1341.540 1758.510 1341.600 ;
        RECT 1756.825 1341.400 1758.510 1341.540 ;
        RECT 1756.825 1341.355 1757.115 1341.400 ;
        RECT 1758.190 1341.340 1758.510 1341.400 ;
        RECT 1303.710 1310.940 1304.030 1311.000 ;
        RECT 1758.190 1310.940 1758.510 1311.000 ;
        RECT 1303.710 1310.800 1758.510 1310.940 ;
        RECT 1303.710 1310.740 1304.030 1310.800 ;
        RECT 1758.190 1310.740 1758.510 1310.800 ;
        RECT 1303.710 554.240 1304.030 554.500 ;
        RECT 1303.800 553.820 1303.940 554.240 ;
        RECT 1303.710 553.560 1304.030 553.820 ;
        RECT 1299.110 20.640 1299.430 20.700 ;
        RECT 1303.710 20.640 1304.030 20.700 ;
        RECT 1299.110 20.500 1304.030 20.640 ;
        RECT 1299.110 20.440 1299.430 20.500 ;
        RECT 1303.710 20.440 1304.030 20.500 ;
      LAYER via ;
        RECT 1756.840 1372.280 1757.100 1372.540 ;
        RECT 1758.220 1341.340 1758.480 1341.600 ;
        RECT 1303.740 1310.740 1304.000 1311.000 ;
        RECT 1758.220 1310.740 1758.480 1311.000 ;
        RECT 1303.740 554.240 1304.000 554.500 ;
        RECT 1303.740 553.560 1304.000 553.820 ;
        RECT 1299.140 20.440 1299.400 20.700 ;
        RECT 1303.740 20.440 1304.000 20.700 ;
      LAYER met2 ;
        RECT 1756.830 2056.475 1757.110 2056.845 ;
        RECT 1756.900 1372.570 1757.040 2056.475 ;
        RECT 1756.840 1372.250 1757.100 1372.570 ;
        RECT 1758.220 1341.310 1758.480 1341.630 ;
        RECT 1758.280 1311.030 1758.420 1341.310 ;
        RECT 1303.740 1310.710 1304.000 1311.030 ;
        RECT 1758.220 1310.710 1758.480 1311.030 ;
        RECT 1303.800 554.530 1303.940 1310.710 ;
        RECT 1303.740 554.210 1304.000 554.530 ;
        RECT 1303.740 553.530 1304.000 553.850 ;
        RECT 1303.800 20.730 1303.940 553.530 ;
        RECT 1299.140 20.410 1299.400 20.730 ;
        RECT 1303.740 20.410 1304.000 20.730 ;
        RECT 1299.200 2.400 1299.340 20.410 ;
        RECT 1298.990 -4.800 1299.550 2.400 ;
      LAYER via2 ;
        RECT 1756.830 2056.520 1757.110 2056.800 ;
      LAYER met3 ;
        RECT 1755.835 2057.575 1759.835 2058.175 ;
        RECT 1756.590 2056.825 1756.890 2057.575 ;
        RECT 1756.590 2056.510 1757.135 2056.825 ;
        RECT 1756.805 2056.495 1757.135 2056.510 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 696.125 1368.925 696.295 1393.575 ;
        RECT 735.225 18.105 735.395 19.295 ;
      LAYER mcon ;
        RECT 696.125 1393.405 696.295 1393.575 ;
        RECT 735.225 19.125 735.395 19.295 ;
      LAYER met1 ;
        RECT 696.050 2377.520 696.370 2377.580 ;
        RECT 852.910 2377.520 853.230 2377.580 ;
        RECT 696.050 2377.380 853.230 2377.520 ;
        RECT 696.050 2377.320 696.370 2377.380 ;
        RECT 852.910 2377.320 853.230 2377.380 ;
        RECT 696.050 1393.560 696.370 1393.620 ;
        RECT 696.050 1393.420 696.565 1393.560 ;
        RECT 696.050 1393.360 696.370 1393.420 ;
        RECT 696.050 1369.080 696.370 1369.140 ;
        RECT 695.855 1368.940 696.370 1369.080 ;
        RECT 696.050 1368.880 696.370 1368.940 ;
        RECT 735.165 19.280 735.455 19.325 ;
        RECT 735.165 19.140 1293.360 19.280 ;
        RECT 735.165 19.095 735.455 19.140 ;
        RECT 1293.220 18.940 1293.360 19.140 ;
        RECT 1317.050 18.940 1317.370 19.000 ;
        RECT 1293.220 18.800 1317.370 18.940 ;
        RECT 1317.050 18.740 1317.370 18.800 ;
        RECT 696.050 18.260 696.370 18.320 ;
        RECT 735.165 18.260 735.455 18.305 ;
        RECT 696.050 18.120 735.455 18.260 ;
        RECT 696.050 18.060 696.370 18.120 ;
        RECT 735.165 18.075 735.455 18.120 ;
      LAYER via ;
        RECT 696.080 2377.320 696.340 2377.580 ;
        RECT 852.940 2377.320 853.200 2377.580 ;
        RECT 696.080 1393.360 696.340 1393.620 ;
        RECT 696.080 1368.880 696.340 1369.140 ;
        RECT 1317.080 18.740 1317.340 19.000 ;
        RECT 696.080 18.060 696.340 18.320 ;
      LAYER met2 ;
        RECT 854.820 2377.690 855.100 2377.880 ;
        RECT 853.000 2377.610 855.100 2377.690 ;
        RECT 696.080 2377.290 696.340 2377.610 ;
        RECT 852.940 2377.550 855.100 2377.610 ;
        RECT 852.940 2377.290 853.200 2377.550 ;
        RECT 696.140 1393.650 696.280 2377.290 ;
        RECT 854.820 2373.880 855.100 2377.550 ;
        RECT 696.080 1393.330 696.340 1393.650 ;
        RECT 696.080 1368.850 696.340 1369.170 ;
        RECT 696.140 18.350 696.280 1368.850 ;
        RECT 1317.080 18.710 1317.340 19.030 ;
        RECT 696.080 18.030 696.340 18.350 ;
        RECT 1317.140 2.400 1317.280 18.710 ;
        RECT 1316.930 -4.800 1317.490 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 731.490 2374.290 731.770 2374.405 ;
        RECT 733.380 2374.290 733.660 2377.880 ;
        RECT 731.490 2374.150 733.660 2374.290 ;
        RECT 731.490 2374.035 731.770 2374.150 ;
        RECT 733.380 2373.880 733.660 2374.150 ;
        RECT 695.150 2373.355 695.430 2373.725 ;
        RECT 695.220 15.485 695.360 2373.355 ;
        RECT 695.150 15.115 695.430 15.485 ;
        RECT 1335.010 15.115 1335.290 15.485 ;
        RECT 1335.080 2.400 1335.220 15.115 ;
        RECT 1334.870 -4.800 1335.430 2.400 ;
      LAYER via2 ;
        RECT 731.490 2374.080 731.770 2374.360 ;
        RECT 695.150 2373.400 695.430 2373.680 ;
        RECT 695.150 15.160 695.430 15.440 ;
        RECT 1335.010 15.160 1335.290 15.440 ;
      LAYER met3 ;
        RECT 731.465 2374.370 731.795 2374.385 ;
        RECT 718.830 2374.070 731.795 2374.370 ;
        RECT 695.125 2373.690 695.455 2373.705 ;
        RECT 718.830 2373.690 719.130 2374.070 ;
        RECT 731.465 2374.055 731.795 2374.070 ;
        RECT 695.125 2373.390 719.130 2373.690 ;
        RECT 695.125 2373.375 695.455 2373.390 ;
        RECT 695.125 15.450 695.455 15.465 ;
        RECT 1334.985 15.450 1335.315 15.465 ;
        RECT 695.125 15.150 1335.315 15.450 ;
        RECT 695.125 15.135 695.455 15.150 ;
        RECT 1334.985 15.135 1335.315 15.150 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 692.370 60.420 692.690 60.480 ;
        RECT 1125.230 60.420 1125.550 60.480 ;
        RECT 692.370 60.280 1125.550 60.420 ;
        RECT 692.370 60.220 692.690 60.280 ;
        RECT 1125.230 60.220 1125.550 60.280 ;
      LAYER via ;
        RECT 692.400 60.220 692.660 60.480 ;
        RECT 1125.260 60.220 1125.520 60.480 ;
      LAYER met2 ;
        RECT 1128.980 1323.690 1129.260 1327.135 ;
        RECT 1125.320 1323.550 1129.260 1323.690 ;
        RECT 1125.320 60.510 1125.460 1323.550 ;
        RECT 1128.980 1323.135 1129.260 1323.550 ;
        RECT 692.400 60.190 692.660 60.510 ;
        RECT 1125.260 60.190 1125.520 60.510 ;
        RECT 692.460 2.400 692.600 60.190 ;
        RECT 692.250 -4.800 692.810 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1358.985 1326.425 1359.155 1330.335 ;
      LAYER mcon ;
        RECT 1358.985 1330.165 1359.155 1330.335 ;
      LAYER met1 ;
        RECT 1358.925 1330.320 1359.215 1330.365 ;
        RECT 1752.210 1330.320 1752.530 1330.380 ;
        RECT 1358.925 1330.180 1752.530 1330.320 ;
        RECT 1358.925 1330.135 1359.215 1330.180 ;
        RECT 1752.210 1330.120 1752.530 1330.180 ;
        RECT 1358.910 1326.580 1359.230 1326.640 ;
        RECT 1358.715 1326.440 1359.230 1326.580 ;
        RECT 1358.910 1326.380 1359.230 1326.440 ;
        RECT 1352.470 20.640 1352.790 20.700 ;
        RECT 1358.910 20.640 1359.230 20.700 ;
        RECT 1352.470 20.500 1359.230 20.640 ;
        RECT 1352.470 20.440 1352.790 20.500 ;
        RECT 1358.910 20.440 1359.230 20.500 ;
      LAYER via ;
        RECT 1752.240 1330.120 1752.500 1330.380 ;
        RECT 1358.940 1326.380 1359.200 1326.640 ;
        RECT 1352.500 20.440 1352.760 20.700 ;
        RECT 1358.940 20.440 1359.200 20.700 ;
      LAYER met2 ;
        RECT 1525.450 2384.235 1525.730 2384.605 ;
        RECT 1525.520 2377.880 1525.660 2384.235 ;
        RECT 1525.500 2373.880 1525.780 2377.880 ;
        RECT 1751.770 2372.930 1752.050 2373.045 ;
        RECT 1751.380 2372.790 1752.050 2372.930 ;
        RECT 1751.380 1330.490 1751.520 2372.790 ;
        RECT 1751.770 2372.675 1752.050 2372.790 ;
        RECT 1751.380 1330.410 1752.440 1330.490 ;
        RECT 1751.380 1330.350 1752.500 1330.410 ;
        RECT 1752.240 1330.090 1752.500 1330.350 ;
        RECT 1358.940 1326.350 1359.200 1326.670 ;
        RECT 1359.000 20.730 1359.140 1326.350 ;
        RECT 1352.500 20.410 1352.760 20.730 ;
        RECT 1358.940 20.410 1359.200 20.730 ;
        RECT 1352.560 2.400 1352.700 20.410 ;
        RECT 1352.350 -4.800 1352.910 2.400 ;
      LAYER via2 ;
        RECT 1525.450 2384.280 1525.730 2384.560 ;
        RECT 1751.770 2372.720 1752.050 2373.000 ;
      LAYER met3 ;
        RECT 1525.425 2384.580 1525.755 2384.585 ;
        RECT 1525.425 2384.570 1526.010 2384.580 ;
        RECT 1525.425 2384.270 1526.210 2384.570 ;
        RECT 1525.425 2384.260 1526.010 2384.270 ;
        RECT 1525.425 2384.255 1525.755 2384.260 ;
        RECT 1525.630 2373.010 1526.010 2373.020 ;
        RECT 1751.745 2373.010 1752.075 2373.025 ;
        RECT 1525.630 2372.710 1752.075 2373.010 ;
        RECT 1525.630 2372.700 1526.010 2372.710 ;
        RECT 1751.745 2372.695 1752.075 2372.710 ;
      LAYER via3 ;
        RECT 1525.660 2384.260 1525.980 2384.580 ;
        RECT 1525.660 2372.700 1525.980 2373.020 ;
      LAYER met4 ;
        RECT 1525.655 2384.255 1525.985 2384.585 ;
        RECT 1525.670 2373.025 1525.970 2384.255 ;
        RECT 1525.655 2372.695 1525.985 2373.025 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1461.970 2379.475 1462.250 2379.845 ;
        RECT 1462.040 2377.880 1462.180 2379.475 ;
        RECT 1462.020 2373.880 1462.300 2377.880 ;
        RECT 1769.250 2371.995 1769.530 2372.365 ;
        RECT 1769.320 1353.045 1769.460 2371.995 ;
        RECT 1769.250 1352.675 1769.530 1353.045 ;
        RECT 1370.430 15.115 1370.710 15.485 ;
        RECT 1370.500 2.400 1370.640 15.115 ;
        RECT 1370.290 -4.800 1370.850 2.400 ;
      LAYER via2 ;
        RECT 1461.970 2379.520 1462.250 2379.800 ;
        RECT 1769.250 2372.040 1769.530 2372.320 ;
        RECT 1769.250 1352.720 1769.530 1353.000 ;
        RECT 1370.430 15.160 1370.710 15.440 ;
      LAYER met3 ;
        RECT 1461.945 2379.820 1462.275 2379.825 ;
        RECT 1461.945 2379.810 1462.530 2379.820 ;
        RECT 1461.945 2379.510 1462.730 2379.810 ;
        RECT 1461.945 2379.500 1462.530 2379.510 ;
        RECT 1461.945 2379.495 1462.275 2379.500 ;
        RECT 1462.150 2372.330 1462.530 2372.340 ;
        RECT 1769.225 2372.330 1769.555 2372.345 ;
        RECT 1462.150 2372.030 1769.555 2372.330 ;
        RECT 1462.150 2372.020 1462.530 2372.030 ;
        RECT 1769.225 2372.015 1769.555 2372.030 ;
        RECT 1764.830 1353.010 1765.210 1353.020 ;
        RECT 1769.225 1353.010 1769.555 1353.025 ;
        RECT 1764.830 1352.710 1769.555 1353.010 ;
        RECT 1764.830 1352.700 1765.210 1352.710 ;
        RECT 1769.225 1352.695 1769.555 1352.710 ;
        RECT 1370.405 15.450 1370.735 15.465 ;
        RECT 1371.990 15.450 1372.370 15.460 ;
        RECT 1370.405 15.150 1372.370 15.450 ;
        RECT 1370.405 15.135 1370.735 15.150 ;
        RECT 1371.990 15.140 1372.370 15.150 ;
      LAYER via3 ;
        RECT 1462.180 2379.500 1462.500 2379.820 ;
        RECT 1462.180 2372.020 1462.500 2372.340 ;
        RECT 1764.860 1352.700 1765.180 1353.020 ;
        RECT 1372.020 15.140 1372.340 15.460 ;
      LAYER met4 ;
        RECT 1462.175 2379.495 1462.505 2379.825 ;
        RECT 1462.190 2372.345 1462.490 2379.495 ;
        RECT 1462.175 2372.015 1462.505 2372.345 ;
        RECT 1764.855 1352.695 1765.185 1353.025 ;
        RECT 1764.870 1348.690 1765.170 1352.695 ;
        RECT 1764.430 1347.510 1765.610 1348.690 ;
        RECT 1371.590 1330.510 1372.770 1331.690 ;
        RECT 1372.030 15.465 1372.330 1330.510 ;
        RECT 1372.015 15.135 1372.345 15.465 ;
      LAYER met5 ;
        RECT 1764.220 1335.300 1765.820 1348.900 ;
        RECT 1371.380 1333.700 1459.460 1335.300 ;
        RECT 1371.380 1330.300 1372.980 1333.700 ;
        RECT 1457.860 1328.500 1459.460 1333.700 ;
        RECT 1465.220 1333.700 1765.820 1335.300 ;
        RECT 1465.220 1328.500 1466.820 1333.700 ;
        RECT 1457.860 1326.900 1466.820 1328.500 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1393.485 1326.425 1393.655 1330.675 ;
      LAYER mcon ;
        RECT 1393.485 1330.505 1393.655 1330.675 ;
      LAYER met1 ;
        RECT 1767.850 1925.320 1768.170 1925.380 ;
        RECT 1779.350 1925.320 1779.670 1925.380 ;
        RECT 1767.850 1925.180 1779.670 1925.320 ;
        RECT 1767.850 1925.120 1768.170 1925.180 ;
        RECT 1779.350 1925.120 1779.670 1925.180 ;
        RECT 1393.425 1330.660 1393.715 1330.705 ;
        RECT 1779.350 1330.660 1779.670 1330.720 ;
        RECT 1393.425 1330.520 1779.670 1330.660 ;
        RECT 1393.425 1330.475 1393.715 1330.520 ;
        RECT 1779.350 1330.460 1779.670 1330.520 ;
        RECT 1393.410 1326.580 1393.730 1326.640 ;
        RECT 1393.215 1326.440 1393.730 1326.580 ;
        RECT 1393.410 1326.380 1393.730 1326.440 ;
        RECT 1388.350 16.560 1388.670 16.620 ;
        RECT 1393.410 16.560 1393.730 16.620 ;
        RECT 1388.350 16.420 1393.730 16.560 ;
        RECT 1388.350 16.360 1388.670 16.420 ;
        RECT 1393.410 16.360 1393.730 16.420 ;
      LAYER via ;
        RECT 1767.880 1925.120 1768.140 1925.380 ;
        RECT 1779.380 1925.120 1779.640 1925.380 ;
        RECT 1779.380 1330.460 1779.640 1330.720 ;
        RECT 1393.440 1326.380 1393.700 1326.640 ;
        RECT 1388.380 16.360 1388.640 16.620 ;
        RECT 1393.440 16.360 1393.700 16.620 ;
      LAYER met2 ;
        RECT 1767.870 1929.995 1768.150 1930.365 ;
        RECT 1767.940 1925.410 1768.080 1929.995 ;
        RECT 1767.880 1925.090 1768.140 1925.410 ;
        RECT 1779.380 1925.090 1779.640 1925.410 ;
        RECT 1779.440 1330.750 1779.580 1925.090 ;
        RECT 1779.380 1330.430 1779.640 1330.750 ;
        RECT 1393.440 1326.350 1393.700 1326.670 ;
        RECT 1393.500 16.650 1393.640 1326.350 ;
        RECT 1388.380 16.330 1388.640 16.650 ;
        RECT 1393.440 16.330 1393.700 16.650 ;
        RECT 1388.440 2.400 1388.580 16.330 ;
        RECT 1388.230 -4.800 1388.790 2.400 ;
      LAYER via2 ;
        RECT 1767.870 1930.040 1768.150 1930.320 ;
      LAYER met3 ;
        RECT 1755.835 1930.330 1759.835 1930.335 ;
        RECT 1767.845 1930.330 1768.175 1930.345 ;
        RECT 1755.835 1930.030 1768.175 1930.330 ;
        RECT 1755.835 1929.735 1759.835 1930.030 ;
        RECT 1767.845 1930.015 1768.175 1930.030 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1403.605 1326.425 1403.775 1332.715 ;
        RECT 1749.525 1325.745 1749.695 1332.715 ;
      LAYER mcon ;
        RECT 1403.605 1332.545 1403.775 1332.715 ;
        RECT 1749.525 1332.545 1749.695 1332.715 ;
      LAYER met1 ;
        RECT 1403.545 1332.700 1403.835 1332.745 ;
        RECT 1749.465 1332.700 1749.755 1332.745 ;
        RECT 1403.545 1332.560 1749.755 1332.700 ;
        RECT 1403.545 1332.515 1403.835 1332.560 ;
        RECT 1749.465 1332.515 1749.755 1332.560 ;
        RECT 1403.530 1326.580 1403.850 1326.640 ;
        RECT 1403.335 1326.440 1403.850 1326.580 ;
        RECT 1403.530 1326.380 1403.850 1326.440 ;
        RECT 1749.450 1325.900 1749.770 1325.960 ;
        RECT 1749.255 1325.760 1749.770 1325.900 ;
        RECT 1749.450 1325.700 1749.770 1325.760 ;
      LAYER via ;
        RECT 1403.560 1326.380 1403.820 1326.640 ;
        RECT 1749.480 1325.700 1749.740 1325.960 ;
      LAYER met2 ;
        RECT 1091.210 2383.555 1091.490 2383.925 ;
        RECT 1091.280 2377.880 1091.420 2383.555 ;
        RECT 1091.260 2373.880 1091.540 2377.880 ;
        RECT 1403.560 1326.525 1403.820 1326.670 ;
        RECT 1403.550 1326.155 1403.830 1326.525 ;
        RECT 1749.470 1326.155 1749.750 1326.525 ;
        RECT 1749.540 1325.990 1749.680 1326.155 ;
        RECT 1749.480 1325.670 1749.740 1325.990 ;
        RECT 1406.310 15.115 1406.590 15.485 ;
        RECT 1406.380 2.400 1406.520 15.115 ;
        RECT 1406.170 -4.800 1406.730 2.400 ;
      LAYER via2 ;
        RECT 1091.210 2383.600 1091.490 2383.880 ;
        RECT 1403.550 1326.200 1403.830 1326.480 ;
        RECT 1749.470 1326.200 1749.750 1326.480 ;
        RECT 1406.310 15.160 1406.590 15.440 ;
      LAYER met3 ;
        RECT 1091.185 2383.890 1091.515 2383.905 ;
        RECT 1749.190 2383.890 1749.570 2383.900 ;
        RECT 1091.185 2383.590 1749.570 2383.890 ;
        RECT 1091.185 2383.575 1091.515 2383.590 ;
        RECT 1749.190 2383.580 1749.570 2383.590 ;
        RECT 1403.525 1326.500 1403.855 1326.505 ;
        RECT 1749.445 1326.500 1749.775 1326.505 ;
        RECT 1403.270 1326.490 1403.855 1326.500 ;
        RECT 1403.070 1326.190 1403.855 1326.490 ;
        RECT 1403.270 1326.180 1403.855 1326.190 ;
        RECT 1749.190 1326.490 1749.775 1326.500 ;
        RECT 1749.190 1326.190 1750.000 1326.490 ;
        RECT 1749.190 1326.180 1749.775 1326.190 ;
        RECT 1403.525 1326.175 1403.855 1326.180 ;
        RECT 1749.445 1326.175 1749.775 1326.180 ;
        RECT 1403.270 15.450 1403.650 15.460 ;
        RECT 1406.285 15.450 1406.615 15.465 ;
        RECT 1403.270 15.150 1406.615 15.450 ;
        RECT 1403.270 15.140 1403.650 15.150 ;
        RECT 1406.285 15.135 1406.615 15.150 ;
      LAYER via3 ;
        RECT 1749.220 2383.580 1749.540 2383.900 ;
        RECT 1403.300 1326.180 1403.620 1326.500 ;
        RECT 1749.220 1326.180 1749.540 1326.500 ;
        RECT 1403.300 15.140 1403.620 15.460 ;
      LAYER met4 ;
        RECT 1749.215 2383.575 1749.545 2383.905 ;
        RECT 1749.230 1326.505 1749.530 2383.575 ;
        RECT 1403.295 1326.175 1403.625 1326.505 ;
        RECT 1749.215 1326.175 1749.545 1326.505 ;
        RECT 1403.310 15.465 1403.610 1326.175 ;
        RECT 1403.295 15.135 1403.625 15.465 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1054.850 68.920 1055.170 68.980 ;
        RECT 1421.470 68.920 1421.790 68.980 ;
        RECT 1054.850 68.780 1421.790 68.920 ;
        RECT 1054.850 68.720 1055.170 68.780 ;
        RECT 1421.470 68.720 1421.790 68.780 ;
      LAYER via ;
        RECT 1054.880 68.720 1055.140 68.980 ;
        RECT 1421.500 68.720 1421.760 68.980 ;
      LAYER met2 ;
        RECT 1053.540 1323.690 1053.820 1327.135 ;
        RECT 1053.540 1323.550 1055.080 1323.690 ;
        RECT 1053.540 1323.135 1053.820 1323.550 ;
        RECT 1054.940 69.010 1055.080 1323.550 ;
        RECT 1054.880 68.690 1055.140 69.010 ;
        RECT 1421.500 68.690 1421.760 69.010 ;
        RECT 1421.560 3.130 1421.700 68.690 ;
        RECT 1421.560 2.990 1424.000 3.130 ;
        RECT 1423.860 2.400 1424.000 2.990 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 721.425 997.645 721.595 1089.955 ;
        RECT 720.965 804.525 721.135 855.355 ;
        RECT 721.425 572.645 721.595 622.455 ;
        RECT 721.425 476.085 721.595 524.195 ;
        RECT 721.885 379.525 722.055 451.435 ;
        RECT 720.965 193.885 721.135 245.055 ;
      LAYER mcon ;
        RECT 721.425 1089.785 721.595 1089.955 ;
        RECT 720.965 855.185 721.135 855.355 ;
        RECT 721.425 622.285 721.595 622.455 ;
        RECT 721.425 524.025 721.595 524.195 ;
        RECT 721.885 451.265 722.055 451.435 ;
        RECT 720.965 244.885 721.135 245.055 ;
      LAYER met1 ;
        RECT 717.210 1729.140 717.530 1729.200 ;
        RECT 720.430 1729.140 720.750 1729.200 ;
        RECT 717.210 1729.000 720.750 1729.140 ;
        RECT 717.210 1728.940 717.530 1729.000 ;
        RECT 720.430 1728.940 720.750 1729.000 ;
        RECT 719.510 1567.640 719.830 1567.700 ;
        RECT 720.430 1567.640 720.750 1567.700 ;
        RECT 719.510 1567.500 720.750 1567.640 ;
        RECT 719.510 1567.440 719.830 1567.500 ;
        RECT 720.430 1567.440 720.750 1567.500 ;
        RECT 719.510 1524.800 719.830 1524.860 ;
        RECT 720.430 1524.800 720.750 1524.860 ;
        RECT 719.510 1524.660 720.750 1524.800 ;
        RECT 719.510 1524.600 719.830 1524.660 ;
        RECT 720.430 1524.600 720.750 1524.660 ;
        RECT 721.810 1187.180 722.130 1187.240 ;
        RECT 722.270 1187.180 722.590 1187.240 ;
        RECT 721.810 1187.040 722.590 1187.180 ;
        RECT 721.810 1186.980 722.130 1187.040 ;
        RECT 722.270 1186.980 722.590 1187.040 ;
        RECT 721.350 1138.560 721.670 1138.620 ;
        RECT 722.270 1138.560 722.590 1138.620 ;
        RECT 721.350 1138.420 722.590 1138.560 ;
        RECT 721.350 1138.360 721.670 1138.420 ;
        RECT 722.270 1138.360 722.590 1138.420 ;
        RECT 721.350 1089.940 721.670 1090.000 ;
        RECT 721.155 1089.800 721.670 1089.940 ;
        RECT 721.350 1089.740 721.670 1089.800 ;
        RECT 721.350 997.800 721.670 997.860 ;
        RECT 721.155 997.660 721.670 997.800 ;
        RECT 721.350 997.600 721.670 997.660 ;
        RECT 720.905 855.340 721.195 855.385 ;
        RECT 721.350 855.340 721.670 855.400 ;
        RECT 720.905 855.200 721.670 855.340 ;
        RECT 720.905 855.155 721.195 855.200 ;
        RECT 721.350 855.140 721.670 855.200 ;
        RECT 720.890 804.680 721.210 804.740 ;
        RECT 720.695 804.540 721.210 804.680 ;
        RECT 720.890 804.480 721.210 804.540 ;
        RECT 720.890 759.460 721.210 759.520 ;
        RECT 720.890 759.320 721.580 759.460 ;
        RECT 720.890 759.260 721.210 759.320 ;
        RECT 721.440 759.180 721.580 759.320 ;
        RECT 721.350 758.920 721.670 759.180 ;
        RECT 721.350 686.700 721.670 686.760 ;
        RECT 722.270 686.700 722.590 686.760 ;
        RECT 721.350 686.560 722.590 686.700 ;
        RECT 721.350 686.500 721.670 686.560 ;
        RECT 722.270 686.500 722.590 686.560 ;
        RECT 721.365 622.440 721.655 622.485 ;
        RECT 722.270 622.440 722.590 622.500 ;
        RECT 721.365 622.300 722.590 622.440 ;
        RECT 721.365 622.255 721.655 622.300 ;
        RECT 722.270 622.240 722.590 622.300 ;
        RECT 721.365 572.800 721.655 572.845 ;
        RECT 722.730 572.800 723.050 572.860 ;
        RECT 721.365 572.660 723.050 572.800 ;
        RECT 721.365 572.615 721.655 572.660 ;
        RECT 722.730 572.600 723.050 572.660 ;
        RECT 722.730 531.660 723.050 531.720 ;
        RECT 721.900 531.520 723.050 531.660 ;
        RECT 721.900 531.380 722.040 531.520 ;
        RECT 722.730 531.460 723.050 531.520 ;
        RECT 721.810 531.120 722.130 531.380 ;
        RECT 721.365 524.180 721.655 524.225 ;
        RECT 721.810 524.180 722.130 524.240 ;
        RECT 721.365 524.040 722.130 524.180 ;
        RECT 721.365 523.995 721.655 524.040 ;
        RECT 721.810 523.980 722.130 524.040 ;
        RECT 721.350 476.240 721.670 476.300 ;
        RECT 721.155 476.100 721.670 476.240 ;
        RECT 721.350 476.040 721.670 476.100 ;
        RECT 721.350 451.420 721.670 451.480 ;
        RECT 721.825 451.420 722.115 451.465 ;
        RECT 721.350 451.280 722.115 451.420 ;
        RECT 721.350 451.220 721.670 451.280 ;
        RECT 721.825 451.235 722.115 451.280 ;
        RECT 721.810 379.680 722.130 379.740 ;
        RECT 721.615 379.540 722.130 379.680 ;
        RECT 721.810 379.480 722.130 379.540 ;
        RECT 720.905 245.040 721.195 245.085 ;
        RECT 721.350 245.040 721.670 245.100 ;
        RECT 720.905 244.900 721.670 245.040 ;
        RECT 720.905 244.855 721.195 244.900 ;
        RECT 721.350 244.840 721.670 244.900 ;
        RECT 720.890 194.040 721.210 194.100 ;
        RECT 720.695 193.900 721.210 194.040 ;
        RECT 720.890 193.840 721.210 193.900 ;
        RECT 720.890 186.020 721.210 186.280 ;
        RECT 720.980 185.880 721.120 186.020 ;
        RECT 721.350 185.880 721.670 185.940 ;
        RECT 720.980 185.740 721.670 185.880 ;
        RECT 721.350 185.680 721.670 185.740 ;
        RECT 721.350 137.940 721.670 138.000 ;
        RECT 720.980 137.800 721.670 137.940 ;
        RECT 720.980 137.660 721.120 137.800 ;
        RECT 721.350 137.740 721.670 137.800 ;
        RECT 720.890 137.400 721.210 137.660 ;
        RECT 720.890 53.620 721.210 53.680 ;
        RECT 1441.710 53.620 1442.030 53.680 ;
        RECT 720.890 53.480 1442.030 53.620 ;
        RECT 720.890 53.420 721.210 53.480 ;
        RECT 1441.710 53.420 1442.030 53.480 ;
      LAYER via ;
        RECT 717.240 1728.940 717.500 1729.200 ;
        RECT 720.460 1728.940 720.720 1729.200 ;
        RECT 719.540 1567.440 719.800 1567.700 ;
        RECT 720.460 1567.440 720.720 1567.700 ;
        RECT 719.540 1524.600 719.800 1524.860 ;
        RECT 720.460 1524.600 720.720 1524.860 ;
        RECT 721.840 1186.980 722.100 1187.240 ;
        RECT 722.300 1186.980 722.560 1187.240 ;
        RECT 721.380 1138.360 721.640 1138.620 ;
        RECT 722.300 1138.360 722.560 1138.620 ;
        RECT 721.380 1089.740 721.640 1090.000 ;
        RECT 721.380 997.600 721.640 997.860 ;
        RECT 721.380 855.140 721.640 855.400 ;
        RECT 720.920 804.480 721.180 804.740 ;
        RECT 720.920 759.260 721.180 759.520 ;
        RECT 721.380 758.920 721.640 759.180 ;
        RECT 721.380 686.500 721.640 686.760 ;
        RECT 722.300 686.500 722.560 686.760 ;
        RECT 722.300 622.240 722.560 622.500 ;
        RECT 722.760 572.600 723.020 572.860 ;
        RECT 722.760 531.460 723.020 531.720 ;
        RECT 721.840 531.120 722.100 531.380 ;
        RECT 721.840 523.980 722.100 524.240 ;
        RECT 721.380 476.040 721.640 476.300 ;
        RECT 721.380 451.220 721.640 451.480 ;
        RECT 721.840 379.480 722.100 379.740 ;
        RECT 721.380 244.840 721.640 245.100 ;
        RECT 720.920 193.840 721.180 194.100 ;
        RECT 720.920 186.020 721.180 186.280 ;
        RECT 721.380 185.680 721.640 185.940 ;
        RECT 721.380 137.740 721.640 138.000 ;
        RECT 720.920 137.400 721.180 137.660 ;
        RECT 720.920 53.420 721.180 53.680 ;
        RECT 1441.740 53.420 1442.000 53.680 ;
      LAYER met2 ;
        RECT 717.230 1734.155 717.510 1734.525 ;
        RECT 717.300 1729.230 717.440 1734.155 ;
        RECT 717.240 1728.910 717.500 1729.230 ;
        RECT 720.460 1728.910 720.720 1729.230 ;
        RECT 720.520 1724.210 720.660 1728.910 ;
        RECT 720.520 1724.070 721.120 1724.210 ;
        RECT 719.540 1567.410 719.800 1567.730 ;
        RECT 720.460 1567.640 720.720 1567.730 ;
        RECT 720.980 1567.640 721.120 1724.070 ;
        RECT 720.460 1567.500 721.120 1567.640 ;
        RECT 720.460 1567.410 720.720 1567.500 ;
        RECT 719.600 1524.890 719.740 1567.410 ;
        RECT 719.540 1524.570 719.800 1524.890 ;
        RECT 720.460 1524.800 720.720 1524.890 ;
        RECT 720.460 1524.660 721.120 1524.800 ;
        RECT 720.460 1524.570 720.720 1524.660 ;
        RECT 720.980 1307.370 721.120 1524.660 ;
        RECT 720.980 1307.230 722.040 1307.370 ;
        RECT 721.900 1255.690 722.040 1307.230 ;
        RECT 721.900 1255.550 722.500 1255.690 ;
        RECT 722.360 1187.270 722.500 1255.550 ;
        RECT 721.840 1186.950 722.100 1187.270 ;
        RECT 722.300 1186.950 722.560 1187.270 ;
        RECT 721.900 1173.410 722.040 1186.950 ;
        RECT 721.440 1173.270 722.040 1173.410 ;
        RECT 721.440 1152.445 721.580 1173.270 ;
        RECT 721.370 1152.075 721.650 1152.445 ;
        RECT 722.290 1152.075 722.570 1152.445 ;
        RECT 722.360 1138.650 722.500 1152.075 ;
        RECT 721.380 1138.330 721.640 1138.650 ;
        RECT 722.300 1138.330 722.560 1138.650 ;
        RECT 721.440 1090.030 721.580 1138.330 ;
        RECT 721.380 1089.710 721.640 1090.030 ;
        RECT 721.380 997.570 721.640 997.890 ;
        RECT 721.440 855.430 721.580 997.570 ;
        RECT 721.380 855.110 721.640 855.430 ;
        RECT 720.920 804.450 721.180 804.770 ;
        RECT 720.980 759.550 721.120 804.450 ;
        RECT 720.920 759.230 721.180 759.550 ;
        RECT 721.380 758.890 721.640 759.210 ;
        RECT 721.440 686.790 721.580 758.890 ;
        RECT 721.380 686.470 721.640 686.790 ;
        RECT 722.300 686.470 722.560 686.790 ;
        RECT 722.360 622.530 722.500 686.470 ;
        RECT 722.300 622.210 722.560 622.530 ;
        RECT 722.760 572.570 723.020 572.890 ;
        RECT 722.820 531.750 722.960 572.570 ;
        RECT 722.760 531.430 723.020 531.750 ;
        RECT 721.840 531.090 722.100 531.410 ;
        RECT 721.900 524.270 722.040 531.090 ;
        RECT 721.840 523.950 722.100 524.270 ;
        RECT 721.380 476.010 721.640 476.330 ;
        RECT 721.440 451.510 721.580 476.010 ;
        RECT 721.380 451.190 721.640 451.510 ;
        RECT 721.840 379.450 722.100 379.770 ;
        RECT 721.900 303.690 722.040 379.450 ;
        RECT 721.440 303.550 722.040 303.690 ;
        RECT 721.440 245.130 721.580 303.550 ;
        RECT 721.380 244.810 721.640 245.130 ;
        RECT 720.920 193.810 721.180 194.130 ;
        RECT 720.980 186.310 721.120 193.810 ;
        RECT 720.920 185.990 721.180 186.310 ;
        RECT 721.380 185.650 721.640 185.970 ;
        RECT 721.440 138.030 721.580 185.650 ;
        RECT 721.380 137.710 721.640 138.030 ;
        RECT 720.920 137.370 721.180 137.690 ;
        RECT 720.980 53.710 721.120 137.370 ;
        RECT 720.920 53.390 721.180 53.710 ;
        RECT 1441.740 53.390 1442.000 53.710 ;
        RECT 1441.800 2.400 1441.940 53.390 ;
        RECT 1441.590 -4.800 1442.150 2.400 ;
      LAYER via2 ;
        RECT 717.230 1734.200 717.510 1734.480 ;
        RECT 721.370 1152.120 721.650 1152.400 ;
        RECT 722.290 1152.120 722.570 1152.400 ;
      LAYER met3 ;
        RECT 715.810 1736.615 719.810 1737.215 ;
        RECT 716.990 1734.505 717.290 1736.615 ;
        RECT 716.990 1734.190 717.535 1734.505 ;
        RECT 717.205 1734.175 717.535 1734.190 ;
        RECT 721.345 1152.410 721.675 1152.425 ;
        RECT 722.265 1152.410 722.595 1152.425 ;
        RECT 721.345 1152.110 722.595 1152.410 ;
        RECT 721.345 1152.095 721.675 1152.110 ;
        RECT 722.265 1152.095 722.595 1152.110 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1628.470 2394.520 1628.790 2394.580 ;
        RECT 1676.310 2394.520 1676.630 2394.580 ;
        RECT 1628.470 2394.380 1676.630 2394.520 ;
        RECT 1628.470 2394.320 1628.790 2394.380 ;
        RECT 1676.310 2394.320 1676.630 2394.380 ;
        RECT 1435.270 2394.180 1435.590 2394.240 ;
        RECT 1483.110 2394.180 1483.430 2394.240 ;
        RECT 1435.270 2394.040 1483.430 2394.180 ;
        RECT 1435.270 2393.980 1435.590 2394.040 ;
        RECT 1483.110 2393.980 1483.430 2394.040 ;
        RECT 1531.870 2394.180 1532.190 2394.240 ;
        RECT 1554.870 2394.180 1555.190 2394.240 ;
        RECT 1531.870 2394.040 1555.190 2394.180 ;
        RECT 1531.870 2393.980 1532.190 2394.040 ;
        RECT 1554.870 2393.980 1555.190 2394.040 ;
        RECT 1281.630 2393.500 1281.950 2393.560 ;
        RECT 1289.910 2393.500 1290.230 2393.560 ;
        RECT 1281.630 2393.360 1290.230 2393.500 ;
        RECT 1281.630 2393.300 1281.950 2393.360 ;
        RECT 1289.910 2393.300 1290.230 2393.360 ;
        RECT 1247.590 2388.740 1247.910 2388.800 ;
        RECT 1254.030 2388.740 1254.350 2388.800 ;
        RECT 1247.590 2388.600 1254.350 2388.740 ;
        RECT 1247.590 2388.540 1247.910 2388.600 ;
        RECT 1254.030 2388.540 1254.350 2388.600 ;
      LAYER via ;
        RECT 1628.500 2394.320 1628.760 2394.580 ;
        RECT 1676.340 2394.320 1676.600 2394.580 ;
        RECT 1435.300 2393.980 1435.560 2394.240 ;
        RECT 1483.140 2393.980 1483.400 2394.240 ;
        RECT 1531.900 2393.980 1532.160 2394.240 ;
        RECT 1554.900 2393.980 1555.160 2394.240 ;
        RECT 1281.660 2393.300 1281.920 2393.560 ;
        RECT 1289.940 2393.300 1290.200 2393.560 ;
        RECT 1247.620 2388.540 1247.880 2388.800 ;
        RECT 1254.060 2388.540 1254.320 2388.800 ;
      LAYER met2 ;
        RECT 1628.500 2394.290 1628.760 2394.610 ;
        RECT 1676.340 2394.290 1676.600 2394.610 ;
        RECT 1435.300 2393.950 1435.560 2394.270 ;
        RECT 1483.140 2393.950 1483.400 2394.270 ;
        RECT 1531.900 2393.950 1532.160 2394.270 ;
        RECT 1554.900 2393.950 1555.160 2394.270 ;
        RECT 1281.660 2393.270 1281.920 2393.590 ;
        RECT 1289.940 2393.445 1290.200 2393.590 ;
        RECT 1435.360 2393.445 1435.500 2393.950 ;
        RECT 1483.200 2393.445 1483.340 2393.950 ;
        RECT 1531.960 2393.445 1532.100 2393.950 ;
        RECT 1281.720 2389.365 1281.860 2393.270 ;
        RECT 1289.930 2393.075 1290.210 2393.445 ;
        RECT 1338.690 2393.075 1338.970 2393.445 ;
        RECT 1386.530 2393.075 1386.810 2393.445 ;
        RECT 1435.290 2393.075 1435.570 2393.445 ;
        RECT 1483.130 2393.075 1483.410 2393.445 ;
        RECT 1531.890 2393.075 1532.170 2393.445 ;
        RECT 1338.760 2390.725 1338.900 2393.075 ;
        RECT 1386.600 2390.725 1386.740 2393.075 ;
        RECT 1554.960 2392.765 1555.100 2393.950 ;
        RECT 1628.560 2393.445 1628.700 2394.290 ;
        RECT 1676.400 2393.445 1676.540 2394.290 ;
        RECT 1628.490 2393.075 1628.770 2393.445 ;
        RECT 1676.330 2393.075 1676.610 2393.445 ;
        RECT 1699.790 2393.075 1700.070 2393.445 ;
        RECT 1554.890 2392.395 1555.170 2392.765 ;
        RECT 1338.690 2390.355 1338.970 2390.725 ;
        RECT 1386.530 2390.355 1386.810 2390.725 ;
        RECT 1254.050 2388.995 1254.330 2389.365 ;
        RECT 1281.650 2388.995 1281.930 2389.365 ;
        RECT 1699.860 2389.250 1700.000 2393.075 ;
        RECT 1701.630 2389.930 1701.910 2390.045 ;
        RECT 1701.240 2389.790 1701.910 2389.930 ;
        RECT 1701.240 2389.250 1701.380 2389.790 ;
        RECT 1701.630 2389.675 1701.910 2389.790 ;
        RECT 1699.860 2389.110 1701.380 2389.250 ;
        RECT 1254.120 2388.830 1254.260 2388.995 ;
        RECT 1247.620 2388.510 1247.880 2388.830 ;
        RECT 1254.060 2388.510 1254.320 2388.830 ;
        RECT 1247.680 2377.880 1247.820 2388.510 ;
        RECT 1247.660 2373.880 1247.940 2377.880 ;
        RECT 1459.670 18.515 1459.950 18.885 ;
        RECT 1459.740 2.400 1459.880 18.515 ;
        RECT 1459.530 -4.800 1460.090 2.400 ;
      LAYER via2 ;
        RECT 1289.930 2393.120 1290.210 2393.400 ;
        RECT 1338.690 2393.120 1338.970 2393.400 ;
        RECT 1386.530 2393.120 1386.810 2393.400 ;
        RECT 1435.290 2393.120 1435.570 2393.400 ;
        RECT 1483.130 2393.120 1483.410 2393.400 ;
        RECT 1531.890 2393.120 1532.170 2393.400 ;
        RECT 1628.490 2393.120 1628.770 2393.400 ;
        RECT 1676.330 2393.120 1676.610 2393.400 ;
        RECT 1699.790 2393.120 1700.070 2393.400 ;
        RECT 1554.890 2392.440 1555.170 2392.720 ;
        RECT 1338.690 2390.400 1338.970 2390.680 ;
        RECT 1386.530 2390.400 1386.810 2390.680 ;
        RECT 1254.050 2389.040 1254.330 2389.320 ;
        RECT 1281.650 2389.040 1281.930 2389.320 ;
        RECT 1701.630 2389.720 1701.910 2390.000 ;
        RECT 1459.670 18.560 1459.950 18.840 ;
      LAYER met3 ;
        RECT 1289.905 2393.410 1290.235 2393.425 ;
        RECT 1338.665 2393.410 1338.995 2393.425 ;
        RECT 1289.905 2393.110 1338.995 2393.410 ;
        RECT 1289.905 2393.095 1290.235 2393.110 ;
        RECT 1338.665 2393.095 1338.995 2393.110 ;
        RECT 1386.505 2393.410 1386.835 2393.425 ;
        RECT 1435.265 2393.410 1435.595 2393.425 ;
        RECT 1386.505 2393.110 1435.595 2393.410 ;
        RECT 1386.505 2393.095 1386.835 2393.110 ;
        RECT 1435.265 2393.095 1435.595 2393.110 ;
        RECT 1483.105 2393.410 1483.435 2393.425 ;
        RECT 1531.865 2393.410 1532.195 2393.425 ;
        RECT 1628.465 2393.410 1628.795 2393.425 ;
        RECT 1483.105 2393.110 1532.195 2393.410 ;
        RECT 1483.105 2393.095 1483.435 2393.110 ;
        RECT 1531.865 2393.095 1532.195 2393.110 ;
        RECT 1582.710 2393.110 1628.795 2393.410 ;
        RECT 1554.865 2392.730 1555.195 2392.745 ;
        RECT 1582.710 2392.730 1583.010 2393.110 ;
        RECT 1628.465 2393.095 1628.795 2393.110 ;
        RECT 1676.305 2393.410 1676.635 2393.425 ;
        RECT 1699.765 2393.410 1700.095 2393.425 ;
        RECT 1676.305 2393.110 1700.095 2393.410 ;
        RECT 1676.305 2393.095 1676.635 2393.110 ;
        RECT 1699.765 2393.095 1700.095 2393.110 ;
        RECT 1554.865 2392.430 1583.010 2392.730 ;
        RECT 1554.865 2392.415 1555.195 2392.430 ;
        RECT 1338.665 2390.690 1338.995 2390.705 ;
        RECT 1386.505 2390.690 1386.835 2390.705 ;
        RECT 1338.665 2390.390 1386.835 2390.690 ;
        RECT 1338.665 2390.375 1338.995 2390.390 ;
        RECT 1386.505 2390.375 1386.835 2390.390 ;
        RECT 1701.605 2390.010 1701.935 2390.025 ;
        RECT 1710.550 2390.010 1710.930 2390.020 ;
        RECT 1701.605 2389.710 1710.930 2390.010 ;
        RECT 1701.605 2389.695 1701.935 2389.710 ;
        RECT 1710.550 2389.700 1710.930 2389.710 ;
        RECT 1254.025 2389.330 1254.355 2389.345 ;
        RECT 1281.625 2389.330 1281.955 2389.345 ;
        RECT 1254.025 2389.030 1281.955 2389.330 ;
        RECT 1254.025 2389.015 1254.355 2389.030 ;
        RECT 1281.625 2389.015 1281.955 2389.030 ;
        RECT 1711.470 2369.610 1711.850 2369.620 ;
        RECT 1770.350 2369.610 1770.730 2369.620 ;
        RECT 1711.470 2369.310 1770.730 2369.610 ;
        RECT 1711.470 2369.300 1711.850 2369.310 ;
        RECT 1770.350 2369.300 1770.730 2369.310 ;
        RECT 1764.830 1355.050 1765.210 1355.060 ;
        RECT 1770.350 1355.050 1770.730 1355.060 ;
        RECT 1764.830 1354.750 1770.730 1355.050 ;
        RECT 1764.830 1354.740 1765.210 1354.750 ;
        RECT 1770.350 1354.740 1770.730 1354.750 ;
        RECT 1459.645 18.850 1459.975 18.865 ;
        RECT 1462.150 18.850 1462.530 18.860 ;
        RECT 1459.645 18.550 1462.530 18.850 ;
        RECT 1459.645 18.535 1459.975 18.550 ;
        RECT 1462.150 18.540 1462.530 18.550 ;
      LAYER via3 ;
        RECT 1710.580 2389.700 1710.900 2390.020 ;
        RECT 1711.500 2369.300 1711.820 2369.620 ;
        RECT 1770.380 2369.300 1770.700 2369.620 ;
        RECT 1764.860 1354.740 1765.180 1355.060 ;
        RECT 1770.380 1354.740 1770.700 1355.060 ;
        RECT 1462.180 18.540 1462.500 18.860 ;
      LAYER met4 ;
        RECT 1710.575 2389.695 1710.905 2390.025 ;
        RECT 1710.590 2388.650 1710.890 2389.695 ;
        RECT 1710.590 2388.350 1711.810 2388.650 ;
        RECT 1711.510 2369.625 1711.810 2388.350 ;
        RECT 1711.495 2369.295 1711.825 2369.625 ;
        RECT 1770.375 2369.295 1770.705 2369.625 ;
        RECT 1764.430 1354.310 1765.610 1355.490 ;
        RECT 1770.390 1355.065 1770.690 2369.295 ;
        RECT 1770.375 1354.735 1770.705 1355.065 ;
        RECT 1461.750 1330.510 1462.930 1331.690 ;
        RECT 1462.190 18.865 1462.490 1330.510 ;
        RECT 1462.175 18.535 1462.505 18.865 ;
      LAYER met5 ;
        RECT 1764.220 1352.300 1765.820 1355.700 ;
        RECT 1760.540 1350.700 1765.820 1352.300 ;
        RECT 1760.540 1338.700 1762.140 1350.700 ;
        RECT 1461.540 1337.100 1762.140 1338.700 ;
        RECT 1461.540 1330.300 1463.140 1337.100 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1483.185 1326.425 1483.355 1331.015 ;
      LAYER mcon ;
        RECT 1483.185 1330.845 1483.355 1331.015 ;
      LAYER met1 ;
        RECT 1722.310 2391.800 1722.630 2391.860 ;
        RECT 1783.030 2391.800 1783.350 2391.860 ;
        RECT 1722.310 2391.660 1783.350 2391.800 ;
        RECT 1722.310 2391.600 1722.630 2391.660 ;
        RECT 1783.030 2391.600 1783.350 2391.660 ;
        RECT 1483.125 1331.000 1483.415 1331.045 ;
        RECT 1783.030 1331.000 1783.350 1331.060 ;
        RECT 1483.125 1330.860 1783.350 1331.000 ;
        RECT 1483.125 1330.815 1483.415 1330.860 ;
        RECT 1783.030 1330.800 1783.350 1330.860 ;
        RECT 1483.110 1326.580 1483.430 1326.640 ;
        RECT 1482.915 1326.440 1483.430 1326.580 ;
        RECT 1483.110 1326.380 1483.430 1326.440 ;
        RECT 1477.590 20.640 1477.910 20.700 ;
        RECT 1483.110 20.640 1483.430 20.700 ;
        RECT 1477.590 20.500 1483.430 20.640 ;
        RECT 1477.590 20.440 1477.910 20.500 ;
        RECT 1483.110 20.440 1483.430 20.500 ;
      LAYER via ;
        RECT 1722.340 2391.600 1722.600 2391.860 ;
        RECT 1783.060 2391.600 1783.320 2391.860 ;
        RECT 1783.060 1330.800 1783.320 1331.060 ;
        RECT 1483.140 1326.380 1483.400 1326.640 ;
        RECT 1477.620 20.440 1477.880 20.700 ;
        RECT 1483.140 20.440 1483.400 20.700 ;
      LAYER met2 ;
        RECT 1722.340 2391.570 1722.600 2391.890 ;
        RECT 1783.060 2391.570 1783.320 2391.890 ;
        RECT 1722.400 2377.880 1722.540 2391.570 ;
        RECT 1722.380 2373.880 1722.660 2377.880 ;
        RECT 1783.120 1331.090 1783.260 2391.570 ;
        RECT 1783.060 1330.770 1783.320 1331.090 ;
        RECT 1483.140 1326.350 1483.400 1326.670 ;
        RECT 1483.200 20.730 1483.340 1326.350 ;
        RECT 1477.620 20.410 1477.880 20.730 ;
        RECT 1483.140 20.410 1483.400 20.730 ;
        RECT 1477.680 2.400 1477.820 20.410 ;
        RECT 1477.470 -4.800 1478.030 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 712.685 1553.545 712.855 1562.895 ;
        RECT 717.745 1333.225 717.915 1404.115 ;
        RECT 1491.465 1326.425 1491.635 1333.395 ;
      LAYER mcon ;
        RECT 712.685 1562.725 712.855 1562.895 ;
        RECT 717.745 1403.945 717.915 1404.115 ;
        RECT 1491.465 1333.225 1491.635 1333.395 ;
      LAYER met1 ;
        RECT 713.990 1798.160 714.310 1798.220 ;
        RECT 717.210 1798.160 717.530 1798.220 ;
        RECT 713.990 1798.020 717.530 1798.160 ;
        RECT 713.990 1797.960 714.310 1798.020 ;
        RECT 717.210 1797.960 717.530 1798.020 ;
        RECT 713.990 1657.060 714.310 1657.120 ;
        RECT 717.210 1657.060 717.530 1657.120 ;
        RECT 713.990 1656.920 717.530 1657.060 ;
        RECT 713.990 1656.860 714.310 1656.920 ;
        RECT 717.210 1656.860 717.530 1656.920 ;
        RECT 712.625 1562.880 712.915 1562.925 ;
        RECT 717.210 1562.880 717.530 1562.940 ;
        RECT 712.625 1562.740 717.530 1562.880 ;
        RECT 712.625 1562.695 712.915 1562.740 ;
        RECT 717.210 1562.680 717.530 1562.740 ;
        RECT 712.610 1553.700 712.930 1553.760 ;
        RECT 712.415 1553.560 712.930 1553.700 ;
        RECT 712.610 1553.500 712.930 1553.560 ;
        RECT 717.210 1404.100 717.530 1404.160 ;
        RECT 717.685 1404.100 717.975 1404.145 ;
        RECT 717.210 1403.960 717.975 1404.100 ;
        RECT 717.210 1403.900 717.530 1403.960 ;
        RECT 717.685 1403.915 717.975 1403.960 ;
        RECT 717.685 1333.380 717.975 1333.425 ;
        RECT 1491.405 1333.380 1491.695 1333.425 ;
        RECT 717.685 1333.240 1491.695 1333.380 ;
        RECT 717.685 1333.195 717.975 1333.240 ;
        RECT 1491.405 1333.195 1491.695 1333.240 ;
        RECT 1491.390 1326.580 1491.710 1326.640 ;
        RECT 1491.195 1326.440 1491.710 1326.580 ;
        RECT 1491.390 1326.380 1491.710 1326.440 ;
      LAYER via ;
        RECT 714.020 1797.960 714.280 1798.220 ;
        RECT 717.240 1797.960 717.500 1798.220 ;
        RECT 714.020 1656.860 714.280 1657.120 ;
        RECT 717.240 1656.860 717.500 1657.120 ;
        RECT 717.240 1562.680 717.500 1562.940 ;
        RECT 712.640 1553.500 712.900 1553.760 ;
        RECT 717.240 1403.900 717.500 1404.160 ;
        RECT 1491.420 1326.380 1491.680 1326.640 ;
      LAYER met2 ;
        RECT 813.830 2382.195 814.110 2382.565 ;
        RECT 813.900 2376.445 814.040 2382.195 ;
        RECT 813.830 2376.075 814.110 2376.445 ;
        RECT 893.410 2376.330 893.690 2376.445 ;
        RECT 895.300 2376.330 895.580 2377.880 ;
        RECT 893.410 2376.190 895.580 2376.330 ;
        RECT 893.410 2376.075 893.690 2376.190 ;
        RECT 895.300 2373.880 895.580 2376.190 ;
        RECT 718.610 2242.115 718.890 2242.485 ;
        RECT 718.680 2154.765 718.820 2242.115 ;
        RECT 718.610 2154.395 718.890 2154.765 ;
        RECT 717.690 2101.355 717.970 2101.725 ;
        RECT 717.760 2084.045 717.900 2101.355 ;
        RECT 717.690 2083.675 717.970 2084.045 ;
        RECT 717.230 1950.395 717.510 1950.765 ;
        RECT 717.300 1939.205 717.440 1950.395 ;
        RECT 717.230 1938.835 717.510 1939.205 ;
        RECT 717.230 1927.275 717.510 1927.645 ;
        RECT 717.300 1798.250 717.440 1927.275 ;
        RECT 714.020 1797.930 714.280 1798.250 ;
        RECT 717.240 1797.930 717.500 1798.250 ;
        RECT 714.080 1657.150 714.220 1797.930 ;
        RECT 714.020 1656.830 714.280 1657.150 ;
        RECT 717.240 1656.830 717.500 1657.150 ;
        RECT 717.300 1562.970 717.440 1656.830 ;
        RECT 717.240 1562.650 717.500 1562.970 ;
        RECT 712.640 1553.470 712.900 1553.790 ;
        RECT 712.700 1552.285 712.840 1553.470 ;
        RECT 712.630 1551.915 712.910 1552.285 ;
        RECT 717.230 1404.355 717.510 1404.725 ;
        RECT 717.300 1404.190 717.440 1404.355 ;
        RECT 717.240 1403.870 717.500 1404.190 ;
        RECT 1491.420 1326.350 1491.680 1326.670 ;
        RECT 1491.480 1325.845 1491.620 1326.350 ;
        RECT 1491.410 1325.475 1491.690 1325.845 ;
        RECT 1495.550 18.515 1495.830 18.885 ;
        RECT 1495.620 2.400 1495.760 18.515 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
      LAYER via2 ;
        RECT 813.830 2382.240 814.110 2382.520 ;
        RECT 813.830 2376.120 814.110 2376.400 ;
        RECT 893.410 2376.120 893.690 2376.400 ;
        RECT 718.610 2242.160 718.890 2242.440 ;
        RECT 718.610 2154.440 718.890 2154.720 ;
        RECT 717.690 2101.400 717.970 2101.680 ;
        RECT 717.690 2083.720 717.970 2084.000 ;
        RECT 717.230 1950.440 717.510 1950.720 ;
        RECT 717.230 1938.880 717.510 1939.160 ;
        RECT 717.230 1927.320 717.510 1927.600 ;
        RECT 712.630 1551.960 712.910 1552.240 ;
        RECT 717.230 1404.400 717.510 1404.680 ;
        RECT 1491.410 1325.520 1491.690 1325.800 ;
        RECT 1495.550 18.560 1495.830 18.840 ;
      LAYER met3 ;
        RECT 765.710 2382.530 766.090 2382.540 ;
        RECT 813.805 2382.530 814.135 2382.545 ;
        RECT 765.710 2382.230 814.135 2382.530 ;
        RECT 765.710 2382.220 766.090 2382.230 ;
        RECT 813.805 2382.215 814.135 2382.230 ;
        RECT 717.870 2376.410 718.250 2376.420 ;
        RECT 765.710 2376.410 766.090 2376.420 ;
        RECT 717.870 2376.110 766.090 2376.410 ;
        RECT 717.870 2376.100 718.250 2376.110 ;
        RECT 765.710 2376.100 766.090 2376.110 ;
        RECT 813.805 2376.410 814.135 2376.425 ;
        RECT 820.910 2376.410 821.290 2376.420 ;
        RECT 813.805 2376.110 821.290 2376.410 ;
        RECT 813.805 2376.095 814.135 2376.110 ;
        RECT 820.910 2376.100 821.290 2376.110 ;
        RECT 821.830 2376.410 822.210 2376.420 ;
        RECT 893.385 2376.410 893.715 2376.425 ;
        RECT 821.830 2376.110 893.715 2376.410 ;
        RECT 821.830 2376.100 822.210 2376.110 ;
        RECT 893.385 2376.095 893.715 2376.110 ;
        RECT 718.790 2289.740 719.170 2290.060 ;
        RECT 718.830 2288.020 719.130 2289.740 ;
        RECT 718.790 2287.700 719.170 2288.020 ;
        RECT 718.585 2242.460 718.915 2242.465 ;
        RECT 718.585 2242.450 719.170 2242.460 ;
        RECT 718.360 2242.150 719.170 2242.450 ;
        RECT 718.585 2242.140 719.170 2242.150 ;
        RECT 718.585 2242.135 718.915 2242.140 ;
        RECT 717.870 2154.730 718.250 2154.740 ;
        RECT 718.585 2154.730 718.915 2154.745 ;
        RECT 717.870 2154.430 718.915 2154.730 ;
        RECT 717.870 2154.420 718.250 2154.430 ;
        RECT 718.585 2154.415 718.915 2154.430 ;
        RECT 717.665 2101.700 717.995 2101.705 ;
        RECT 717.665 2101.690 718.250 2101.700 ;
        RECT 717.440 2101.390 718.250 2101.690 ;
        RECT 717.665 2101.380 718.250 2101.390 ;
        RECT 717.665 2101.375 717.995 2101.380 ;
        RECT 717.665 2084.020 717.995 2084.025 ;
        RECT 717.665 2084.010 718.250 2084.020 ;
        RECT 717.440 2083.710 718.250 2084.010 ;
        RECT 717.665 2083.700 718.250 2083.710 ;
        RECT 717.665 2083.695 717.995 2083.700 ;
        RECT 717.870 1955.860 718.250 1956.180 ;
        RECT 717.910 1955.490 718.210 1955.860 ;
        RECT 718.790 1955.490 719.170 1955.500 ;
        RECT 717.910 1955.190 719.170 1955.490 ;
        RECT 718.790 1955.180 719.170 1955.190 ;
        RECT 717.205 1950.730 717.535 1950.745 ;
        RECT 718.790 1950.730 719.170 1950.740 ;
        RECT 717.205 1950.430 719.170 1950.730 ;
        RECT 717.205 1950.415 717.535 1950.430 ;
        RECT 718.790 1950.420 719.170 1950.430 ;
        RECT 717.205 1939.170 717.535 1939.185 ;
        RECT 718.790 1939.170 719.170 1939.180 ;
        RECT 717.205 1938.870 719.170 1939.170 ;
        RECT 717.205 1938.855 717.535 1938.870 ;
        RECT 718.790 1938.860 719.170 1938.870 ;
        RECT 717.205 1927.610 717.535 1927.625 ;
        RECT 718.790 1927.610 719.170 1927.620 ;
        RECT 717.205 1927.310 719.170 1927.610 ;
        RECT 717.205 1927.295 717.535 1927.310 ;
        RECT 718.790 1927.300 719.170 1927.310 ;
        RECT 712.605 1552.250 712.935 1552.265 ;
        RECT 716.030 1552.250 716.410 1552.260 ;
        RECT 712.605 1551.950 716.410 1552.250 ;
        RECT 712.605 1551.935 712.935 1551.950 ;
        RECT 716.030 1551.940 716.410 1551.950 ;
        RECT 717.205 1404.690 717.535 1404.705 ;
        RECT 718.790 1404.690 719.170 1404.700 ;
        RECT 717.205 1404.390 719.170 1404.690 ;
        RECT 717.205 1404.375 717.535 1404.390 ;
        RECT 718.790 1404.380 719.170 1404.390 ;
        RECT 1491.385 1325.810 1491.715 1325.825 ;
        RECT 1493.430 1325.810 1493.810 1325.820 ;
        RECT 1491.385 1325.510 1493.810 1325.810 ;
        RECT 1491.385 1325.495 1491.715 1325.510 ;
        RECT 1493.430 1325.500 1493.810 1325.510 ;
        RECT 1493.430 18.850 1493.810 18.860 ;
        RECT 1495.525 18.850 1495.855 18.865 ;
        RECT 1493.430 18.550 1495.855 18.850 ;
        RECT 1493.430 18.540 1493.810 18.550 ;
        RECT 1495.525 18.535 1495.855 18.550 ;
      LAYER via3 ;
        RECT 765.740 2382.220 766.060 2382.540 ;
        RECT 717.900 2376.100 718.220 2376.420 ;
        RECT 765.740 2376.100 766.060 2376.420 ;
        RECT 820.940 2376.100 821.260 2376.420 ;
        RECT 821.860 2376.100 822.180 2376.420 ;
        RECT 718.820 2289.740 719.140 2290.060 ;
        RECT 718.820 2287.700 719.140 2288.020 ;
        RECT 718.820 2242.140 719.140 2242.460 ;
        RECT 717.900 2154.420 718.220 2154.740 ;
        RECT 717.900 2101.380 718.220 2101.700 ;
        RECT 717.900 2083.700 718.220 2084.020 ;
        RECT 717.900 1955.860 718.220 1956.180 ;
        RECT 718.820 1955.180 719.140 1955.500 ;
        RECT 718.820 1950.420 719.140 1950.740 ;
        RECT 718.820 1938.860 719.140 1939.180 ;
        RECT 718.820 1927.300 719.140 1927.620 ;
        RECT 716.060 1551.940 716.380 1552.260 ;
        RECT 718.820 1404.380 719.140 1404.700 ;
        RECT 1493.460 1325.500 1493.780 1325.820 ;
        RECT 1493.460 18.540 1493.780 18.860 ;
      LAYER met4 ;
        RECT 765.735 2382.215 766.065 2382.545 ;
        RECT 765.750 2376.425 766.050 2382.215 ;
        RECT 717.895 2376.095 718.225 2376.425 ;
        RECT 765.735 2376.095 766.065 2376.425 ;
        RECT 820.935 2376.095 821.265 2376.425 ;
        RECT 821.855 2376.095 822.185 2376.425 ;
        RECT 717.910 2313.850 718.210 2376.095 ;
        RECT 820.950 2375.050 821.250 2376.095 ;
        RECT 821.870 2375.050 822.170 2376.095 ;
        RECT 820.950 2374.750 822.170 2375.050 ;
        RECT 717.910 2313.550 720.050 2313.850 ;
        RECT 718.815 2290.050 719.145 2290.065 ;
        RECT 719.750 2290.050 720.050 2313.550 ;
        RECT 718.815 2289.750 720.050 2290.050 ;
        RECT 718.815 2289.735 719.145 2289.750 ;
        RECT 718.815 2287.695 719.145 2288.025 ;
        RECT 718.830 2283.250 719.130 2287.695 ;
        RECT 718.830 2282.950 720.050 2283.250 ;
        RECT 718.815 2242.450 719.145 2242.465 ;
        RECT 719.750 2242.450 720.050 2282.950 ;
        RECT 718.815 2242.150 720.050 2242.450 ;
        RECT 718.815 2242.135 719.145 2242.150 ;
        RECT 717.895 2154.415 718.225 2154.745 ;
        RECT 717.910 2101.705 718.210 2154.415 ;
        RECT 717.895 2101.375 718.225 2101.705 ;
        RECT 717.895 2083.695 718.225 2084.025 ;
        RECT 717.910 1956.185 718.210 2083.695 ;
        RECT 717.895 1955.855 718.225 1956.185 ;
        RECT 718.815 1955.175 719.145 1955.505 ;
        RECT 718.830 1950.745 719.130 1955.175 ;
        RECT 718.815 1950.415 719.145 1950.745 ;
        RECT 718.815 1938.855 719.145 1939.185 ;
        RECT 718.830 1927.625 719.130 1938.855 ;
        RECT 718.815 1927.295 719.145 1927.625 ;
        RECT 716.055 1551.935 716.385 1552.265 ;
        RECT 716.070 1474.490 716.370 1551.935 ;
        RECT 721.150 1476.770 722.330 1477.890 ;
        RECT 721.150 1476.710 723.730 1476.770 ;
        RECT 721.590 1476.470 723.730 1476.710 ;
        RECT 715.630 1473.310 716.810 1474.490 ;
        RECT 723.430 1426.450 723.730 1476.470 ;
        RECT 718.830 1426.150 723.730 1426.450 ;
        RECT 718.830 1404.705 719.130 1426.150 ;
        RECT 718.815 1404.375 719.145 1404.705 ;
        RECT 1493.455 1325.495 1493.785 1325.825 ;
        RECT 1493.470 18.865 1493.770 1325.495 ;
        RECT 1493.455 18.535 1493.785 18.865 ;
      LAYER met5 ;
        RECT 715.420 1476.500 722.540 1478.100 ;
        RECT 715.420 1473.100 717.020 1476.500 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1234.710 74.360 1235.030 74.420 ;
        RECT 1511.170 74.360 1511.490 74.420 ;
        RECT 1234.710 74.220 1511.490 74.360 ;
        RECT 1234.710 74.160 1235.030 74.220 ;
        RECT 1511.170 74.160 1511.490 74.220 ;
      LAYER via ;
        RECT 1234.740 74.160 1235.000 74.420 ;
        RECT 1511.200 74.160 1511.460 74.420 ;
      LAYER met2 ;
        RECT 1232.940 1323.690 1233.220 1327.135 ;
        RECT 1232.940 1323.550 1234.940 1323.690 ;
        RECT 1232.940 1323.135 1233.220 1323.550 ;
        RECT 1234.800 74.450 1234.940 1323.550 ;
        RECT 1234.740 74.130 1235.000 74.450 ;
        RECT 1511.200 74.130 1511.460 74.450 ;
        RECT 1511.260 7.210 1511.400 74.130 ;
        RECT 1511.260 7.070 1513.240 7.210 ;
        RECT 1513.100 2.400 1513.240 7.070 ;
        RECT 1512.890 -4.800 1513.450 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 707.550 20.640 707.870 20.700 ;
        RECT 710.310 20.640 710.630 20.700 ;
        RECT 707.550 20.500 710.630 20.640 ;
        RECT 707.550 20.440 707.870 20.500 ;
        RECT 710.310 20.440 710.630 20.500 ;
      LAYER via ;
        RECT 707.580 20.440 707.840 20.700 ;
        RECT 710.340 20.440 710.600 20.700 ;
      LAYER met2 ;
        RECT 707.570 1437.675 707.850 1438.045 ;
        RECT 707.640 20.730 707.780 1437.675 ;
        RECT 707.580 20.410 707.840 20.730 ;
        RECT 710.340 20.410 710.600 20.730 ;
        RECT 710.400 2.400 710.540 20.410 ;
        RECT 710.190 -4.800 710.750 2.400 ;
      LAYER via2 ;
        RECT 707.570 1437.720 707.850 1438.000 ;
      LAYER met3 ;
        RECT 707.545 1438.010 707.875 1438.025 ;
        RECT 715.810 1438.010 719.810 1438.015 ;
        RECT 707.545 1437.710 719.810 1438.010 ;
        RECT 707.545 1437.695 707.875 1437.710 ;
        RECT 715.810 1437.415 719.810 1437.710 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 705.250 1286.800 705.570 1286.860 ;
        RECT 1524.970 1286.800 1525.290 1286.860 ;
        RECT 705.250 1286.660 1525.290 1286.800 ;
        RECT 705.250 1286.600 705.570 1286.660 ;
        RECT 1524.970 1286.600 1525.290 1286.660 ;
        RECT 1524.970 37.640 1525.290 37.700 ;
        RECT 1530.950 37.640 1531.270 37.700 ;
        RECT 1524.970 37.500 1531.270 37.640 ;
        RECT 1524.970 37.440 1525.290 37.500 ;
        RECT 1530.950 37.440 1531.270 37.500 ;
      LAYER via ;
        RECT 705.280 1286.600 705.540 1286.860 ;
        RECT 1525.000 1286.600 1525.260 1286.860 ;
        RECT 1525.000 37.440 1525.260 37.700 ;
        RECT 1530.980 37.440 1531.240 37.700 ;
      LAYER met2 ;
        RECT 705.270 1728.715 705.550 1729.085 ;
        RECT 705.340 1393.845 705.480 1728.715 ;
        RECT 705.270 1393.475 705.550 1393.845 ;
        RECT 705.270 1392.115 705.550 1392.485 ;
        RECT 705.340 1286.890 705.480 1392.115 ;
        RECT 705.280 1286.570 705.540 1286.890 ;
        RECT 1525.000 1286.570 1525.260 1286.890 ;
        RECT 1525.060 37.730 1525.200 1286.570 ;
        RECT 1525.000 37.410 1525.260 37.730 ;
        RECT 1530.980 37.410 1531.240 37.730 ;
        RECT 1531.040 2.400 1531.180 37.410 ;
        RECT 1530.830 -4.800 1531.390 2.400 ;
      LAYER via2 ;
        RECT 705.270 1728.760 705.550 1729.040 ;
        RECT 705.270 1393.520 705.550 1393.800 ;
        RECT 705.270 1392.160 705.550 1392.440 ;
      LAYER met3 ;
        RECT 705.245 1729.050 705.575 1729.065 ;
        RECT 715.810 1729.050 719.810 1729.055 ;
        RECT 705.245 1728.750 719.810 1729.050 ;
        RECT 705.245 1728.735 705.575 1728.750 ;
        RECT 715.810 1728.455 719.810 1728.750 ;
        RECT 705.245 1393.810 705.575 1393.825 ;
        RECT 705.030 1393.495 705.575 1393.810 ;
        RECT 705.030 1392.465 705.330 1393.495 ;
        RECT 705.030 1392.150 705.575 1392.465 ;
        RECT 705.245 1392.135 705.575 1392.150 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1547.125 1326.425 1547.295 1329.655 ;
      LAYER mcon ;
        RECT 1547.125 1329.485 1547.295 1329.655 ;
      LAYER met1 ;
        RECT 714.910 1329.640 715.230 1329.700 ;
        RECT 1547.065 1329.640 1547.355 1329.685 ;
        RECT 714.910 1329.500 1547.355 1329.640 ;
        RECT 714.910 1329.440 715.230 1329.500 ;
        RECT 1547.065 1329.455 1547.355 1329.500 ;
        RECT 1547.050 1326.580 1547.370 1326.640 ;
        RECT 1546.855 1326.440 1547.370 1326.580 ;
        RECT 1547.050 1326.380 1547.370 1326.440 ;
      LAYER via ;
        RECT 714.940 1329.440 715.200 1329.700 ;
        RECT 1547.080 1326.380 1547.340 1326.640 ;
      LAYER met2 ;
        RECT 714.930 2301.275 715.210 2301.645 ;
        RECT 715.000 1329.730 715.140 2301.275 ;
        RECT 714.940 1329.410 715.200 1329.730 ;
        RECT 1547.080 1326.350 1547.340 1326.670 ;
        RECT 1547.140 7.210 1547.280 1326.350 ;
        RECT 1547.140 7.070 1549.120 7.210 ;
        RECT 1548.980 2.400 1549.120 7.070 ;
        RECT 1548.770 -4.800 1549.330 2.400 ;
      LAYER via2 ;
        RECT 714.930 2301.320 715.210 2301.600 ;
      LAYER met3 ;
        RECT 714.905 2301.610 715.235 2301.625 ;
        RECT 715.810 2301.610 719.810 2301.615 ;
        RECT 714.905 2301.310 719.810 2301.610 ;
        RECT 714.905 2301.295 715.235 2301.310 ;
        RECT 715.810 2301.015 719.810 2301.310 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1140.870 1311.280 1141.190 1311.340 ;
        RECT 1144.550 1311.280 1144.870 1311.340 ;
        RECT 1140.870 1311.140 1144.870 1311.280 ;
        RECT 1140.870 1311.080 1141.190 1311.140 ;
        RECT 1144.550 1311.080 1144.870 1311.140 ;
        RECT 1144.550 74.020 1144.870 74.080 ;
        RECT 1566.370 74.020 1566.690 74.080 ;
        RECT 1144.550 73.880 1566.690 74.020 ;
        RECT 1144.550 73.820 1144.870 73.880 ;
        RECT 1566.370 73.820 1566.690 73.880 ;
      LAYER via ;
        RECT 1140.900 1311.080 1141.160 1311.340 ;
        RECT 1144.580 1311.080 1144.840 1311.340 ;
        RECT 1144.580 73.820 1144.840 74.080 ;
        RECT 1566.400 73.820 1566.660 74.080 ;
      LAYER met2 ;
        RECT 1140.940 1323.135 1141.220 1327.135 ;
        RECT 1140.960 1311.370 1141.100 1323.135 ;
        RECT 1140.900 1311.050 1141.160 1311.370 ;
        RECT 1144.580 1311.050 1144.840 1311.370 ;
        RECT 1144.640 74.110 1144.780 1311.050 ;
        RECT 1144.580 73.790 1144.840 74.110 ;
        RECT 1566.400 73.790 1566.660 74.110 ;
        RECT 1566.460 3.130 1566.600 73.790 ;
        RECT 1566.460 2.990 1567.060 3.130 ;
        RECT 1566.920 2.400 1567.060 2.990 ;
        RECT 1566.710 -4.800 1567.270 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1586.685 1326.425 1586.855 1329.655 ;
      LAYER mcon ;
        RECT 1586.685 1329.485 1586.855 1329.655 ;
      LAYER met1 ;
        RECT 1772.910 2190.520 1773.230 2190.580 ;
        RECT 1785.790 2190.520 1786.110 2190.580 ;
        RECT 1772.910 2190.380 1786.110 2190.520 ;
        RECT 1772.910 2190.320 1773.230 2190.380 ;
        RECT 1785.790 2190.320 1786.110 2190.380 ;
        RECT 1586.625 1329.640 1586.915 1329.685 ;
        RECT 1785.790 1329.640 1786.110 1329.700 ;
        RECT 1586.625 1329.500 1786.110 1329.640 ;
        RECT 1586.625 1329.455 1586.915 1329.500 ;
        RECT 1785.790 1329.440 1786.110 1329.500 ;
        RECT 1586.610 1326.580 1586.930 1326.640 ;
        RECT 1586.415 1326.440 1586.930 1326.580 ;
        RECT 1586.610 1326.380 1586.930 1326.440 ;
        RECT 1584.770 2.960 1585.090 3.020 ;
        RECT 1586.610 2.960 1586.930 3.020 ;
        RECT 1584.770 2.820 1586.930 2.960 ;
        RECT 1584.770 2.760 1585.090 2.820 ;
        RECT 1586.610 2.760 1586.930 2.820 ;
      LAYER via ;
        RECT 1772.940 2190.320 1773.200 2190.580 ;
        RECT 1785.820 2190.320 1786.080 2190.580 ;
        RECT 1785.820 1329.440 1786.080 1329.700 ;
        RECT 1586.640 1326.380 1586.900 1326.640 ;
        RECT 1584.800 2.760 1585.060 3.020 ;
        RECT 1586.640 2.760 1586.900 3.020 ;
      LAYER met2 ;
        RECT 1772.930 2193.835 1773.210 2194.205 ;
        RECT 1773.000 2190.610 1773.140 2193.835 ;
        RECT 1772.940 2190.290 1773.200 2190.610 ;
        RECT 1785.820 2190.290 1786.080 2190.610 ;
        RECT 1785.880 1329.730 1786.020 2190.290 ;
        RECT 1785.820 1329.410 1786.080 1329.730 ;
        RECT 1586.640 1326.350 1586.900 1326.670 ;
        RECT 1586.700 3.050 1586.840 1326.350 ;
        RECT 1584.800 2.730 1585.060 3.050 ;
        RECT 1586.640 2.730 1586.900 3.050 ;
        RECT 1584.860 2.400 1585.000 2.730 ;
        RECT 1584.650 -4.800 1585.210 2.400 ;
      LAYER via2 ;
        RECT 1772.930 2193.880 1773.210 2194.160 ;
      LAYER met3 ;
        RECT 1755.835 2194.170 1759.835 2194.175 ;
        RECT 1772.905 2194.170 1773.235 2194.185 ;
        RECT 1755.835 2193.870 1773.235 2194.170 ;
        RECT 1755.835 2193.575 1759.835 2193.870 ;
        RECT 1772.905 2193.855 1773.235 2193.870 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 710.385 1309.085 710.555 1328.295 ;
      LAYER mcon ;
        RECT 710.385 1328.125 710.555 1328.295 ;
      LAYER met1 ;
        RECT 710.310 1328.280 710.630 1328.340 ;
        RECT 710.115 1328.140 710.630 1328.280 ;
        RECT 710.310 1328.080 710.630 1328.140 ;
        RECT 710.325 1309.240 710.615 1309.285 ;
        RECT 710.325 1309.100 742.740 1309.240 ;
        RECT 710.325 1309.055 710.615 1309.100 ;
        RECT 742.600 1308.900 742.740 1309.100 ;
        RECT 1600.870 1308.900 1601.190 1308.960 ;
        RECT 742.600 1308.760 1601.190 1308.900 ;
        RECT 1600.870 1308.700 1601.190 1308.760 ;
      LAYER via ;
        RECT 710.340 1328.080 710.600 1328.340 ;
        RECT 1600.900 1308.700 1601.160 1308.960 ;
      LAYER met2 ;
        RECT 710.330 1523.355 710.610 1523.725 ;
        RECT 710.400 1328.370 710.540 1523.355 ;
        RECT 710.340 1328.050 710.600 1328.370 ;
        RECT 1600.900 1308.670 1601.160 1308.990 ;
        RECT 1600.960 3.130 1601.100 1308.670 ;
        RECT 1600.960 2.990 1602.480 3.130 ;
        RECT 1602.340 2.400 1602.480 2.990 ;
        RECT 1602.130 -4.800 1602.690 2.400 ;
      LAYER via2 ;
        RECT 710.330 1523.400 710.610 1523.680 ;
      LAYER met3 ;
        RECT 710.305 1523.690 710.635 1523.705 ;
        RECT 715.810 1523.690 719.810 1523.695 ;
        RECT 710.305 1523.390 719.810 1523.690 ;
        RECT 710.305 1523.375 710.635 1523.390 ;
        RECT 715.810 1523.095 719.810 1523.390 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1577.870 2374.120 1578.190 2374.180 ;
        RECT 1774.750 2374.120 1775.070 2374.180 ;
        RECT 1577.870 2373.980 1775.070 2374.120 ;
        RECT 1577.870 2373.920 1578.190 2373.980 ;
        RECT 1774.750 2373.920 1775.070 2373.980 ;
        RECT 1620.190 16.900 1620.510 16.960 ;
        RECT 1774.750 16.900 1775.070 16.960 ;
        RECT 1620.190 16.760 1775.070 16.900 ;
        RECT 1620.190 16.700 1620.510 16.760 ;
        RECT 1774.750 16.700 1775.070 16.760 ;
      LAYER via ;
        RECT 1577.900 2373.920 1578.160 2374.180 ;
        RECT 1774.780 2373.920 1775.040 2374.180 ;
        RECT 1620.220 16.700 1620.480 16.960 ;
        RECT 1774.780 16.700 1775.040 16.960 ;
      LAYER met2 ;
        RECT 1577.940 2374.210 1578.220 2377.880 ;
        RECT 1577.900 2373.890 1578.220 2374.210 ;
        RECT 1774.780 2373.890 1775.040 2374.210 ;
        RECT 1577.940 2373.880 1578.220 2373.890 ;
        RECT 1774.840 16.990 1774.980 2373.890 ;
        RECT 1620.220 16.670 1620.480 16.990 ;
        RECT 1774.780 16.670 1775.040 16.990 ;
        RECT 1620.280 2.400 1620.420 16.670 ;
        RECT 1620.070 -4.800 1620.630 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1754.125 2377.875 1754.295 2378.215 ;
        RECT 1753.205 2377.705 1754.295 2377.875 ;
      LAYER mcon ;
        RECT 1754.125 2378.045 1754.295 2378.215 ;
      LAYER met1 ;
        RECT 1754.065 2378.200 1754.355 2378.245 ;
        RECT 1780.730 2378.200 1781.050 2378.260 ;
        RECT 1754.065 2378.060 1781.050 2378.200 ;
        RECT 1754.065 2378.015 1754.355 2378.060 ;
        RECT 1780.730 2378.000 1781.050 2378.060 ;
        RECT 1386.050 2377.860 1386.370 2377.920 ;
        RECT 1753.145 2377.860 1753.435 2377.905 ;
        RECT 1386.050 2377.720 1753.435 2377.860 ;
        RECT 1386.050 2377.660 1386.370 2377.720 ;
        RECT 1753.145 2377.675 1753.435 2377.720 ;
        RECT 1638.130 15.880 1638.450 15.940 ;
        RECT 1780.270 15.880 1780.590 15.940 ;
        RECT 1638.130 15.740 1780.590 15.880 ;
        RECT 1638.130 15.680 1638.450 15.740 ;
        RECT 1780.270 15.680 1780.590 15.740 ;
      LAYER via ;
        RECT 1780.760 2378.000 1781.020 2378.260 ;
        RECT 1386.080 2377.660 1386.340 2377.920 ;
        RECT 1638.160 15.680 1638.420 15.940 ;
        RECT 1780.300 15.680 1780.560 15.940 ;
      LAYER met2 ;
        RECT 1780.760 2377.970 1781.020 2378.290 ;
        RECT 1386.080 2377.690 1386.340 2377.950 ;
        RECT 1386.580 2377.690 1386.860 2377.880 ;
        RECT 1386.080 2377.630 1386.860 2377.690 ;
        RECT 1386.140 2377.550 1386.860 2377.630 ;
        RECT 1386.580 2373.880 1386.860 2377.550 ;
        RECT 1780.820 21.490 1780.960 2377.970 ;
        RECT 1780.360 21.350 1780.960 21.490 ;
        RECT 1780.360 15.970 1780.500 21.350 ;
        RECT 1638.160 15.650 1638.420 15.970 ;
        RECT 1780.300 15.650 1780.560 15.970 ;
        RECT 1638.220 2.400 1638.360 15.650 ;
        RECT 1638.010 -4.800 1638.570 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1757.805 1340.705 1757.975 1342.575 ;
        RECT 1733.425 1326.425 1733.595 1327.615 ;
      LAYER mcon ;
        RECT 1757.805 1342.405 1757.975 1342.575 ;
        RECT 1733.425 1327.445 1733.595 1327.615 ;
      LAYER met1 ;
        RECT 1757.730 1342.560 1758.050 1342.620 ;
        RECT 1757.535 1342.420 1758.050 1342.560 ;
        RECT 1757.730 1342.360 1758.050 1342.420 ;
        RECT 1756.810 1340.860 1757.130 1340.920 ;
        RECT 1757.745 1340.860 1758.035 1340.905 ;
        RECT 1756.810 1340.720 1758.035 1340.860 ;
        RECT 1756.810 1340.660 1757.130 1340.720 ;
        RECT 1757.745 1340.675 1758.035 1340.720 ;
        RECT 1733.365 1327.600 1733.655 1327.645 ;
        RECT 1756.350 1327.600 1756.670 1327.660 ;
        RECT 1733.365 1327.460 1756.670 1327.600 ;
        RECT 1733.365 1327.415 1733.655 1327.460 ;
        RECT 1756.350 1327.400 1756.670 1327.460 ;
        RECT 1662.510 1326.580 1662.830 1326.640 ;
        RECT 1733.365 1326.580 1733.655 1326.625 ;
        RECT 1662.510 1326.440 1733.655 1326.580 ;
        RECT 1662.510 1326.380 1662.830 1326.440 ;
        RECT 1733.365 1326.395 1733.655 1326.440 ;
        RECT 1656.070 18.940 1656.390 19.000 ;
        RECT 1662.510 18.940 1662.830 19.000 ;
        RECT 1656.070 18.800 1662.830 18.940 ;
        RECT 1656.070 18.740 1656.390 18.800 ;
        RECT 1662.510 18.740 1662.830 18.800 ;
      LAYER via ;
        RECT 1757.760 1342.360 1758.020 1342.620 ;
        RECT 1756.840 1340.660 1757.100 1340.920 ;
        RECT 1756.380 1327.400 1756.640 1327.660 ;
        RECT 1662.540 1326.380 1662.800 1326.640 ;
        RECT 1656.100 18.740 1656.360 19.000 ;
        RECT 1662.540 18.740 1662.800 19.000 ;
      LAYER met2 ;
        RECT 1758.210 1636.235 1758.490 1636.605 ;
        RECT 1758.280 1623.570 1758.420 1636.235 ;
        RECT 1757.820 1623.430 1758.420 1623.570 ;
        RECT 1757.820 1342.650 1757.960 1623.430 ;
        RECT 1757.760 1342.330 1758.020 1342.650 ;
        RECT 1756.840 1340.630 1757.100 1340.950 ;
        RECT 1756.900 1328.450 1757.040 1340.630 ;
        RECT 1756.440 1328.310 1757.040 1328.450 ;
        RECT 1756.440 1327.690 1756.580 1328.310 ;
        RECT 1756.380 1327.370 1756.640 1327.690 ;
        RECT 1662.540 1326.350 1662.800 1326.670 ;
        RECT 1662.600 19.030 1662.740 1326.350 ;
        RECT 1656.100 18.710 1656.360 19.030 ;
        RECT 1662.540 18.710 1662.800 19.030 ;
        RECT 1656.160 2.400 1656.300 18.710 ;
        RECT 1655.950 -4.800 1656.510 2.400 ;
      LAYER via2 ;
        RECT 1758.210 1636.280 1758.490 1636.560 ;
      LAYER met3 ;
        RECT 1755.835 1638.695 1759.835 1639.295 ;
        RECT 1758.430 1636.585 1758.730 1638.695 ;
        RECT 1758.185 1636.270 1758.730 1636.585 ;
        RECT 1758.185 1636.255 1758.515 1636.270 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1181.350 1311.280 1181.670 1311.340 ;
        RECT 1185.490 1311.280 1185.810 1311.340 ;
        RECT 1181.350 1311.140 1185.810 1311.280 ;
        RECT 1181.350 1311.080 1181.670 1311.140 ;
        RECT 1185.490 1311.080 1185.810 1311.140 ;
        RECT 1185.490 73.680 1185.810 73.740 ;
        RECT 1669.870 73.680 1670.190 73.740 ;
        RECT 1185.490 73.540 1670.190 73.680 ;
        RECT 1185.490 73.480 1185.810 73.540 ;
        RECT 1669.870 73.480 1670.190 73.540 ;
      LAYER via ;
        RECT 1181.380 1311.080 1181.640 1311.340 ;
        RECT 1185.520 1311.080 1185.780 1311.340 ;
        RECT 1185.520 73.480 1185.780 73.740 ;
        RECT 1669.900 73.480 1670.160 73.740 ;
      LAYER met2 ;
        RECT 1181.420 1323.135 1181.700 1327.135 ;
        RECT 1181.440 1311.370 1181.580 1323.135 ;
        RECT 1181.380 1311.050 1181.640 1311.370 ;
        RECT 1185.520 1311.050 1185.780 1311.370 ;
        RECT 1185.580 73.770 1185.720 1311.050 ;
        RECT 1185.520 73.450 1185.780 73.770 ;
        RECT 1669.900 73.450 1670.160 73.770 ;
        RECT 1669.960 7.210 1670.100 73.450 ;
        RECT 1669.960 7.070 1673.780 7.210 ;
        RECT 1673.640 2.400 1673.780 7.070 ;
        RECT 1673.430 -4.800 1673.990 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1690.645 1326.085 1690.815 1329.315 ;
      LAYER mcon ;
        RECT 1690.645 1329.145 1690.815 1329.315 ;
      LAYER met1 ;
        RECT 704.330 1355.140 704.650 1355.200 ;
        RECT 706.170 1355.140 706.490 1355.200 ;
        RECT 704.330 1355.000 706.490 1355.140 ;
        RECT 704.330 1354.940 704.650 1355.000 ;
        RECT 706.170 1354.940 706.490 1355.000 ;
        RECT 706.170 1329.300 706.490 1329.360 ;
        RECT 1690.585 1329.300 1690.875 1329.345 ;
        RECT 706.170 1329.160 1690.875 1329.300 ;
        RECT 706.170 1329.100 706.490 1329.160 ;
        RECT 1690.585 1329.115 1690.875 1329.160 ;
        RECT 1690.570 1326.240 1690.890 1326.300 ;
        RECT 1690.375 1326.100 1690.890 1326.240 ;
        RECT 1690.570 1326.040 1690.890 1326.100 ;
      LAYER via ;
        RECT 704.360 1354.940 704.620 1355.200 ;
        RECT 706.200 1354.940 706.460 1355.200 ;
        RECT 706.200 1329.100 706.460 1329.360 ;
        RECT 1690.600 1326.040 1690.860 1326.300 ;
      LAYER met2 ;
        RECT 704.350 1531.515 704.630 1531.885 ;
        RECT 704.420 1393.845 704.560 1531.515 ;
        RECT 704.350 1393.475 704.630 1393.845 ;
        RECT 704.350 1392.795 704.630 1393.165 ;
        RECT 704.420 1355.230 704.560 1392.795 ;
        RECT 704.360 1354.910 704.620 1355.230 ;
        RECT 706.200 1354.910 706.460 1355.230 ;
        RECT 706.260 1329.390 706.400 1354.910 ;
        RECT 706.200 1329.070 706.460 1329.390 ;
        RECT 1690.600 1326.010 1690.860 1326.330 ;
        RECT 1690.660 16.730 1690.800 1326.010 ;
        RECT 1690.660 16.590 1691.720 16.730 ;
        RECT 1691.580 2.400 1691.720 16.590 ;
        RECT 1691.370 -4.800 1691.930 2.400 ;
      LAYER via2 ;
        RECT 704.350 1531.560 704.630 1531.840 ;
        RECT 704.350 1393.520 704.630 1393.800 ;
        RECT 704.350 1392.840 704.630 1393.120 ;
      LAYER met3 ;
        RECT 704.325 1531.850 704.655 1531.865 ;
        RECT 715.810 1531.850 719.810 1531.855 ;
        RECT 704.325 1531.550 719.810 1531.850 ;
        RECT 704.325 1531.535 704.655 1531.550 ;
        RECT 715.810 1531.255 719.810 1531.550 ;
        RECT 704.325 1393.495 704.655 1393.825 ;
        RECT 704.340 1393.145 704.640 1393.495 ;
        RECT 704.325 1392.815 704.655 1393.145 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1756.425 1325.745 1756.595 1349.375 ;
      LAYER mcon ;
        RECT 1756.425 1349.205 1756.595 1349.375 ;
      LAYER met1 ;
        RECT 1756.365 1349.360 1756.655 1349.405 ;
        RECT 1756.810 1349.360 1757.130 1349.420 ;
        RECT 1756.365 1349.220 1757.130 1349.360 ;
        RECT 1756.365 1349.175 1756.655 1349.220 ;
        RECT 1756.810 1349.160 1757.130 1349.220 ;
        RECT 1756.350 1325.900 1756.670 1325.960 ;
        RECT 1756.155 1325.760 1756.670 1325.900 ;
        RECT 1756.350 1325.700 1756.670 1325.760 ;
      LAYER via ;
        RECT 1756.840 1349.160 1757.100 1349.420 ;
        RECT 1756.380 1325.700 1756.640 1325.960 ;
      LAYER met2 ;
        RECT 1756.830 1367.635 1757.110 1368.005 ;
        RECT 1756.900 1349.450 1757.040 1367.635 ;
        RECT 1756.840 1349.130 1757.100 1349.450 ;
        RECT 1756.380 1325.670 1756.640 1325.990 ;
        RECT 1756.440 1325.165 1756.580 1325.670 ;
        RECT 1756.370 1324.795 1756.650 1325.165 ;
        RECT 729.190 51.155 729.470 51.525 ;
        RECT 729.260 18.770 729.400 51.155 ;
        RECT 728.340 18.630 729.400 18.770 ;
        RECT 728.340 2.400 728.480 18.630 ;
        RECT 728.130 -4.800 728.690 2.400 ;
      LAYER via2 ;
        RECT 1756.830 1367.680 1757.110 1367.960 ;
        RECT 1756.370 1324.840 1756.650 1325.120 ;
        RECT 729.190 51.200 729.470 51.480 ;
      LAYER met3 ;
        RECT 1755.835 2133.735 1759.835 2134.335 ;
        RECT 1756.590 2132.300 1756.890 2133.735 ;
        RECT 1756.550 2131.980 1756.930 2132.300 ;
        RECT 1758.390 1950.420 1758.770 1950.740 ;
        RECT 1756.550 1949.370 1756.930 1949.380 ;
        RECT 1758.430 1949.370 1758.730 1950.420 ;
        RECT 1756.550 1949.070 1758.730 1949.370 ;
        RECT 1756.550 1949.060 1756.930 1949.070 ;
        RECT 1756.805 1367.980 1757.135 1367.985 ;
        RECT 1756.550 1367.970 1757.135 1367.980 ;
        RECT 1756.550 1367.670 1757.360 1367.970 ;
        RECT 1756.550 1367.660 1757.135 1367.670 ;
        RECT 1756.805 1367.655 1757.135 1367.660 ;
        RECT 1753.830 1325.140 1755.050 1325.300 ;
        RECT 1753.790 1325.130 1755.050 1325.140 ;
        RECT 1756.345 1325.130 1756.675 1325.145 ;
        RECT 1753.790 1325.000 1756.675 1325.130 ;
        RECT 1753.790 1324.820 1754.170 1325.000 ;
        RECT 1754.750 1324.830 1756.675 1325.000 ;
        RECT 1756.345 1324.815 1756.675 1324.830 ;
        RECT 1753.790 910.330 1754.170 910.340 ;
        RECT 1752.910 910.030 1754.170 910.330 ;
        RECT 1752.910 908.980 1753.210 910.030 ;
        RECT 1753.790 910.020 1754.170 910.030 ;
        RECT 1752.870 908.660 1753.250 908.980 ;
        RECT 1753.790 858.650 1754.170 858.660 ;
        RECT 1756.550 858.650 1756.930 858.660 ;
        RECT 1753.790 858.350 1756.930 858.650 ;
        RECT 1753.790 858.340 1754.170 858.350 ;
        RECT 1756.550 858.340 1756.930 858.350 ;
        RECT 1754.710 403.050 1755.090 403.060 ;
        RECT 1758.390 403.050 1758.770 403.060 ;
        RECT 1754.710 402.750 1758.770 403.050 ;
        RECT 1754.710 402.740 1755.090 402.750 ;
        RECT 1758.390 402.740 1758.770 402.750 ;
        RECT 1753.790 348.650 1754.170 348.660 ;
        RECT 1758.390 348.650 1758.770 348.660 ;
        RECT 1753.790 348.350 1758.770 348.650 ;
        RECT 1753.790 348.340 1754.170 348.350 ;
        RECT 1758.390 348.340 1758.770 348.350 ;
        RECT 1753.790 303.090 1754.170 303.100 ;
        RECT 1755.630 303.090 1756.010 303.100 ;
        RECT 1753.790 302.790 1756.010 303.090 ;
        RECT 1753.790 302.780 1754.170 302.790 ;
        RECT 1755.630 302.780 1756.010 302.790 ;
        RECT 1755.630 158.930 1756.010 158.940 ;
        RECT 1758.390 158.930 1758.770 158.940 ;
        RECT 1755.630 158.630 1758.770 158.930 ;
        RECT 1755.630 158.620 1756.010 158.630 ;
        RECT 1758.390 158.620 1758.770 158.630 ;
        RECT 1754.710 134.450 1755.090 134.460 ;
        RECT 1758.390 134.450 1758.770 134.460 ;
        RECT 1754.710 134.150 1758.770 134.450 ;
        RECT 1754.710 134.140 1755.090 134.150 ;
        RECT 1758.390 134.140 1758.770 134.150 ;
        RECT 729.165 51.490 729.495 51.505 ;
        RECT 1756.550 51.490 1756.930 51.500 ;
        RECT 729.165 51.190 1756.930 51.490 ;
        RECT 729.165 51.175 729.495 51.190 ;
        RECT 1756.550 51.180 1756.930 51.190 ;
      LAYER via3 ;
        RECT 1756.580 2131.980 1756.900 2132.300 ;
        RECT 1758.420 1950.420 1758.740 1950.740 ;
        RECT 1756.580 1949.060 1756.900 1949.380 ;
        RECT 1756.580 1367.660 1756.900 1367.980 ;
        RECT 1753.820 1324.820 1754.140 1325.140 ;
        RECT 1753.820 910.020 1754.140 910.340 ;
        RECT 1752.900 908.660 1753.220 908.980 ;
        RECT 1753.820 858.340 1754.140 858.660 ;
        RECT 1756.580 858.340 1756.900 858.660 ;
        RECT 1754.740 402.740 1755.060 403.060 ;
        RECT 1758.420 402.740 1758.740 403.060 ;
        RECT 1753.820 348.340 1754.140 348.660 ;
        RECT 1758.420 348.340 1758.740 348.660 ;
        RECT 1753.820 302.780 1754.140 303.100 ;
        RECT 1755.660 302.780 1755.980 303.100 ;
        RECT 1755.660 158.620 1755.980 158.940 ;
        RECT 1758.420 158.620 1758.740 158.940 ;
        RECT 1754.740 134.140 1755.060 134.460 ;
        RECT 1758.420 134.140 1758.740 134.460 ;
        RECT 1756.580 51.180 1756.900 51.500 ;
      LAYER met4 ;
        RECT 1756.575 2131.975 1756.905 2132.305 ;
        RECT 1756.590 2072.450 1756.890 2131.975 ;
        RECT 1756.590 2072.150 1758.040 2072.450 ;
        RECT 1757.740 2069.050 1758.040 2072.150 ;
        RECT 1757.510 2068.750 1758.040 2069.050 ;
        RECT 1757.510 2055.450 1757.810 2068.750 ;
        RECT 1752.910 2055.150 1757.810 2055.450 ;
        RECT 1752.910 2027.570 1753.210 2055.150 ;
        RECT 1752.910 2027.270 1758.730 2027.570 ;
        RECT 1758.430 1950.745 1758.730 2027.270 ;
        RECT 1758.415 1950.415 1758.745 1950.745 ;
        RECT 1756.575 1949.055 1756.905 1949.385 ;
        RECT 1756.590 1946.650 1756.890 1949.055 ;
        RECT 1752.910 1946.350 1756.890 1946.650 ;
        RECT 1752.910 1939.850 1753.210 1946.350 ;
        RECT 1751.070 1939.550 1753.210 1939.850 ;
        RECT 1751.070 1926.250 1751.370 1939.550 ;
        RECT 1751.070 1925.950 1754.130 1926.250 ;
        RECT 1753.830 1909.250 1754.130 1925.950 ;
        RECT 1753.830 1908.950 1756.890 1909.250 ;
        RECT 1756.590 1878.650 1756.890 1908.950 ;
        RECT 1756.590 1878.350 1757.580 1878.650 ;
        RECT 1757.280 1875.250 1757.580 1878.350 ;
        RECT 1756.590 1874.950 1757.580 1875.250 ;
        RECT 1756.590 1868.450 1756.890 1874.950 ;
        RECT 1755.670 1868.150 1756.890 1868.450 ;
        RECT 1755.670 1844.650 1755.970 1868.150 ;
        RECT 1753.830 1844.350 1755.970 1844.650 ;
        RECT 1753.830 1841.930 1754.130 1844.350 ;
        RECT 1752.910 1841.630 1754.130 1841.930 ;
        RECT 1752.910 1817.450 1753.210 1841.630 ;
        RECT 1752.910 1817.150 1755.050 1817.450 ;
        RECT 1754.750 1769.850 1755.050 1817.150 ;
        RECT 1753.830 1769.550 1755.050 1769.850 ;
        RECT 1753.830 1579.450 1754.130 1769.550 ;
        RECT 1752.910 1579.150 1754.130 1579.450 ;
        RECT 1752.910 1535.250 1753.210 1579.150 ;
        RECT 1752.910 1534.950 1755.050 1535.250 ;
        RECT 1754.750 1525.050 1755.050 1534.950 ;
        RECT 1753.830 1524.750 1755.050 1525.050 ;
        RECT 1753.830 1406.730 1754.130 1524.750 ;
        RECT 1753.830 1406.430 1755.970 1406.730 ;
        RECT 1755.670 1395.850 1755.970 1406.430 ;
        RECT 1753.830 1395.550 1755.970 1395.850 ;
        RECT 1753.830 1375.450 1754.130 1395.550 ;
        RECT 1753.830 1375.150 1755.050 1375.450 ;
        RECT 1754.750 1368.650 1755.050 1375.150 ;
        RECT 1754.750 1368.350 1756.660 1368.650 ;
        RECT 1756.360 1367.985 1756.660 1368.350 ;
        RECT 1756.360 1367.670 1756.905 1367.985 ;
        RECT 1756.575 1367.655 1756.905 1367.670 ;
        RECT 1753.815 1324.815 1754.145 1325.145 ;
        RECT 1753.830 1293.850 1754.130 1324.815 ;
        RECT 1752.910 1293.550 1754.130 1293.850 ;
        RECT 1752.910 1246.250 1753.210 1293.550 ;
        RECT 1752.910 1245.950 1754.130 1246.250 ;
        RECT 1753.830 910.345 1754.130 1245.950 ;
        RECT 1753.815 910.015 1754.145 910.345 ;
        RECT 1752.895 908.655 1753.225 908.985 ;
        RECT 1752.910 862.050 1753.210 908.655 ;
        RECT 1752.910 861.750 1754.130 862.050 ;
        RECT 1753.830 858.665 1754.130 861.750 ;
        RECT 1753.815 858.335 1754.145 858.665 ;
        RECT 1756.575 858.335 1756.905 858.665 ;
        RECT 1756.590 794.050 1756.890 858.335 ;
        RECT 1753.830 793.750 1756.890 794.050 ;
        RECT 1753.830 712.450 1754.130 793.750 ;
        RECT 1753.830 712.150 1755.970 712.450 ;
        RECT 1755.670 664.850 1755.970 712.150 ;
        RECT 1754.750 664.550 1755.970 664.850 ;
        RECT 1754.750 620.650 1755.050 664.550 ;
        RECT 1754.750 620.350 1755.970 620.650 ;
        RECT 1755.670 569.650 1755.970 620.350 ;
        RECT 1754.750 569.350 1755.970 569.650 ;
        RECT 1754.750 522.050 1755.050 569.350 ;
        RECT 1754.750 521.750 1755.970 522.050 ;
        RECT 1755.670 474.450 1755.970 521.750 ;
        RECT 1754.750 474.150 1755.970 474.450 ;
        RECT 1754.750 403.065 1755.050 474.150 ;
        RECT 1754.735 402.735 1755.065 403.065 ;
        RECT 1758.415 402.735 1758.745 403.065 ;
        RECT 1758.430 348.665 1758.730 402.735 ;
        RECT 1753.815 348.335 1754.145 348.665 ;
        RECT 1758.415 348.335 1758.745 348.665 ;
        RECT 1753.830 303.105 1754.130 348.335 ;
        RECT 1753.815 302.775 1754.145 303.105 ;
        RECT 1755.655 302.775 1755.985 303.105 ;
        RECT 1755.670 280.650 1755.970 302.775 ;
        RECT 1754.750 280.350 1755.970 280.650 ;
        RECT 1754.750 209.250 1755.050 280.350 ;
        RECT 1754.750 208.950 1755.970 209.250 ;
        RECT 1755.670 158.945 1755.970 208.950 ;
        RECT 1755.655 158.615 1755.985 158.945 ;
        RECT 1758.415 158.615 1758.745 158.945 ;
        RECT 1758.430 134.465 1758.730 158.615 ;
        RECT 1754.735 134.135 1755.065 134.465 ;
        RECT 1758.415 134.135 1758.745 134.465 ;
        RECT 1754.750 83.450 1755.050 134.135 ;
        RECT 1754.750 83.150 1756.890 83.450 ;
        RECT 1756.590 51.505 1756.890 83.150 ;
        RECT 1756.575 51.175 1756.905 51.505 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1675.465 689.265 1675.635 717.655 ;
        RECT 1675.465 593.045 1675.635 627.895 ;
        RECT 1675.925 544.765 1676.095 579.615 ;
        RECT 1675.925 483.225 1676.095 531.335 ;
        RECT 1675.925 434.945 1676.095 482.715 ;
        RECT 1676.385 186.405 1676.555 234.515 ;
        RECT 1675.465 89.165 1675.635 131.155 ;
        RECT 1675.465 41.565 1675.635 62.475 ;
      LAYER mcon ;
        RECT 1675.465 717.485 1675.635 717.655 ;
        RECT 1675.465 627.725 1675.635 627.895 ;
        RECT 1675.925 579.445 1676.095 579.615 ;
        RECT 1675.925 531.165 1676.095 531.335 ;
        RECT 1675.925 482.545 1676.095 482.715 ;
        RECT 1676.385 234.345 1676.555 234.515 ;
        RECT 1675.465 130.985 1675.635 131.155 ;
        RECT 1675.465 62.305 1675.635 62.475 ;
      LAYER met1 ;
        RECT 1674.010 1311.280 1674.330 1311.340 ;
        RECT 1676.310 1311.280 1676.630 1311.340 ;
        RECT 1674.010 1311.140 1676.630 1311.280 ;
        RECT 1674.010 1311.080 1674.330 1311.140 ;
        RECT 1676.310 1311.080 1676.630 1311.140 ;
        RECT 1675.850 883.700 1676.170 883.960 ;
        RECT 1675.940 882.940 1676.080 883.700 ;
        RECT 1675.850 882.680 1676.170 882.940 ;
        RECT 1675.390 773.060 1675.710 773.120 ;
        RECT 1675.850 773.060 1676.170 773.120 ;
        RECT 1675.390 772.920 1676.170 773.060 ;
        RECT 1675.390 772.860 1675.710 772.920 ;
        RECT 1675.850 772.860 1676.170 772.920 ;
        RECT 1675.850 738.720 1676.170 738.780 ;
        RECT 1675.480 738.580 1676.170 738.720 ;
        RECT 1675.480 738.100 1675.620 738.580 ;
        RECT 1675.850 738.520 1676.170 738.580 ;
        RECT 1675.390 737.840 1675.710 738.100 ;
        RECT 1675.390 717.640 1675.710 717.700 ;
        RECT 1675.195 717.500 1675.710 717.640 ;
        RECT 1675.390 717.440 1675.710 717.500 ;
        RECT 1675.405 689.420 1675.695 689.465 ;
        RECT 1675.850 689.420 1676.170 689.480 ;
        RECT 1675.405 689.280 1676.170 689.420 ;
        RECT 1675.405 689.235 1675.695 689.280 ;
        RECT 1675.850 689.220 1676.170 689.280 ;
        RECT 1674.930 627.880 1675.250 627.940 ;
        RECT 1675.405 627.880 1675.695 627.925 ;
        RECT 1674.930 627.740 1675.695 627.880 ;
        RECT 1674.930 627.680 1675.250 627.740 ;
        RECT 1675.405 627.695 1675.695 627.740 ;
        RECT 1675.390 593.200 1675.710 593.260 ;
        RECT 1675.195 593.060 1675.710 593.200 ;
        RECT 1675.390 593.000 1675.710 593.060 ;
        RECT 1675.850 579.600 1676.170 579.660 ;
        RECT 1675.655 579.460 1676.170 579.600 ;
        RECT 1675.850 579.400 1676.170 579.460 ;
        RECT 1675.850 544.920 1676.170 544.980 ;
        RECT 1675.655 544.780 1676.170 544.920 ;
        RECT 1675.850 544.720 1676.170 544.780 ;
        RECT 1675.850 531.320 1676.170 531.380 ;
        RECT 1675.655 531.180 1676.170 531.320 ;
        RECT 1675.850 531.120 1676.170 531.180 ;
        RECT 1675.850 483.380 1676.170 483.440 ;
        RECT 1675.655 483.240 1676.170 483.380 ;
        RECT 1675.850 483.180 1676.170 483.240 ;
        RECT 1675.850 482.700 1676.170 482.760 ;
        RECT 1675.655 482.560 1676.170 482.700 ;
        RECT 1675.850 482.500 1676.170 482.560 ;
        RECT 1675.850 435.100 1676.170 435.160 ;
        RECT 1675.655 434.960 1676.170 435.100 ;
        RECT 1675.850 434.900 1676.170 434.960 ;
        RECT 1675.850 400.560 1676.170 400.820 ;
        RECT 1675.940 400.140 1676.080 400.560 ;
        RECT 1675.850 399.880 1676.170 400.140 ;
        RECT 1675.850 241.440 1676.170 241.700 ;
        RECT 1675.390 241.300 1675.710 241.360 ;
        RECT 1675.940 241.300 1676.080 241.440 ;
        RECT 1675.390 241.160 1676.080 241.300 ;
        RECT 1675.390 241.100 1675.710 241.160 ;
        RECT 1676.310 234.500 1676.630 234.560 ;
        RECT 1676.115 234.360 1676.630 234.500 ;
        RECT 1676.310 234.300 1676.630 234.360 ;
        RECT 1676.310 186.560 1676.630 186.620 ;
        RECT 1676.115 186.420 1676.630 186.560 ;
        RECT 1676.310 186.360 1676.630 186.420 ;
        RECT 1675.390 131.140 1675.710 131.200 ;
        RECT 1675.195 131.000 1675.710 131.140 ;
        RECT 1675.390 130.940 1675.710 131.000 ;
        RECT 1675.390 89.320 1675.710 89.380 ;
        RECT 1675.195 89.180 1675.710 89.320 ;
        RECT 1675.390 89.120 1675.710 89.180 ;
        RECT 1675.390 62.460 1675.710 62.520 ;
        RECT 1675.195 62.320 1675.710 62.460 ;
        RECT 1675.390 62.260 1675.710 62.320 ;
        RECT 1675.390 41.720 1675.710 41.780 ;
        RECT 1675.195 41.580 1675.710 41.720 ;
        RECT 1675.390 41.520 1675.710 41.580 ;
        RECT 1675.390 24.040 1675.710 24.100 ;
        RECT 1709.430 24.040 1709.750 24.100 ;
        RECT 1675.390 23.900 1709.750 24.040 ;
        RECT 1675.390 23.840 1675.710 23.900 ;
        RECT 1709.430 23.840 1709.750 23.900 ;
      LAYER via ;
        RECT 1674.040 1311.080 1674.300 1311.340 ;
        RECT 1676.340 1311.080 1676.600 1311.340 ;
        RECT 1675.880 883.700 1676.140 883.960 ;
        RECT 1675.880 882.680 1676.140 882.940 ;
        RECT 1675.420 772.860 1675.680 773.120 ;
        RECT 1675.880 772.860 1676.140 773.120 ;
        RECT 1675.880 738.520 1676.140 738.780 ;
        RECT 1675.420 737.840 1675.680 738.100 ;
        RECT 1675.420 717.440 1675.680 717.700 ;
        RECT 1675.880 689.220 1676.140 689.480 ;
        RECT 1674.960 627.680 1675.220 627.940 ;
        RECT 1675.420 593.000 1675.680 593.260 ;
        RECT 1675.880 579.400 1676.140 579.660 ;
        RECT 1675.880 544.720 1676.140 544.980 ;
        RECT 1675.880 531.120 1676.140 531.380 ;
        RECT 1675.880 483.180 1676.140 483.440 ;
        RECT 1675.880 482.500 1676.140 482.760 ;
        RECT 1675.880 434.900 1676.140 435.160 ;
        RECT 1675.880 400.560 1676.140 400.820 ;
        RECT 1675.880 399.880 1676.140 400.140 ;
        RECT 1675.880 241.440 1676.140 241.700 ;
        RECT 1675.420 241.100 1675.680 241.360 ;
        RECT 1676.340 234.300 1676.600 234.560 ;
        RECT 1676.340 186.360 1676.600 186.620 ;
        RECT 1675.420 130.940 1675.680 131.200 ;
        RECT 1675.420 89.120 1675.680 89.380 ;
        RECT 1675.420 62.260 1675.680 62.520 ;
        RECT 1675.420 41.520 1675.680 41.780 ;
        RECT 1675.420 23.840 1675.680 24.100 ;
        RECT 1709.460 23.840 1709.720 24.100 ;
      LAYER met2 ;
        RECT 1672.700 1323.690 1672.980 1327.135 ;
        RECT 1672.700 1323.550 1674.240 1323.690 ;
        RECT 1672.700 1323.135 1672.980 1323.550 ;
        RECT 1674.100 1311.370 1674.240 1323.550 ;
        RECT 1674.040 1311.050 1674.300 1311.370 ;
        RECT 1676.340 1311.050 1676.600 1311.370 ;
        RECT 1676.400 1269.290 1676.540 1311.050 ;
        RECT 1675.940 1269.150 1676.540 1269.290 ;
        RECT 1675.940 1221.690 1676.080 1269.150 ;
        RECT 1675.480 1221.550 1676.080 1221.690 ;
        RECT 1675.480 1221.010 1675.620 1221.550 ;
        RECT 1675.480 1220.870 1676.080 1221.010 ;
        RECT 1675.940 1173.410 1676.080 1220.870 ;
        RECT 1675.940 1173.270 1676.540 1173.410 ;
        RECT 1676.400 1172.730 1676.540 1173.270 ;
        RECT 1675.940 1172.590 1676.540 1172.730 ;
        RECT 1675.940 1125.130 1676.080 1172.590 ;
        RECT 1675.480 1124.990 1676.080 1125.130 ;
        RECT 1675.480 1124.450 1675.620 1124.990 ;
        RECT 1675.480 1124.310 1676.080 1124.450 ;
        RECT 1675.940 1076.850 1676.080 1124.310 ;
        RECT 1675.940 1076.710 1676.540 1076.850 ;
        RECT 1676.400 1076.170 1676.540 1076.710 ;
        RECT 1675.940 1076.030 1676.540 1076.170 ;
        RECT 1675.940 1028.570 1676.080 1076.030 ;
        RECT 1675.480 1028.430 1676.080 1028.570 ;
        RECT 1675.480 1027.890 1675.620 1028.430 ;
        RECT 1675.480 1027.750 1676.080 1027.890 ;
        RECT 1675.940 980.290 1676.080 1027.750 ;
        RECT 1675.940 980.150 1676.540 980.290 ;
        RECT 1676.400 979.610 1676.540 980.150 ;
        RECT 1675.940 979.470 1676.540 979.610 ;
        RECT 1675.940 932.010 1676.080 979.470 ;
        RECT 1675.480 931.870 1676.080 932.010 ;
        RECT 1675.480 931.330 1675.620 931.870 ;
        RECT 1675.480 931.190 1676.080 931.330 ;
        RECT 1675.940 883.990 1676.080 931.190 ;
        RECT 1675.880 883.670 1676.140 883.990 ;
        RECT 1675.880 882.650 1676.140 882.970 ;
        RECT 1675.940 835.450 1676.080 882.650 ;
        RECT 1675.480 835.310 1676.080 835.450 ;
        RECT 1675.480 834.770 1675.620 835.310 ;
        RECT 1675.480 834.630 1676.080 834.770 ;
        RECT 1675.940 787.170 1676.080 834.630 ;
        RECT 1675.480 787.030 1676.080 787.170 ;
        RECT 1675.480 773.150 1675.620 787.030 ;
        RECT 1675.420 772.830 1675.680 773.150 ;
        RECT 1675.880 772.830 1676.140 773.150 ;
        RECT 1675.940 738.810 1676.080 772.830 ;
        RECT 1675.880 738.490 1676.140 738.810 ;
        RECT 1675.420 737.810 1675.680 738.130 ;
        RECT 1675.480 717.730 1675.620 737.810 ;
        RECT 1675.420 717.410 1675.680 717.730 ;
        RECT 1675.880 689.190 1676.140 689.510 ;
        RECT 1675.940 651.850 1676.080 689.190 ;
        RECT 1675.020 651.710 1676.080 651.850 ;
        RECT 1675.020 627.970 1675.160 651.710 ;
        RECT 1674.960 627.650 1675.220 627.970 ;
        RECT 1675.420 592.970 1675.680 593.290 ;
        RECT 1675.480 579.770 1675.620 592.970 ;
        RECT 1675.480 579.690 1676.080 579.770 ;
        RECT 1675.480 579.630 1676.140 579.690 ;
        RECT 1675.880 579.370 1676.140 579.630 ;
        RECT 1675.940 579.215 1676.080 579.370 ;
        RECT 1675.880 544.690 1676.140 545.010 ;
        RECT 1675.940 531.410 1676.080 544.690 ;
        RECT 1675.880 531.090 1676.140 531.410 ;
        RECT 1675.880 483.150 1676.140 483.470 ;
        RECT 1675.940 482.790 1676.080 483.150 ;
        RECT 1675.880 482.470 1676.140 482.790 ;
        RECT 1675.880 434.870 1676.140 435.190 ;
        RECT 1675.940 400.850 1676.080 434.870 ;
        RECT 1675.880 400.530 1676.140 400.850 ;
        RECT 1675.880 399.850 1676.140 400.170 ;
        RECT 1675.940 351.970 1676.080 399.850 ;
        RECT 1675.480 351.830 1676.080 351.970 ;
        RECT 1675.480 351.290 1675.620 351.830 ;
        RECT 1675.480 351.150 1676.080 351.290 ;
        RECT 1675.940 241.730 1676.080 351.150 ;
        RECT 1675.880 241.410 1676.140 241.730 ;
        RECT 1675.420 241.070 1675.680 241.390 ;
        RECT 1675.480 235.125 1675.620 241.070 ;
        RECT 1675.410 234.755 1675.690 235.125 ;
        RECT 1676.330 234.755 1676.610 235.125 ;
        RECT 1676.400 234.590 1676.540 234.755 ;
        RECT 1676.340 234.270 1676.600 234.590 ;
        RECT 1676.340 186.330 1676.600 186.650 ;
        RECT 1676.400 162.250 1676.540 186.330 ;
        RECT 1675.480 162.110 1676.540 162.250 ;
        RECT 1675.480 131.230 1675.620 162.110 ;
        RECT 1675.420 130.910 1675.680 131.230 ;
        RECT 1675.420 89.090 1675.680 89.410 ;
        RECT 1675.480 62.550 1675.620 89.090 ;
        RECT 1675.420 62.230 1675.680 62.550 ;
        RECT 1675.420 41.490 1675.680 41.810 ;
        RECT 1675.480 24.130 1675.620 41.490 ;
        RECT 1675.420 23.810 1675.680 24.130 ;
        RECT 1709.460 23.810 1709.720 24.130 ;
        RECT 1709.520 2.400 1709.660 23.810 ;
        RECT 1709.310 -4.800 1709.870 2.400 ;
      LAYER via2 ;
        RECT 1675.410 234.800 1675.690 235.080 ;
        RECT 1676.330 234.800 1676.610 235.080 ;
      LAYER met3 ;
        RECT 1675.385 235.090 1675.715 235.105 ;
        RECT 1676.305 235.090 1676.635 235.105 ;
        RECT 1675.385 234.790 1676.635 235.090 ;
        RECT 1675.385 234.775 1675.715 234.790 ;
        RECT 1676.305 234.775 1676.635 234.790 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1341.890 2377.520 1342.210 2377.580 ;
        RECT 1752.670 2377.520 1752.990 2377.580 ;
        RECT 1341.890 2377.380 1752.990 2377.520 ;
        RECT 1341.890 2377.320 1342.210 2377.380 ;
        RECT 1752.670 2377.320 1752.990 2377.380 ;
        RECT 1727.370 14.520 1727.690 14.580 ;
        RECT 1774.290 14.520 1774.610 14.580 ;
        RECT 1727.370 14.380 1774.610 14.520 ;
        RECT 1727.370 14.320 1727.690 14.380 ;
        RECT 1774.290 14.320 1774.610 14.380 ;
      LAYER via ;
        RECT 1341.920 2377.320 1342.180 2377.580 ;
        RECT 1752.700 2377.320 1752.960 2377.580 ;
        RECT 1727.400 14.320 1727.660 14.580 ;
        RECT 1774.320 14.320 1774.580 14.580 ;
      LAYER met2 ;
        RECT 1340.580 2377.690 1340.860 2377.880 ;
        RECT 1340.580 2377.610 1342.120 2377.690 ;
        RECT 1340.580 2377.550 1342.180 2377.610 ;
        RECT 1340.580 2373.880 1340.860 2377.550 ;
        RECT 1341.920 2377.290 1342.180 2377.550 ;
        RECT 1752.700 2377.290 1752.960 2377.610 ;
        RECT 1752.760 2373.725 1752.900 2377.290 ;
        RECT 1752.690 2373.355 1752.970 2373.725 ;
        RECT 1774.310 2373.355 1774.590 2373.725 ;
        RECT 1774.380 14.610 1774.520 2373.355 ;
        RECT 1727.400 14.290 1727.660 14.610 ;
        RECT 1774.320 14.290 1774.580 14.610 ;
        RECT 1727.460 2.400 1727.600 14.290 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
      LAYER via2 ;
        RECT 1752.690 2373.400 1752.970 2373.680 ;
        RECT 1774.310 2373.400 1774.590 2373.680 ;
      LAYER met3 ;
        RECT 1752.665 2373.690 1752.995 2373.705 ;
        RECT 1774.285 2373.690 1774.615 2373.705 ;
        RECT 1752.665 2373.390 1774.615 2373.690 ;
        RECT 1752.665 2373.375 1752.995 2373.390 ;
        RECT 1774.285 2373.375 1774.615 2373.390 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1757.345 1324.725 1757.515 1343.935 ;
        RECT 1744.005 48.365 1744.175 62.815 ;
      LAYER mcon ;
        RECT 1757.345 1343.765 1757.515 1343.935 ;
        RECT 1744.005 62.645 1744.175 62.815 ;
      LAYER met1 ;
        RECT 1757.270 1343.920 1757.590 1343.980 ;
        RECT 1757.075 1343.780 1757.590 1343.920 ;
        RECT 1757.270 1343.720 1757.590 1343.780 ;
        RECT 1744.850 1324.880 1745.170 1324.940 ;
        RECT 1757.285 1324.880 1757.575 1324.925 ;
        RECT 1744.850 1324.740 1757.575 1324.880 ;
        RECT 1744.850 1324.680 1745.170 1324.740 ;
        RECT 1757.285 1324.695 1757.575 1324.740 ;
        RECT 1743.930 717.640 1744.250 717.700 ;
        RECT 1744.850 717.640 1745.170 717.700 ;
        RECT 1743.930 717.500 1745.170 717.640 ;
        RECT 1743.930 717.440 1744.250 717.500 ;
        RECT 1744.850 717.440 1745.170 717.500 ;
        RECT 1743.945 62.800 1744.235 62.845 ;
        RECT 1744.850 62.800 1745.170 62.860 ;
        RECT 1743.945 62.660 1745.170 62.800 ;
        RECT 1743.945 62.615 1744.235 62.660 ;
        RECT 1744.850 62.600 1745.170 62.660 ;
        RECT 1743.930 48.520 1744.250 48.580 ;
        RECT 1743.735 48.380 1744.250 48.520 ;
        RECT 1743.930 48.320 1744.250 48.380 ;
      LAYER via ;
        RECT 1757.300 1343.720 1757.560 1343.980 ;
        RECT 1744.880 1324.680 1745.140 1324.940 ;
        RECT 1743.960 717.440 1744.220 717.700 ;
        RECT 1744.880 717.440 1745.140 717.700 ;
        RECT 1744.880 62.600 1745.140 62.860 ;
        RECT 1743.960 48.320 1744.220 48.580 ;
      LAYER met2 ;
        RECT 1757.290 1823.915 1757.570 1824.285 ;
        RECT 1757.360 1344.010 1757.500 1823.915 ;
        RECT 1757.300 1343.690 1757.560 1344.010 ;
        RECT 1744.880 1324.650 1745.140 1324.970 ;
        RECT 1744.940 717.730 1745.080 1324.650 ;
        RECT 1743.960 717.410 1744.220 717.730 ;
        RECT 1744.880 717.410 1745.140 717.730 ;
        RECT 1744.020 669.645 1744.160 717.410 ;
        RECT 1743.950 669.275 1744.230 669.645 ;
        RECT 1744.870 669.275 1745.150 669.645 ;
        RECT 1744.940 62.890 1745.080 669.275 ;
        RECT 1744.880 62.570 1745.140 62.890 ;
        RECT 1743.960 48.290 1744.220 48.610 ;
        RECT 1744.020 18.090 1744.160 48.290 ;
        RECT 1744.020 17.950 1745.540 18.090 ;
        RECT 1745.400 2.400 1745.540 17.950 ;
        RECT 1745.190 -4.800 1745.750 2.400 ;
      LAYER via2 ;
        RECT 1757.290 1823.960 1757.570 1824.240 ;
        RECT 1743.950 669.320 1744.230 669.600 ;
        RECT 1744.870 669.320 1745.150 669.600 ;
      LAYER met3 ;
        RECT 1755.835 1826.375 1759.835 1826.975 ;
        RECT 1756.590 1824.250 1756.890 1826.375 ;
        RECT 1757.265 1824.250 1757.595 1824.265 ;
        RECT 1756.590 1823.950 1757.595 1824.250 ;
        RECT 1757.265 1823.935 1757.595 1823.950 ;
        RECT 1743.925 669.610 1744.255 669.625 ;
        RECT 1744.845 669.610 1745.175 669.625 ;
        RECT 1743.925 669.310 1745.175 669.610 ;
        RECT 1743.925 669.295 1744.255 669.310 ;
        RECT 1744.845 669.295 1745.175 669.310 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1001.950 1311.280 1002.270 1311.340 ;
        RECT 1006.550 1311.280 1006.870 1311.340 ;
        RECT 1001.950 1311.140 1006.870 1311.280 ;
        RECT 1001.950 1311.080 1002.270 1311.140 ;
        RECT 1006.550 1311.080 1006.870 1311.140 ;
        RECT 1006.550 25.740 1006.870 25.800 ;
        RECT 1762.790 25.740 1763.110 25.800 ;
        RECT 1006.550 25.600 1763.110 25.740 ;
        RECT 1006.550 25.540 1006.870 25.600 ;
        RECT 1762.790 25.540 1763.110 25.600 ;
      LAYER via ;
        RECT 1001.980 1311.080 1002.240 1311.340 ;
        RECT 1006.580 1311.080 1006.840 1311.340 ;
        RECT 1006.580 25.540 1006.840 25.800 ;
        RECT 1762.820 25.540 1763.080 25.800 ;
      LAYER met2 ;
        RECT 1002.020 1323.135 1002.300 1327.135 ;
        RECT 1002.040 1311.370 1002.180 1323.135 ;
        RECT 1001.980 1311.050 1002.240 1311.370 ;
        RECT 1006.580 1311.050 1006.840 1311.370 ;
        RECT 1006.640 25.830 1006.780 1311.050 ;
        RECT 1006.580 25.510 1006.840 25.830 ;
        RECT 1762.820 25.510 1763.080 25.830 ;
        RECT 1762.880 2.400 1763.020 25.510 ;
        RECT 1762.670 -4.800 1763.230 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1507.950 2379.220 1508.270 2379.280 ;
        RECT 1776.590 2379.220 1776.910 2379.280 ;
        RECT 1507.950 2379.080 1776.910 2379.220 ;
        RECT 1507.950 2379.020 1508.270 2379.080 ;
        RECT 1776.590 2379.020 1776.910 2379.080 ;
        RECT 1776.590 20.640 1776.910 20.700 ;
        RECT 1780.730 20.640 1781.050 20.700 ;
        RECT 1776.590 20.500 1781.050 20.640 ;
        RECT 1776.590 20.440 1776.910 20.500 ;
        RECT 1780.730 20.440 1781.050 20.500 ;
      LAYER via ;
        RECT 1507.980 2379.020 1508.240 2379.280 ;
        RECT 1776.620 2379.020 1776.880 2379.280 ;
        RECT 1776.620 20.440 1776.880 20.700 ;
        RECT 1780.760 20.440 1781.020 20.700 ;
      LAYER met2 ;
        RECT 1507.980 2378.990 1508.240 2379.310 ;
        RECT 1776.620 2378.990 1776.880 2379.310 ;
        RECT 1508.040 2377.880 1508.180 2378.990 ;
        RECT 1508.020 2373.880 1508.300 2377.880 ;
        RECT 1776.680 20.730 1776.820 2378.990 ;
        RECT 1776.620 20.410 1776.880 20.730 ;
        RECT 1780.760 20.410 1781.020 20.730 ;
        RECT 1780.820 2.400 1780.960 20.410 ;
        RECT 1780.610 -4.800 1781.170 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1798.745 2.805 1798.915 25.415 ;
      LAYER mcon ;
        RECT 1798.745 25.245 1798.915 25.415 ;
      LAYER met1 ;
        RECT 717.210 1328.620 717.530 1328.680 ;
        RECT 1794.070 1328.620 1794.390 1328.680 ;
        RECT 717.210 1328.480 1794.390 1328.620 ;
        RECT 717.210 1328.420 717.530 1328.480 ;
        RECT 1794.070 1328.420 1794.390 1328.480 ;
        RECT 1794.070 25.400 1794.390 25.460 ;
        RECT 1798.685 25.400 1798.975 25.445 ;
        RECT 1794.070 25.260 1798.975 25.400 ;
        RECT 1794.070 25.200 1794.390 25.260 ;
        RECT 1798.685 25.215 1798.975 25.260 ;
        RECT 1798.670 2.960 1798.990 3.020 ;
        RECT 1798.475 2.820 1798.990 2.960 ;
        RECT 1798.670 2.760 1798.990 2.820 ;
      LAYER via ;
        RECT 717.240 1328.420 717.500 1328.680 ;
        RECT 1794.100 1328.420 1794.360 1328.680 ;
        RECT 1794.100 25.200 1794.360 25.460 ;
        RECT 1798.700 2.760 1798.960 3.020 ;
      LAYER met2 ;
        RECT 717.230 1349.275 717.510 1349.645 ;
        RECT 717.300 1328.710 717.440 1349.275 ;
        RECT 717.240 1328.390 717.500 1328.710 ;
        RECT 1794.100 1328.390 1794.360 1328.710 ;
        RECT 1794.160 25.490 1794.300 1328.390 ;
        RECT 1794.100 25.170 1794.360 25.490 ;
        RECT 1798.700 2.730 1798.960 3.050 ;
        RECT 1798.760 2.400 1798.900 2.730 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
      LAYER via2 ;
        RECT 717.230 1349.320 717.510 1349.600 ;
      LAYER met3 ;
        RECT 715.810 1351.735 719.810 1352.335 ;
        RECT 716.990 1349.625 717.290 1351.735 ;
        RECT 716.990 1349.310 717.535 1349.625 ;
        RECT 717.205 1349.295 717.535 1349.310 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1394.790 1311.280 1395.110 1311.340 ;
        RECT 1399.390 1311.280 1399.710 1311.340 ;
        RECT 1394.790 1311.140 1399.710 1311.280 ;
        RECT 1394.790 1311.080 1395.110 1311.140 ;
        RECT 1399.390 1311.080 1399.710 1311.140 ;
        RECT 1399.390 80.820 1399.710 80.880 ;
        RECT 1814.770 80.820 1815.090 80.880 ;
        RECT 1399.390 80.680 1815.090 80.820 ;
        RECT 1399.390 80.620 1399.710 80.680 ;
        RECT 1814.770 80.620 1815.090 80.680 ;
      LAYER via ;
        RECT 1394.820 1311.080 1395.080 1311.340 ;
        RECT 1399.420 1311.080 1399.680 1311.340 ;
        RECT 1399.420 80.620 1399.680 80.880 ;
        RECT 1814.800 80.620 1815.060 80.880 ;
      LAYER met2 ;
        RECT 1394.860 1323.135 1395.140 1327.135 ;
        RECT 1394.880 1311.370 1395.020 1323.135 ;
        RECT 1394.820 1311.050 1395.080 1311.370 ;
        RECT 1399.420 1311.050 1399.680 1311.370 ;
        RECT 1399.480 80.910 1399.620 1311.050 ;
        RECT 1399.420 80.590 1399.680 80.910 ;
        RECT 1814.800 80.590 1815.060 80.910 ;
        RECT 1814.860 24.210 1815.000 80.590 ;
        RECT 1814.860 24.070 1816.840 24.210 ;
        RECT 1816.700 2.400 1816.840 24.070 ;
        RECT 1816.490 -4.800 1817.050 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1065.430 1317.400 1065.750 1317.460 ;
        RECT 1817.990 1317.400 1818.310 1317.460 ;
        RECT 1065.430 1317.260 1818.310 1317.400 ;
        RECT 1065.430 1317.200 1065.750 1317.260 ;
        RECT 1817.990 1317.200 1818.310 1317.260 ;
        RECT 1817.990 20.640 1818.310 20.700 ;
        RECT 1834.550 20.640 1834.870 20.700 ;
        RECT 1817.990 20.500 1834.870 20.640 ;
        RECT 1817.990 20.440 1818.310 20.500 ;
        RECT 1834.550 20.440 1834.870 20.500 ;
      LAYER via ;
        RECT 1065.460 1317.200 1065.720 1317.460 ;
        RECT 1818.020 1317.200 1818.280 1317.460 ;
        RECT 1818.020 20.440 1818.280 20.700 ;
        RECT 1834.580 20.440 1834.840 20.700 ;
      LAYER met2 ;
        RECT 1065.500 1323.135 1065.780 1327.135 ;
        RECT 1065.520 1317.490 1065.660 1323.135 ;
        RECT 1065.460 1317.170 1065.720 1317.490 ;
        RECT 1818.020 1317.170 1818.280 1317.490 ;
        RECT 1818.080 20.730 1818.220 1317.170 ;
        RECT 1818.020 20.410 1818.280 20.730 ;
        RECT 1834.580 20.410 1834.840 20.730 ;
        RECT 1834.640 2.400 1834.780 20.410 ;
        RECT 1834.430 -4.800 1834.990 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1412.270 1317.060 1412.590 1317.120 ;
        RECT 1832.250 1317.060 1832.570 1317.120 ;
        RECT 1412.270 1316.920 1832.570 1317.060 ;
        RECT 1412.270 1316.860 1412.590 1316.920 ;
        RECT 1832.250 1316.860 1832.570 1316.920 ;
        RECT 1832.250 15.880 1832.570 15.940 ;
        RECT 1852.030 15.880 1852.350 15.940 ;
        RECT 1832.250 15.740 1852.350 15.880 ;
        RECT 1832.250 15.680 1832.570 15.740 ;
        RECT 1852.030 15.680 1852.350 15.740 ;
      LAYER via ;
        RECT 1412.300 1316.860 1412.560 1317.120 ;
        RECT 1832.280 1316.860 1832.540 1317.120 ;
        RECT 1832.280 15.680 1832.540 15.940 ;
        RECT 1852.060 15.680 1852.320 15.940 ;
      LAYER met2 ;
        RECT 1412.340 1323.135 1412.620 1327.135 ;
        RECT 1412.360 1317.150 1412.500 1323.135 ;
        RECT 1412.300 1316.830 1412.560 1317.150 ;
        RECT 1832.280 1316.830 1832.540 1317.150 ;
        RECT 1832.340 15.970 1832.480 1316.830 ;
        RECT 1832.280 15.650 1832.540 15.970 ;
        RECT 1852.060 15.650 1852.320 15.970 ;
        RECT 1852.120 2.400 1852.260 15.650 ;
        RECT 1851.910 -4.800 1852.470 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1505.190 1313.660 1505.510 1313.720 ;
        RECT 1831.790 1313.660 1832.110 1313.720 ;
        RECT 1505.190 1313.520 1832.110 1313.660 ;
        RECT 1505.190 1313.460 1505.510 1313.520 ;
        RECT 1831.790 1313.460 1832.110 1313.520 ;
        RECT 1831.790 19.960 1832.110 20.020 ;
        RECT 1869.970 19.960 1870.290 20.020 ;
        RECT 1831.790 19.820 1870.290 19.960 ;
        RECT 1831.790 19.760 1832.110 19.820 ;
        RECT 1869.970 19.760 1870.290 19.820 ;
      LAYER via ;
        RECT 1505.220 1313.460 1505.480 1313.720 ;
        RECT 1831.820 1313.460 1832.080 1313.720 ;
        RECT 1831.820 19.760 1832.080 20.020 ;
        RECT 1870.000 19.760 1870.260 20.020 ;
      LAYER met2 ;
        RECT 1505.260 1323.135 1505.540 1327.135 ;
        RECT 1505.280 1313.750 1505.420 1323.135 ;
        RECT 1505.220 1313.430 1505.480 1313.750 ;
        RECT 1831.820 1313.430 1832.080 1313.750 ;
        RECT 1831.880 20.050 1832.020 1313.430 ;
        RECT 1831.820 19.730 1832.080 20.050 ;
        RECT 1870.000 19.730 1870.260 20.050 ;
        RECT 1870.060 2.400 1870.200 19.730 ;
        RECT 1869.850 -4.800 1870.410 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 697.965 1368.925 698.135 1393.575 ;
        RECT 745.805 531.505 745.975 579.615 ;
        RECT 745.805 418.285 745.975 483.055 ;
        RECT 745.805 341.445 745.975 386.155 ;
        RECT 745.805 224.825 745.975 289.595 ;
        RECT 745.805 51.765 745.975 96.475 ;
      LAYER mcon ;
        RECT 697.965 1393.405 698.135 1393.575 ;
        RECT 745.805 579.445 745.975 579.615 ;
        RECT 745.805 482.885 745.975 483.055 ;
        RECT 745.805 385.985 745.975 386.155 ;
        RECT 745.805 289.425 745.975 289.595 ;
        RECT 745.805 96.305 745.975 96.475 ;
      LAYER met1 ;
        RECT 697.890 2391.800 698.210 2391.860 ;
        RECT 1224.590 2391.800 1224.910 2391.860 ;
        RECT 697.890 2391.660 1224.910 2391.800 ;
        RECT 697.890 2391.600 698.210 2391.660 ;
        RECT 1224.590 2391.600 1224.910 2391.660 ;
        RECT 697.890 1393.560 698.210 1393.620 ;
        RECT 697.890 1393.420 698.405 1393.560 ;
        RECT 697.890 1393.360 698.210 1393.420 ;
        RECT 697.890 1369.080 698.210 1369.140 ;
        RECT 697.695 1368.940 698.210 1369.080 ;
        RECT 697.890 1368.880 698.210 1368.940 ;
        RECT 697.890 1327.600 698.210 1327.660 ;
        RECT 697.890 1327.460 726.640 1327.600 ;
        RECT 697.890 1327.400 698.210 1327.460 ;
        RECT 726.500 1326.580 726.640 1327.460 ;
        RECT 745.730 1326.580 746.050 1326.640 ;
        RECT 726.500 1326.440 746.050 1326.580 ;
        RECT 745.730 1326.380 746.050 1326.440 ;
        RECT 745.730 676.160 746.050 676.220 ;
        RECT 746.650 676.160 746.970 676.220 ;
        RECT 745.730 676.020 746.970 676.160 ;
        RECT 745.730 675.960 746.050 676.020 ;
        RECT 746.650 675.960 746.970 676.020 ;
        RECT 745.730 579.600 746.050 579.660 ;
        RECT 745.535 579.460 746.050 579.600 ;
        RECT 745.730 579.400 746.050 579.460 ;
        RECT 745.730 531.660 746.050 531.720 ;
        RECT 745.535 531.520 746.050 531.660 ;
        RECT 745.730 531.460 746.050 531.520 ;
        RECT 745.730 483.040 746.050 483.100 ;
        RECT 745.535 482.900 746.050 483.040 ;
        RECT 745.730 482.840 746.050 482.900 ;
        RECT 745.730 418.440 746.050 418.500 ;
        RECT 745.535 418.300 746.050 418.440 ;
        RECT 745.730 418.240 746.050 418.300 ;
        RECT 745.730 386.140 746.050 386.200 ;
        RECT 745.535 386.000 746.050 386.140 ;
        RECT 745.730 385.940 746.050 386.000 ;
        RECT 745.730 341.600 746.050 341.660 ;
        RECT 745.535 341.460 746.050 341.600 ;
        RECT 745.730 341.400 746.050 341.460 ;
        RECT 745.730 289.580 746.050 289.640 ;
        RECT 745.535 289.440 746.050 289.580 ;
        RECT 745.730 289.380 746.050 289.440 ;
        RECT 745.730 224.980 746.050 225.040 ;
        RECT 745.535 224.840 746.050 224.980 ;
        RECT 745.730 224.780 746.050 224.840 ;
        RECT 745.730 96.460 746.050 96.520 ;
        RECT 745.535 96.320 746.050 96.460 ;
        RECT 745.730 96.260 746.050 96.320 ;
        RECT 745.730 51.920 746.050 51.980 ;
        RECT 745.535 51.780 746.050 51.920 ;
        RECT 745.730 51.720 746.050 51.780 ;
      LAYER via ;
        RECT 697.920 2391.600 698.180 2391.860 ;
        RECT 1224.620 2391.600 1224.880 2391.860 ;
        RECT 697.920 1393.360 698.180 1393.620 ;
        RECT 697.920 1368.880 698.180 1369.140 ;
        RECT 697.920 1327.400 698.180 1327.660 ;
        RECT 745.760 1326.380 746.020 1326.640 ;
        RECT 745.760 675.960 746.020 676.220 ;
        RECT 746.680 675.960 746.940 676.220 ;
        RECT 745.760 579.400 746.020 579.660 ;
        RECT 745.760 531.460 746.020 531.720 ;
        RECT 745.760 482.840 746.020 483.100 ;
        RECT 745.760 418.240 746.020 418.500 ;
        RECT 745.760 385.940 746.020 386.200 ;
        RECT 745.760 341.400 746.020 341.660 ;
        RECT 745.760 289.380 746.020 289.640 ;
        RECT 745.760 224.780 746.020 225.040 ;
        RECT 745.760 96.260 746.020 96.520 ;
        RECT 745.760 51.720 746.020 51.980 ;
      LAYER met2 ;
        RECT 697.920 2391.570 698.180 2391.890 ;
        RECT 1224.620 2391.570 1224.880 2391.890 ;
        RECT 697.980 1393.650 698.120 2391.570 ;
        RECT 1224.680 2377.880 1224.820 2391.570 ;
        RECT 1224.660 2373.880 1224.940 2377.880 ;
        RECT 697.920 1393.330 698.180 1393.650 ;
        RECT 697.920 1368.850 698.180 1369.170 ;
        RECT 697.980 1327.690 698.120 1368.850 ;
        RECT 697.920 1327.370 698.180 1327.690 ;
        RECT 745.760 1326.350 746.020 1326.670 ;
        RECT 745.820 870.245 745.960 1326.350 ;
        RECT 745.750 869.875 746.030 870.245 ;
        RECT 745.750 868.515 746.030 868.885 ;
        RECT 745.820 773.685 745.960 868.515 ;
        RECT 745.750 773.315 746.030 773.685 ;
        RECT 745.750 772.635 746.030 773.005 ;
        RECT 745.820 677.125 745.960 772.635 ;
        RECT 745.750 676.755 746.030 677.125 ;
        RECT 745.750 676.075 746.030 676.445 ;
        RECT 745.760 675.930 746.020 676.075 ;
        RECT 746.680 675.930 746.940 676.250 ;
        RECT 746.740 631.450 746.880 675.930 ;
        RECT 745.820 631.310 746.880 631.450 ;
        RECT 745.820 579.690 745.960 631.310 ;
        RECT 745.760 579.370 746.020 579.690 ;
        RECT 745.760 531.430 746.020 531.750 ;
        RECT 745.820 483.130 745.960 531.430 ;
        RECT 745.760 482.810 746.020 483.130 ;
        RECT 745.760 418.210 746.020 418.530 ;
        RECT 745.820 386.230 745.960 418.210 ;
        RECT 745.760 385.910 746.020 386.230 ;
        RECT 745.760 341.370 746.020 341.690 ;
        RECT 745.820 289.670 745.960 341.370 ;
        RECT 745.760 289.350 746.020 289.670 ;
        RECT 745.760 224.750 746.020 225.070 ;
        RECT 745.820 96.550 745.960 224.750 ;
        RECT 745.760 96.230 746.020 96.550 ;
        RECT 745.760 51.690 746.020 52.010 ;
        RECT 745.820 14.180 745.960 51.690 ;
        RECT 745.360 14.040 745.960 14.180 ;
        RECT 745.360 13.330 745.500 14.040 ;
        RECT 745.360 13.190 746.420 13.330 ;
        RECT 746.280 2.400 746.420 13.190 ;
        RECT 746.070 -4.800 746.630 2.400 ;
      LAYER via2 ;
        RECT 745.750 869.920 746.030 870.200 ;
        RECT 745.750 868.560 746.030 868.840 ;
        RECT 745.750 773.360 746.030 773.640 ;
        RECT 745.750 772.680 746.030 772.960 ;
        RECT 745.750 676.800 746.030 677.080 ;
        RECT 745.750 676.120 746.030 676.400 ;
      LAYER met3 ;
        RECT 745.725 870.210 746.055 870.225 ;
        RECT 745.510 869.895 746.055 870.210 ;
        RECT 745.510 868.865 745.810 869.895 ;
        RECT 745.510 868.550 746.055 868.865 ;
        RECT 745.725 868.535 746.055 868.550 ;
        RECT 745.725 773.650 746.055 773.665 ;
        RECT 745.510 773.335 746.055 773.650 ;
        RECT 745.510 772.985 745.810 773.335 ;
        RECT 745.510 772.670 746.055 772.985 ;
        RECT 745.725 772.655 746.055 772.670 ;
        RECT 745.725 677.090 746.055 677.105 ;
        RECT 745.510 676.775 746.055 677.090 ;
        RECT 745.510 676.425 745.810 676.775 ;
        RECT 745.510 676.110 746.055 676.425 ;
        RECT 745.725 676.095 746.055 676.110 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 717.210 1356.840 717.530 1356.900 ;
        RECT 719.510 1356.840 719.830 1356.900 ;
        RECT 717.210 1356.700 719.830 1356.840 ;
        RECT 717.210 1356.640 717.530 1356.700 ;
        RECT 719.510 1356.640 719.830 1356.700 ;
        RECT 1887.910 51.920 1888.230 51.980 ;
        RECT 746.280 51.780 1888.230 51.920 ;
        RECT 719.510 51.580 719.830 51.640 ;
        RECT 746.280 51.580 746.420 51.780 ;
        RECT 1887.910 51.720 1888.230 51.780 ;
        RECT 719.510 51.440 746.420 51.580 ;
        RECT 719.510 51.380 719.830 51.440 ;
      LAYER via ;
        RECT 717.240 1356.640 717.500 1356.900 ;
        RECT 719.540 1356.640 719.800 1356.900 ;
        RECT 719.540 51.380 719.800 51.640 ;
        RECT 1887.940 51.720 1888.200 51.980 ;
      LAYER met2 ;
        RECT 717.230 1366.955 717.510 1367.325 ;
        RECT 717.300 1356.930 717.440 1366.955 ;
        RECT 717.240 1356.610 717.500 1356.930 ;
        RECT 719.540 1356.610 719.800 1356.930 ;
        RECT 719.600 51.670 719.740 1356.610 ;
        RECT 1887.940 51.690 1888.200 52.010 ;
        RECT 719.540 51.350 719.800 51.670 ;
        RECT 1888.000 2.400 1888.140 51.690 ;
        RECT 1887.790 -4.800 1888.350 2.400 ;
      LAYER via2 ;
        RECT 717.230 1367.000 717.510 1367.280 ;
      LAYER met3 ;
        RECT 715.810 1369.415 719.810 1370.015 ;
        RECT 716.990 1367.305 717.290 1369.415 ;
        RECT 716.990 1366.990 717.535 1367.305 ;
        RECT 717.205 1366.975 717.535 1366.990 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1772.910 1842.700 1773.230 1842.760 ;
        RECT 1873.650 1842.700 1873.970 1842.760 ;
        RECT 1772.910 1842.560 1873.970 1842.700 ;
        RECT 1772.910 1842.500 1773.230 1842.560 ;
        RECT 1873.650 1842.500 1873.970 1842.560 ;
        RECT 1873.650 19.960 1873.970 20.020 ;
        RECT 1905.850 19.960 1906.170 20.020 ;
        RECT 1873.650 19.820 1906.170 19.960 ;
        RECT 1873.650 19.760 1873.970 19.820 ;
        RECT 1905.850 19.760 1906.170 19.820 ;
      LAYER via ;
        RECT 1772.940 1842.500 1773.200 1842.760 ;
        RECT 1873.680 1842.500 1873.940 1842.760 ;
        RECT 1873.680 19.760 1873.940 20.020 ;
        RECT 1905.880 19.760 1906.140 20.020 ;
      LAYER met2 ;
        RECT 1772.930 1844.315 1773.210 1844.685 ;
        RECT 1773.000 1842.790 1773.140 1844.315 ;
        RECT 1772.940 1842.470 1773.200 1842.790 ;
        RECT 1873.680 1842.470 1873.940 1842.790 ;
        RECT 1873.740 20.050 1873.880 1842.470 ;
        RECT 1873.680 19.730 1873.940 20.050 ;
        RECT 1905.880 19.730 1906.140 20.050 ;
        RECT 1905.940 2.400 1906.080 19.730 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
      LAYER via2 ;
        RECT 1772.930 1844.360 1773.210 1844.640 ;
      LAYER met3 ;
        RECT 1755.835 1844.650 1759.835 1844.655 ;
        RECT 1772.905 1844.650 1773.235 1844.665 ;
        RECT 1755.835 1844.350 1773.235 1844.650 ;
        RECT 1755.835 1844.055 1759.835 1844.350 ;
        RECT 1772.905 1844.335 1773.235 1844.350 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1603.630 1314.000 1603.950 1314.060 ;
        RECT 1907.690 1314.000 1908.010 1314.060 ;
        RECT 1603.630 1313.860 1908.010 1314.000 ;
        RECT 1603.630 1313.800 1603.950 1313.860 ;
        RECT 1907.690 1313.800 1908.010 1313.860 ;
        RECT 1907.690 20.300 1908.010 20.360 ;
        RECT 1923.330 20.300 1923.650 20.360 ;
        RECT 1907.690 20.160 1923.650 20.300 ;
        RECT 1907.690 20.100 1908.010 20.160 ;
        RECT 1923.330 20.100 1923.650 20.160 ;
      LAYER via ;
        RECT 1603.660 1313.800 1603.920 1314.060 ;
        RECT 1907.720 1313.800 1907.980 1314.060 ;
        RECT 1907.720 20.100 1907.980 20.360 ;
        RECT 1923.360 20.100 1923.620 20.360 ;
      LAYER met2 ;
        RECT 1603.700 1323.135 1603.980 1327.135 ;
        RECT 1603.720 1314.090 1603.860 1323.135 ;
        RECT 1603.660 1313.770 1603.920 1314.090 ;
        RECT 1907.720 1313.770 1907.980 1314.090 ;
        RECT 1907.780 20.390 1907.920 1313.770 ;
        RECT 1907.720 20.070 1907.980 20.390 ;
        RECT 1923.360 20.070 1923.620 20.390 ;
        RECT 1923.420 2.400 1923.560 20.070 ;
        RECT 1923.210 -4.800 1923.770 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1772.450 1338.820 1772.770 1338.880 ;
        RECT 1915.050 1338.820 1915.370 1338.880 ;
        RECT 1772.450 1338.680 1915.370 1338.820 ;
        RECT 1772.450 1338.620 1772.770 1338.680 ;
        RECT 1915.050 1338.620 1915.370 1338.680 ;
        RECT 1915.050 19.960 1915.370 20.020 ;
        RECT 1941.270 19.960 1941.590 20.020 ;
        RECT 1915.050 19.820 1941.590 19.960 ;
        RECT 1915.050 19.760 1915.370 19.820 ;
        RECT 1941.270 19.760 1941.590 19.820 ;
      LAYER via ;
        RECT 1772.480 1338.620 1772.740 1338.880 ;
        RECT 1915.080 1338.620 1915.340 1338.880 ;
        RECT 1915.080 19.760 1915.340 20.020 ;
        RECT 1941.300 19.760 1941.560 20.020 ;
      LAYER met2 ;
        RECT 1772.470 1339.755 1772.750 1340.125 ;
        RECT 1772.540 1338.910 1772.680 1339.755 ;
        RECT 1772.480 1338.590 1772.740 1338.910 ;
        RECT 1915.080 1338.590 1915.340 1338.910 ;
        RECT 1915.140 20.050 1915.280 1338.590 ;
        RECT 1915.080 19.730 1915.340 20.050 ;
        RECT 1941.300 19.730 1941.560 20.050 ;
        RECT 1941.360 2.400 1941.500 19.730 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
      LAYER via2 ;
        RECT 1772.470 1339.800 1772.750 1340.080 ;
      LAYER met3 ;
        RECT 1755.835 1340.090 1759.835 1340.095 ;
        RECT 1772.445 1340.090 1772.775 1340.105 ;
        RECT 1755.835 1339.790 1772.775 1340.090 ;
        RECT 1755.835 1339.495 1759.835 1339.790 ;
        RECT 1772.445 1339.775 1772.775 1339.790 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1667.110 1312.980 1667.430 1313.040 ;
        RECT 1921.490 1312.980 1921.810 1313.040 ;
        RECT 1667.110 1312.840 1921.810 1312.980 ;
        RECT 1667.110 1312.780 1667.430 1312.840 ;
        RECT 1921.490 1312.780 1921.810 1312.840 ;
        RECT 1921.490 16.560 1921.810 16.620 ;
        RECT 1959.210 16.560 1959.530 16.620 ;
        RECT 1921.490 16.420 1959.530 16.560 ;
        RECT 1921.490 16.360 1921.810 16.420 ;
        RECT 1959.210 16.360 1959.530 16.420 ;
      LAYER via ;
        RECT 1667.140 1312.780 1667.400 1313.040 ;
        RECT 1921.520 1312.780 1921.780 1313.040 ;
        RECT 1921.520 16.360 1921.780 16.620 ;
        RECT 1959.240 16.360 1959.500 16.620 ;
      LAYER met2 ;
        RECT 1667.180 1323.135 1667.460 1327.135 ;
        RECT 1667.200 1313.070 1667.340 1323.135 ;
        RECT 1667.140 1312.750 1667.400 1313.070 ;
        RECT 1921.520 1312.750 1921.780 1313.070 ;
        RECT 1921.580 16.650 1921.720 1312.750 ;
        RECT 1921.520 16.330 1921.780 16.650 ;
        RECT 1959.240 16.330 1959.500 16.650 ;
        RECT 1959.300 2.400 1959.440 16.330 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1074.650 2378.115 1074.930 2378.485 ;
        RECT 1758.670 2378.115 1758.950 2378.485 ;
        RECT 1074.720 2377.880 1074.860 2378.115 ;
        RECT 1074.700 2373.880 1074.980 2377.880 ;
        RECT 1758.740 2360.125 1758.880 2378.115 ;
        RECT 1758.670 2359.755 1758.950 2360.125 ;
        RECT 1777.530 1669.555 1777.810 1669.925 ;
        RECT 1777.600 1581.525 1777.740 1669.555 ;
        RECT 1777.530 1581.155 1777.810 1581.525 ;
        RECT 1779.830 1386.675 1780.110 1387.045 ;
        RECT 1779.900 1353.725 1780.040 1386.675 ;
        RECT 1779.830 1353.355 1780.110 1353.725 ;
        RECT 1778.910 1227.555 1779.190 1227.925 ;
        RECT 1778.980 1204.125 1779.120 1227.555 ;
        RECT 1778.910 1203.755 1779.190 1204.125 ;
        RECT 1777.070 1152.075 1777.350 1152.445 ;
        RECT 1777.140 1104.845 1777.280 1152.075 ;
        RECT 1777.070 1104.475 1777.350 1104.845 ;
        RECT 1778.450 1048.035 1778.730 1048.405 ;
        RECT 1778.520 1000.805 1778.660 1048.035 ;
        RECT 1778.450 1000.435 1778.730 1000.805 ;
        RECT 1776.150 999.755 1776.430 1000.125 ;
        RECT 1776.220 952.525 1776.360 999.755 ;
        RECT 1776.150 952.155 1776.430 952.525 ;
        RECT 1777.070 950.795 1777.350 951.165 ;
        RECT 1777.140 904.245 1777.280 950.795 ;
        RECT 1777.070 903.875 1777.350 904.245 ;
        RECT 1777.990 613.515 1778.270 613.885 ;
        RECT 1778.060 566.965 1778.200 613.515 ;
        RECT 1777.990 566.595 1778.270 566.965 ;
        RECT 1777.990 516.275 1778.270 516.645 ;
        RECT 1778.060 428.925 1778.200 516.275 ;
        RECT 1777.990 428.555 1778.270 428.925 ;
        RECT 1779.830 396.595 1780.110 396.965 ;
        RECT 1779.900 373.845 1780.040 396.595 ;
        RECT 1779.830 373.475 1780.110 373.845 ;
        RECT 1779.830 372.115 1780.110 372.485 ;
        RECT 1779.900 325.565 1780.040 372.115 ;
        RECT 1779.830 325.195 1780.110 325.565 ;
        RECT 1779.830 304.115 1780.110 304.485 ;
        RECT 1779.900 282.725 1780.040 304.115 ;
        RECT 1779.830 282.355 1780.110 282.725 ;
        RECT 1777.990 88.555 1778.270 88.925 ;
        RECT 1778.060 47.445 1778.200 88.555 ;
        RECT 1777.990 47.075 1778.270 47.445 ;
        RECT 1977.170 15.795 1977.450 16.165 ;
        RECT 1977.240 2.400 1977.380 15.795 ;
        RECT 1977.030 -4.800 1977.590 2.400 ;
      LAYER via2 ;
        RECT 1074.650 2378.160 1074.930 2378.440 ;
        RECT 1758.670 2378.160 1758.950 2378.440 ;
        RECT 1758.670 2359.800 1758.950 2360.080 ;
        RECT 1777.530 1669.600 1777.810 1669.880 ;
        RECT 1777.530 1581.200 1777.810 1581.480 ;
        RECT 1779.830 1386.720 1780.110 1387.000 ;
        RECT 1779.830 1353.400 1780.110 1353.680 ;
        RECT 1778.910 1227.600 1779.190 1227.880 ;
        RECT 1778.910 1203.800 1779.190 1204.080 ;
        RECT 1777.070 1152.120 1777.350 1152.400 ;
        RECT 1777.070 1104.520 1777.350 1104.800 ;
        RECT 1778.450 1048.080 1778.730 1048.360 ;
        RECT 1778.450 1000.480 1778.730 1000.760 ;
        RECT 1776.150 999.800 1776.430 1000.080 ;
        RECT 1776.150 952.200 1776.430 952.480 ;
        RECT 1777.070 950.840 1777.350 951.120 ;
        RECT 1777.070 903.920 1777.350 904.200 ;
        RECT 1777.990 613.560 1778.270 613.840 ;
        RECT 1777.990 566.640 1778.270 566.920 ;
        RECT 1777.990 516.320 1778.270 516.600 ;
        RECT 1777.990 428.600 1778.270 428.880 ;
        RECT 1779.830 396.640 1780.110 396.920 ;
        RECT 1779.830 373.520 1780.110 373.800 ;
        RECT 1779.830 372.160 1780.110 372.440 ;
        RECT 1779.830 325.240 1780.110 325.520 ;
        RECT 1779.830 304.160 1780.110 304.440 ;
        RECT 1779.830 282.400 1780.110 282.680 ;
        RECT 1777.990 88.600 1778.270 88.880 ;
        RECT 1777.990 47.120 1778.270 47.400 ;
        RECT 1977.170 15.840 1977.450 16.120 ;
      LAYER met3 ;
        RECT 1074.625 2378.450 1074.955 2378.465 ;
        RECT 1758.645 2378.450 1758.975 2378.465 ;
        RECT 1074.625 2378.150 1758.975 2378.450 ;
        RECT 1074.625 2378.135 1074.955 2378.150 ;
        RECT 1758.645 2378.135 1758.975 2378.150 ;
        RECT 1758.645 2360.090 1758.975 2360.105 ;
        RECT 1774.950 2360.090 1775.330 2360.100 ;
        RECT 1758.645 2359.790 1775.330 2360.090 ;
        RECT 1758.645 2359.775 1758.975 2359.790 ;
        RECT 1774.950 2359.780 1775.330 2359.790 ;
        RECT 1774.950 2309.770 1775.330 2309.780 ;
        RECT 1777.710 2309.770 1778.090 2309.780 ;
        RECT 1774.950 2309.470 1778.090 2309.770 ;
        RECT 1774.950 2309.460 1775.330 2309.470 ;
        RECT 1777.710 2309.460 1778.090 2309.470 ;
        RECT 1777.710 2223.410 1778.090 2223.420 ;
        RECT 1775.910 2223.110 1778.090 2223.410 ;
        RECT 1775.910 2221.380 1776.210 2223.110 ;
        RECT 1777.710 2223.100 1778.090 2223.110 ;
        RECT 1775.870 2221.060 1776.250 2221.380 ;
        RECT 1775.870 2125.490 1776.250 2125.500 ;
        RECT 1777.710 2125.490 1778.090 2125.500 ;
        RECT 1775.870 2125.190 1778.090 2125.490 ;
        RECT 1775.870 2125.180 1776.250 2125.190 ;
        RECT 1777.710 2125.180 1778.090 2125.190 ;
        RECT 1775.870 2001.730 1776.250 2001.740 ;
        RECT 1777.710 2001.730 1778.090 2001.740 ;
        RECT 1775.870 2001.430 1778.090 2001.730 ;
        RECT 1775.870 2001.420 1776.250 2001.430 ;
        RECT 1777.710 2001.420 1778.090 2001.430 ;
        RECT 1775.870 1949.370 1776.250 1949.380 ;
        RECT 1777.710 1949.370 1778.090 1949.380 ;
        RECT 1775.870 1949.070 1778.090 1949.370 ;
        RECT 1775.870 1949.060 1776.250 1949.070 ;
        RECT 1777.710 1949.060 1778.090 1949.070 ;
        RECT 1774.950 1859.610 1775.330 1859.620 ;
        RECT 1777.710 1859.610 1778.090 1859.620 ;
        RECT 1774.950 1859.310 1778.090 1859.610 ;
        RECT 1774.950 1859.300 1775.330 1859.310 ;
        RECT 1777.710 1859.300 1778.090 1859.310 ;
        RECT 1775.870 1724.660 1776.250 1724.980 ;
        RECT 1774.950 1724.290 1775.330 1724.300 ;
        RECT 1775.910 1724.290 1776.210 1724.660 ;
        RECT 1774.950 1723.990 1776.210 1724.290 ;
        RECT 1774.950 1723.980 1775.330 1723.990 ;
        RECT 1775.870 1669.890 1776.250 1669.900 ;
        RECT 1777.505 1669.890 1777.835 1669.905 ;
        RECT 1775.870 1669.590 1777.835 1669.890 ;
        RECT 1775.870 1669.580 1776.250 1669.590 ;
        RECT 1777.505 1669.575 1777.835 1669.590 ;
        RECT 1777.505 1581.490 1777.835 1581.505 ;
        RECT 1774.990 1581.190 1777.835 1581.490 ;
        RECT 1774.990 1580.820 1775.290 1581.190 ;
        RECT 1777.505 1581.175 1777.835 1581.190 ;
        RECT 1774.950 1580.500 1775.330 1580.820 ;
        RECT 1774.950 1473.370 1775.330 1473.380 ;
        RECT 1777.710 1473.370 1778.090 1473.380 ;
        RECT 1774.950 1473.070 1778.090 1473.370 ;
        RECT 1774.950 1473.060 1775.330 1473.070 ;
        RECT 1777.710 1473.060 1778.090 1473.070 ;
        RECT 1777.710 1387.010 1778.090 1387.020 ;
        RECT 1779.805 1387.010 1780.135 1387.025 ;
        RECT 1777.710 1386.710 1780.135 1387.010 ;
        RECT 1777.710 1386.700 1778.090 1386.710 ;
        RECT 1779.805 1386.695 1780.135 1386.710 ;
        RECT 1777.710 1353.690 1778.090 1353.700 ;
        RECT 1779.805 1353.690 1780.135 1353.705 ;
        RECT 1777.710 1353.390 1780.135 1353.690 ;
        RECT 1777.710 1353.380 1778.090 1353.390 ;
        RECT 1779.805 1353.375 1780.135 1353.390 ;
        RECT 1778.885 1227.900 1779.215 1227.905 ;
        RECT 1778.630 1227.890 1779.215 1227.900 ;
        RECT 1778.630 1227.590 1779.440 1227.890 ;
        RECT 1778.630 1227.580 1779.215 1227.590 ;
        RECT 1778.885 1227.575 1779.215 1227.580 ;
        RECT 1778.885 1204.100 1779.215 1204.105 ;
        RECT 1778.630 1204.090 1779.215 1204.100 ;
        RECT 1778.430 1203.790 1779.215 1204.090 ;
        RECT 1778.630 1203.780 1779.215 1203.790 ;
        RECT 1778.885 1203.775 1779.215 1203.780 ;
        RECT 1777.045 1152.410 1777.375 1152.425 ;
        RECT 1778.630 1152.410 1779.010 1152.420 ;
        RECT 1777.045 1152.110 1779.010 1152.410 ;
        RECT 1777.045 1152.095 1777.375 1152.110 ;
        RECT 1778.630 1152.100 1779.010 1152.110 ;
        RECT 1777.045 1104.810 1777.375 1104.825 ;
        RECT 1777.710 1104.810 1778.090 1104.820 ;
        RECT 1777.045 1104.510 1778.090 1104.810 ;
        RECT 1777.045 1104.495 1777.375 1104.510 ;
        RECT 1777.710 1104.500 1778.090 1104.510 ;
        RECT 1778.630 1049.730 1779.010 1049.740 ;
        RECT 1777.750 1049.430 1779.010 1049.730 ;
        RECT 1777.750 1049.060 1778.050 1049.430 ;
        RECT 1778.630 1049.420 1779.010 1049.430 ;
        RECT 1777.710 1048.740 1778.090 1049.060 ;
        RECT 1777.710 1048.370 1778.090 1048.380 ;
        RECT 1778.425 1048.370 1778.755 1048.385 ;
        RECT 1777.710 1048.070 1778.755 1048.370 ;
        RECT 1777.710 1048.060 1778.090 1048.070 ;
        RECT 1778.425 1048.055 1778.755 1048.070 ;
        RECT 1777.710 1000.770 1778.090 1000.780 ;
        RECT 1778.425 1000.770 1778.755 1000.785 ;
        RECT 1777.710 1000.470 1778.755 1000.770 ;
        RECT 1777.710 1000.460 1778.090 1000.470 ;
        RECT 1778.425 1000.455 1778.755 1000.470 ;
        RECT 1776.125 1000.090 1776.455 1000.105 ;
        RECT 1777.710 1000.090 1778.090 1000.100 ;
        RECT 1776.125 999.790 1778.090 1000.090 ;
        RECT 1776.125 999.775 1776.455 999.790 ;
        RECT 1777.710 999.780 1778.090 999.790 ;
        RECT 1776.125 952.500 1776.455 952.505 ;
        RECT 1775.870 952.490 1776.455 952.500 ;
        RECT 1775.670 952.190 1776.455 952.490 ;
        RECT 1775.870 952.180 1776.455 952.190 ;
        RECT 1776.125 952.175 1776.455 952.180 ;
        RECT 1775.870 951.500 1776.250 951.820 ;
        RECT 1775.910 951.130 1776.210 951.500 ;
        RECT 1777.045 951.130 1777.375 951.145 ;
        RECT 1775.910 950.830 1777.375 951.130 ;
        RECT 1777.045 950.815 1777.375 950.830 ;
        RECT 1777.045 904.210 1777.375 904.225 ;
        RECT 1777.710 904.210 1778.090 904.220 ;
        RECT 1777.045 903.910 1778.090 904.210 ;
        RECT 1777.045 903.895 1777.375 903.910 ;
        RECT 1777.710 903.900 1778.090 903.910 ;
        RECT 1778.630 883.810 1779.010 883.820 ;
        RECT 1777.750 883.510 1779.010 883.810 ;
        RECT 1777.750 883.140 1778.050 883.510 ;
        RECT 1778.630 883.500 1779.010 883.510 ;
        RECT 1777.710 882.820 1778.090 883.140 ;
        RECT 1777.710 772.660 1778.090 772.980 ;
        RECT 1777.750 772.290 1778.050 772.660 ;
        RECT 1778.630 772.290 1779.010 772.300 ;
        RECT 1777.750 771.990 1779.010 772.290 ;
        RECT 1778.630 771.980 1779.010 771.990 ;
        RECT 1777.710 690.380 1778.090 690.700 ;
        RECT 1777.750 689.330 1778.050 690.380 ;
        RECT 1778.630 689.330 1779.010 689.340 ;
        RECT 1777.750 689.030 1779.010 689.330 ;
        RECT 1778.630 689.020 1779.010 689.030 ;
        RECT 1777.710 628.130 1778.090 628.140 ;
        RECT 1778.630 628.130 1779.010 628.140 ;
        RECT 1777.710 627.830 1779.010 628.130 ;
        RECT 1777.710 627.820 1778.090 627.830 ;
        RECT 1778.630 627.820 1779.010 627.830 ;
        RECT 1777.965 613.860 1778.295 613.865 ;
        RECT 1777.710 613.850 1778.295 613.860 ;
        RECT 1777.710 613.550 1778.520 613.850 ;
        RECT 1777.710 613.540 1778.295 613.550 ;
        RECT 1777.965 613.535 1778.295 613.540 ;
        RECT 1777.965 566.930 1778.295 566.945 ;
        RECT 1777.750 566.615 1778.295 566.930 ;
        RECT 1777.750 566.260 1778.050 566.615 ;
        RECT 1777.710 565.940 1778.090 566.260 ;
        RECT 1777.710 516.980 1778.090 517.300 ;
        RECT 1777.750 516.625 1778.050 516.980 ;
        RECT 1777.750 516.310 1778.295 516.625 ;
        RECT 1777.965 516.295 1778.295 516.310 ;
        RECT 1777.965 428.890 1778.295 428.905 ;
        RECT 1778.630 428.890 1779.010 428.900 ;
        RECT 1777.965 428.590 1779.010 428.890 ;
        RECT 1777.965 428.575 1778.295 428.590 ;
        RECT 1778.630 428.580 1779.010 428.590 ;
        RECT 1778.630 427.530 1779.010 427.540 ;
        RECT 1777.750 427.230 1779.010 427.530 ;
        RECT 1777.750 426.860 1778.050 427.230 ;
        RECT 1778.630 427.220 1779.010 427.230 ;
        RECT 1777.710 426.540 1778.090 426.860 ;
        RECT 1777.710 396.930 1778.090 396.940 ;
        RECT 1779.805 396.930 1780.135 396.945 ;
        RECT 1777.710 396.630 1780.135 396.930 ;
        RECT 1777.710 396.620 1778.090 396.630 ;
        RECT 1779.805 396.615 1780.135 396.630 ;
        RECT 1779.805 373.820 1780.135 373.825 ;
        RECT 1779.550 373.810 1780.135 373.820 ;
        RECT 1779.550 373.510 1780.360 373.810 ;
        RECT 1779.550 373.500 1780.135 373.510 ;
        RECT 1779.805 373.495 1780.135 373.500 ;
        RECT 1779.805 372.460 1780.135 372.465 ;
        RECT 1779.550 372.450 1780.135 372.460 ;
        RECT 1779.550 372.150 1780.360 372.450 ;
        RECT 1779.550 372.140 1780.135 372.150 ;
        RECT 1779.805 372.135 1780.135 372.140 ;
        RECT 1779.805 325.530 1780.135 325.545 ;
        RECT 1779.590 325.215 1780.135 325.530 ;
        RECT 1779.590 324.860 1779.890 325.215 ;
        RECT 1779.550 324.540 1779.930 324.860 ;
        RECT 1779.805 304.460 1780.135 304.465 ;
        RECT 1779.550 304.450 1780.135 304.460 ;
        RECT 1779.550 304.150 1780.360 304.450 ;
        RECT 1779.550 304.140 1780.135 304.150 ;
        RECT 1779.805 304.135 1780.135 304.140 ;
        RECT 1779.805 282.700 1780.135 282.705 ;
        RECT 1779.550 282.690 1780.135 282.700 ;
        RECT 1779.350 282.390 1780.135 282.690 ;
        RECT 1779.550 282.380 1780.135 282.390 ;
        RECT 1779.805 282.375 1780.135 282.380 ;
        RECT 1779.550 234.100 1779.930 234.420 ;
        RECT 1777.710 233.050 1778.090 233.060 ;
        RECT 1779.590 233.050 1779.890 234.100 ;
        RECT 1777.710 232.750 1779.890 233.050 ;
        RECT 1777.710 232.740 1778.090 232.750 ;
        RECT 1777.710 89.260 1778.090 89.580 ;
        RECT 1777.750 88.905 1778.050 89.260 ;
        RECT 1777.750 88.590 1778.295 88.905 ;
        RECT 1777.965 88.575 1778.295 88.590 ;
        RECT 1777.965 47.410 1778.295 47.425 ;
        RECT 1778.630 47.410 1779.010 47.420 ;
        RECT 1777.965 47.110 1779.010 47.410 ;
        RECT 1777.965 47.095 1778.295 47.110 ;
        RECT 1778.630 47.100 1779.010 47.110 ;
        RECT 1778.630 16.130 1779.010 16.140 ;
        RECT 1977.145 16.130 1977.475 16.145 ;
        RECT 1778.630 15.830 1977.475 16.130 ;
        RECT 1778.630 15.820 1779.010 15.830 ;
        RECT 1977.145 15.815 1977.475 15.830 ;
      LAYER via3 ;
        RECT 1774.980 2359.780 1775.300 2360.100 ;
        RECT 1774.980 2309.460 1775.300 2309.780 ;
        RECT 1777.740 2309.460 1778.060 2309.780 ;
        RECT 1777.740 2223.100 1778.060 2223.420 ;
        RECT 1775.900 2221.060 1776.220 2221.380 ;
        RECT 1775.900 2125.180 1776.220 2125.500 ;
        RECT 1777.740 2125.180 1778.060 2125.500 ;
        RECT 1775.900 2001.420 1776.220 2001.740 ;
        RECT 1777.740 2001.420 1778.060 2001.740 ;
        RECT 1775.900 1949.060 1776.220 1949.380 ;
        RECT 1777.740 1949.060 1778.060 1949.380 ;
        RECT 1774.980 1859.300 1775.300 1859.620 ;
        RECT 1777.740 1859.300 1778.060 1859.620 ;
        RECT 1775.900 1724.660 1776.220 1724.980 ;
        RECT 1774.980 1723.980 1775.300 1724.300 ;
        RECT 1775.900 1669.580 1776.220 1669.900 ;
        RECT 1774.980 1580.500 1775.300 1580.820 ;
        RECT 1774.980 1473.060 1775.300 1473.380 ;
        RECT 1777.740 1473.060 1778.060 1473.380 ;
        RECT 1777.740 1386.700 1778.060 1387.020 ;
        RECT 1777.740 1353.380 1778.060 1353.700 ;
        RECT 1778.660 1227.580 1778.980 1227.900 ;
        RECT 1778.660 1203.780 1778.980 1204.100 ;
        RECT 1778.660 1152.100 1778.980 1152.420 ;
        RECT 1777.740 1104.500 1778.060 1104.820 ;
        RECT 1778.660 1049.420 1778.980 1049.740 ;
        RECT 1777.740 1048.740 1778.060 1049.060 ;
        RECT 1777.740 1048.060 1778.060 1048.380 ;
        RECT 1777.740 1000.460 1778.060 1000.780 ;
        RECT 1777.740 999.780 1778.060 1000.100 ;
        RECT 1775.900 952.180 1776.220 952.500 ;
        RECT 1775.900 951.500 1776.220 951.820 ;
        RECT 1777.740 903.900 1778.060 904.220 ;
        RECT 1778.660 883.500 1778.980 883.820 ;
        RECT 1777.740 882.820 1778.060 883.140 ;
        RECT 1777.740 772.660 1778.060 772.980 ;
        RECT 1778.660 771.980 1778.980 772.300 ;
        RECT 1777.740 690.380 1778.060 690.700 ;
        RECT 1778.660 689.020 1778.980 689.340 ;
        RECT 1777.740 627.820 1778.060 628.140 ;
        RECT 1778.660 627.820 1778.980 628.140 ;
        RECT 1777.740 613.540 1778.060 613.860 ;
        RECT 1777.740 565.940 1778.060 566.260 ;
        RECT 1777.740 516.980 1778.060 517.300 ;
        RECT 1778.660 428.580 1778.980 428.900 ;
        RECT 1778.660 427.220 1778.980 427.540 ;
        RECT 1777.740 426.540 1778.060 426.860 ;
        RECT 1777.740 396.620 1778.060 396.940 ;
        RECT 1779.580 373.500 1779.900 373.820 ;
        RECT 1779.580 372.140 1779.900 372.460 ;
        RECT 1779.580 324.540 1779.900 324.860 ;
        RECT 1779.580 304.140 1779.900 304.460 ;
        RECT 1779.580 282.380 1779.900 282.700 ;
        RECT 1779.580 234.100 1779.900 234.420 ;
        RECT 1777.740 232.740 1778.060 233.060 ;
        RECT 1777.740 89.260 1778.060 89.580 ;
        RECT 1778.660 47.100 1778.980 47.420 ;
        RECT 1778.660 15.820 1778.980 16.140 ;
      LAYER met4 ;
        RECT 1774.975 2359.775 1775.305 2360.105 ;
        RECT 1774.990 2309.785 1775.290 2359.775 ;
        RECT 1774.975 2309.455 1775.305 2309.785 ;
        RECT 1777.735 2309.455 1778.065 2309.785 ;
        RECT 1777.750 2223.425 1778.050 2309.455 ;
        RECT 1777.735 2223.095 1778.065 2223.425 ;
        RECT 1775.895 2221.055 1776.225 2221.385 ;
        RECT 1775.910 2125.505 1776.210 2221.055 ;
        RECT 1775.895 2125.175 1776.225 2125.505 ;
        RECT 1777.735 2125.175 1778.065 2125.505 ;
        RECT 1777.750 2001.745 1778.050 2125.175 ;
        RECT 1775.895 2001.415 1776.225 2001.745 ;
        RECT 1777.735 2001.415 1778.065 2001.745 ;
        RECT 1775.910 1949.385 1776.210 2001.415 ;
        RECT 1775.895 1949.055 1776.225 1949.385 ;
        RECT 1777.735 1949.055 1778.065 1949.385 ;
        RECT 1777.750 1859.625 1778.050 1949.055 ;
        RECT 1774.975 1859.295 1775.305 1859.625 ;
        RECT 1777.735 1859.295 1778.065 1859.625 ;
        RECT 1774.990 1763.050 1775.290 1859.295 ;
        RECT 1774.990 1762.750 1776.210 1763.050 ;
        RECT 1775.910 1724.985 1776.210 1762.750 ;
        RECT 1775.895 1724.655 1776.225 1724.985 ;
        RECT 1774.975 1723.975 1775.305 1724.305 ;
        RECT 1774.990 1678.050 1775.290 1723.975 ;
        RECT 1774.990 1677.750 1776.210 1678.050 ;
        RECT 1775.910 1669.905 1776.210 1677.750 ;
        RECT 1775.895 1669.575 1776.225 1669.905 ;
        RECT 1774.975 1580.495 1775.305 1580.825 ;
        RECT 1774.990 1473.385 1775.290 1580.495 ;
        RECT 1774.975 1473.055 1775.305 1473.385 ;
        RECT 1777.735 1473.055 1778.065 1473.385 ;
        RECT 1777.750 1387.025 1778.050 1473.055 ;
        RECT 1777.735 1386.695 1778.065 1387.025 ;
        RECT 1777.735 1353.375 1778.065 1353.705 ;
        RECT 1777.750 1283.650 1778.050 1353.375 ;
        RECT 1777.750 1283.350 1778.970 1283.650 ;
        RECT 1778.670 1227.905 1778.970 1283.350 ;
        RECT 1778.655 1227.575 1778.985 1227.905 ;
        RECT 1778.655 1203.775 1778.985 1204.105 ;
        RECT 1778.670 1152.425 1778.970 1203.775 ;
        RECT 1778.655 1152.095 1778.985 1152.425 ;
        RECT 1777.735 1104.495 1778.065 1104.825 ;
        RECT 1777.750 1096.650 1778.050 1104.495 ;
        RECT 1777.750 1096.350 1778.970 1096.650 ;
        RECT 1778.670 1049.745 1778.970 1096.350 ;
        RECT 1778.655 1049.415 1778.985 1049.745 ;
        RECT 1777.735 1048.735 1778.065 1049.065 ;
        RECT 1777.750 1048.385 1778.050 1048.735 ;
        RECT 1777.735 1048.055 1778.065 1048.385 ;
        RECT 1777.735 1000.455 1778.065 1000.785 ;
        RECT 1777.750 1000.105 1778.050 1000.455 ;
        RECT 1777.735 999.775 1778.065 1000.105 ;
        RECT 1775.895 952.175 1776.225 952.505 ;
        RECT 1775.910 951.825 1776.210 952.175 ;
        RECT 1775.895 951.495 1776.225 951.825 ;
        RECT 1777.735 903.895 1778.065 904.225 ;
        RECT 1777.750 902.850 1778.050 903.895 ;
        RECT 1777.750 902.550 1778.970 902.850 ;
        RECT 1778.670 883.825 1778.970 902.550 ;
        RECT 1778.655 883.495 1778.985 883.825 ;
        RECT 1777.735 882.815 1778.065 883.145 ;
        RECT 1777.750 772.985 1778.050 882.815 ;
        RECT 1777.735 772.655 1778.065 772.985 ;
        RECT 1778.655 771.975 1778.985 772.305 ;
        RECT 1778.670 736.250 1778.970 771.975 ;
        RECT 1777.750 735.950 1778.970 736.250 ;
        RECT 1777.750 690.705 1778.050 735.950 ;
        RECT 1777.735 690.375 1778.065 690.705 ;
        RECT 1778.655 689.015 1778.985 689.345 ;
        RECT 1778.670 628.145 1778.970 689.015 ;
        RECT 1777.735 627.815 1778.065 628.145 ;
        RECT 1778.655 627.815 1778.985 628.145 ;
        RECT 1777.750 613.865 1778.050 627.815 ;
        RECT 1777.735 613.535 1778.065 613.865 ;
        RECT 1777.735 565.935 1778.065 566.265 ;
        RECT 1777.750 517.305 1778.050 565.935 ;
        RECT 1777.735 516.975 1778.065 517.305 ;
        RECT 1778.655 428.575 1778.985 428.905 ;
        RECT 1778.670 427.545 1778.970 428.575 ;
        RECT 1778.655 427.215 1778.985 427.545 ;
        RECT 1777.735 426.535 1778.065 426.865 ;
        RECT 1777.750 396.945 1778.050 426.535 ;
        RECT 1777.735 396.615 1778.065 396.945 ;
        RECT 1779.575 373.495 1779.905 373.825 ;
        RECT 1779.590 372.465 1779.890 373.495 ;
        RECT 1779.575 372.135 1779.905 372.465 ;
        RECT 1779.575 324.535 1779.905 324.865 ;
        RECT 1779.590 304.465 1779.890 324.535 ;
        RECT 1779.575 304.135 1779.905 304.465 ;
        RECT 1779.575 282.375 1779.905 282.705 ;
        RECT 1779.590 234.425 1779.890 282.375 ;
        RECT 1779.575 234.095 1779.905 234.425 ;
        RECT 1777.735 232.735 1778.065 233.065 ;
        RECT 1777.750 89.585 1778.050 232.735 ;
        RECT 1777.735 89.255 1778.065 89.585 ;
        RECT 1778.655 47.095 1778.985 47.425 ;
        RECT 1778.670 16.145 1778.970 47.095 ;
        RECT 1778.655 15.815 1778.985 16.145 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1699.310 2392.480 1699.630 2392.540 ;
        RECT 1976.690 2392.480 1977.010 2392.540 ;
        RECT 1699.310 2392.340 1977.010 2392.480 ;
        RECT 1699.310 2392.280 1699.630 2392.340 ;
        RECT 1976.690 2392.280 1977.010 2392.340 ;
        RECT 1976.690 19.620 1977.010 19.680 ;
        RECT 1995.090 19.620 1995.410 19.680 ;
        RECT 1976.690 19.480 1995.410 19.620 ;
        RECT 1976.690 19.420 1977.010 19.480 ;
        RECT 1995.090 19.420 1995.410 19.480 ;
      LAYER via ;
        RECT 1699.340 2392.280 1699.600 2392.540 ;
        RECT 1976.720 2392.280 1976.980 2392.540 ;
        RECT 1976.720 19.420 1976.980 19.680 ;
        RECT 1995.120 19.420 1995.380 19.680 ;
      LAYER met2 ;
        RECT 1699.340 2392.250 1699.600 2392.570 ;
        RECT 1976.720 2392.250 1976.980 2392.570 ;
        RECT 1699.400 2377.880 1699.540 2392.250 ;
        RECT 1699.380 2373.880 1699.660 2377.880 ;
        RECT 1976.780 19.710 1976.920 2392.250 ;
        RECT 1976.720 19.390 1976.980 19.710 ;
        RECT 1995.120 19.390 1995.380 19.710 ;
        RECT 1995.180 2.400 1995.320 19.390 ;
        RECT 1994.970 -4.800 1995.530 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1146.390 1316.380 1146.710 1316.440 ;
        RECT 1997.390 1316.380 1997.710 1316.440 ;
        RECT 1146.390 1316.240 1997.710 1316.380 ;
        RECT 1146.390 1316.180 1146.710 1316.240 ;
        RECT 1997.390 1316.180 1997.710 1316.240 ;
        RECT 1997.390 20.640 1997.710 20.700 ;
        RECT 2012.570 20.640 2012.890 20.700 ;
        RECT 1997.390 20.500 2012.890 20.640 ;
        RECT 1997.390 20.440 1997.710 20.500 ;
        RECT 2012.570 20.440 2012.890 20.500 ;
      LAYER via ;
        RECT 1146.420 1316.180 1146.680 1316.440 ;
        RECT 1997.420 1316.180 1997.680 1316.440 ;
        RECT 1997.420 20.440 1997.680 20.700 ;
        RECT 2012.600 20.440 2012.860 20.700 ;
      LAYER met2 ;
        RECT 1146.460 1323.135 1146.740 1327.135 ;
        RECT 1146.480 1316.470 1146.620 1323.135 ;
        RECT 1146.420 1316.150 1146.680 1316.470 ;
        RECT 1997.420 1316.150 1997.680 1316.470 ;
        RECT 1997.480 20.730 1997.620 1316.150 ;
        RECT 1997.420 20.410 1997.680 20.730 ;
        RECT 2012.600 20.410 2012.860 20.730 ;
        RECT 2012.660 2.400 2012.800 20.410 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1545.670 1316.720 1545.990 1316.780 ;
        RECT 2004.290 1316.720 2004.610 1316.780 ;
        RECT 1545.670 1316.580 2004.610 1316.720 ;
        RECT 1545.670 1316.520 1545.990 1316.580 ;
        RECT 2004.290 1316.520 2004.610 1316.580 ;
        RECT 2004.290 20.300 2004.610 20.360 ;
        RECT 2030.510 20.300 2030.830 20.360 ;
        RECT 2004.290 20.160 2030.830 20.300 ;
        RECT 2004.290 20.100 2004.610 20.160 ;
        RECT 2030.510 20.100 2030.830 20.160 ;
      LAYER via ;
        RECT 1545.700 1316.520 1545.960 1316.780 ;
        RECT 2004.320 1316.520 2004.580 1316.780 ;
        RECT 2004.320 20.100 2004.580 20.360 ;
        RECT 2030.540 20.100 2030.800 20.360 ;
      LAYER met2 ;
        RECT 1545.740 1323.135 1546.020 1327.135 ;
        RECT 1545.760 1316.810 1545.900 1323.135 ;
        RECT 1545.700 1316.490 1545.960 1316.810 ;
        RECT 2004.320 1316.490 2004.580 1316.810 ;
        RECT 2004.380 20.390 2004.520 1316.490 ;
        RECT 2004.320 20.070 2004.580 20.390 ;
        RECT 2030.540 20.070 2030.800 20.390 ;
        RECT 2030.600 2.400 2030.740 20.070 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 759.070 1311.620 759.390 1311.680 ;
        RECT 764.590 1311.620 764.910 1311.680 ;
        RECT 759.070 1311.480 764.910 1311.620 ;
        RECT 759.070 1311.420 759.390 1311.480 ;
        RECT 764.590 1311.420 764.910 1311.480 ;
        RECT 764.590 66.880 764.910 66.940 ;
        RECT 2042.470 66.880 2042.790 66.940 ;
        RECT 764.590 66.740 2042.790 66.880 ;
        RECT 764.590 66.680 764.910 66.740 ;
        RECT 2042.470 66.680 2042.790 66.740 ;
        RECT 2042.470 37.640 2042.790 37.700 ;
        RECT 2048.450 37.640 2048.770 37.700 ;
        RECT 2042.470 37.500 2048.770 37.640 ;
        RECT 2042.470 37.440 2042.790 37.500 ;
        RECT 2048.450 37.440 2048.770 37.500 ;
      LAYER via ;
        RECT 759.100 1311.420 759.360 1311.680 ;
        RECT 764.620 1311.420 764.880 1311.680 ;
        RECT 764.620 66.680 764.880 66.940 ;
        RECT 2042.500 66.680 2042.760 66.940 ;
        RECT 2042.500 37.440 2042.760 37.700 ;
        RECT 2048.480 37.440 2048.740 37.700 ;
      LAYER met2 ;
        RECT 759.140 1323.135 759.420 1327.135 ;
        RECT 759.160 1311.710 759.300 1323.135 ;
        RECT 759.100 1311.390 759.360 1311.710 ;
        RECT 764.620 1311.390 764.880 1311.710 ;
        RECT 764.680 66.970 764.820 1311.390 ;
        RECT 764.620 66.650 764.880 66.970 ;
        RECT 2042.500 66.650 2042.760 66.970 ;
        RECT 2042.560 37.730 2042.700 66.650 ;
        RECT 2042.500 37.410 2042.760 37.730 ;
        RECT 2048.480 37.410 2048.740 37.730 ;
        RECT 2048.540 2.400 2048.680 37.410 ;
        RECT 2048.330 -4.800 2048.890 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1727.905 1329.145 1728.995 1329.315 ;
        RECT 765.585 1326.085 765.755 1328.975 ;
        RECT 855.745 1326.085 855.915 1328.975 ;
        RECT 903.585 1326.085 903.755 1328.975 ;
        RECT 944.065 1327.785 944.235 1328.975 ;
        RECT 1000.185 1327.785 1000.355 1328.975 ;
        RECT 1048.945 1327.785 1049.115 1328.975 ;
        RECT 1100.465 1327.785 1100.635 1328.975 ;
        RECT 1145.545 1327.785 1145.715 1328.975 ;
        RECT 1193.385 1327.785 1193.555 1328.975 ;
        RECT 1242.145 1327.785 1242.315 1328.975 ;
        RECT 1289.985 1327.785 1290.155 1328.975 ;
        RECT 1338.745 1327.785 1338.915 1328.975 ;
        RECT 1386.585 1327.785 1386.755 1328.975 ;
        RECT 1435.345 1327.785 1435.515 1328.975 ;
        RECT 1507.565 1327.785 1507.735 1328.975 ;
        RECT 1535.165 1327.105 1535.335 1328.975 ;
        RECT 1579.785 1327.275 1579.955 1328.975 ;
        RECT 1579.325 1327.105 1579.955 1327.275 ;
        RECT 1628.545 1326.085 1628.715 1328.975 ;
        RECT 1680.525 1326.085 1680.695 1328.975 ;
        RECT 1727.905 1328.805 1728.075 1329.145 ;
        RECT 1728.825 1327.785 1728.995 1329.145 ;
        RECT 1751.825 1329.145 1752.455 1329.315 ;
        RECT 1751.825 1327.785 1751.995 1329.145 ;
      LAYER mcon ;
        RECT 765.585 1328.805 765.755 1328.975 ;
        RECT 855.745 1328.805 855.915 1328.975 ;
        RECT 903.585 1328.805 903.755 1328.975 ;
        RECT 944.065 1328.805 944.235 1328.975 ;
        RECT 1000.185 1328.805 1000.355 1328.975 ;
        RECT 1048.945 1328.805 1049.115 1328.975 ;
        RECT 1100.465 1328.805 1100.635 1328.975 ;
        RECT 1145.545 1328.805 1145.715 1328.975 ;
        RECT 1193.385 1328.805 1193.555 1328.975 ;
        RECT 1242.145 1328.805 1242.315 1328.975 ;
        RECT 1289.985 1328.805 1290.155 1328.975 ;
        RECT 1338.745 1328.805 1338.915 1328.975 ;
        RECT 1386.585 1328.805 1386.755 1328.975 ;
        RECT 1435.345 1328.805 1435.515 1328.975 ;
        RECT 1507.565 1328.805 1507.735 1328.975 ;
        RECT 1535.165 1328.805 1535.335 1328.975 ;
        RECT 1579.785 1328.805 1579.955 1328.975 ;
        RECT 1628.545 1328.805 1628.715 1328.975 ;
        RECT 1680.525 1328.805 1680.695 1328.975 ;
        RECT 1752.285 1329.145 1752.455 1329.315 ;
      LAYER met1 ;
        RECT 1768.310 1566.620 1768.630 1566.680 ;
        RECT 1778.890 1566.620 1779.210 1566.680 ;
        RECT 1768.310 1566.480 1779.210 1566.620 ;
        RECT 1768.310 1566.420 1768.630 1566.480 ;
        RECT 1778.890 1566.420 1779.210 1566.480 ;
        RECT 1752.225 1329.300 1752.515 1329.345 ;
        RECT 1778.890 1329.300 1779.210 1329.360 ;
        RECT 1752.225 1329.160 1779.210 1329.300 ;
        RECT 1752.225 1329.115 1752.515 1329.160 ;
        RECT 1778.890 1329.100 1779.210 1329.160 ;
        RECT 765.525 1328.960 765.815 1329.005 ;
        RECT 855.685 1328.960 855.975 1329.005 ;
        RECT 765.525 1328.820 855.975 1328.960 ;
        RECT 765.525 1328.775 765.815 1328.820 ;
        RECT 855.685 1328.775 855.975 1328.820 ;
        RECT 903.525 1328.960 903.815 1329.005 ;
        RECT 944.005 1328.960 944.295 1329.005 ;
        RECT 903.525 1328.820 944.295 1328.960 ;
        RECT 903.525 1328.775 903.815 1328.820 ;
        RECT 944.005 1328.775 944.295 1328.820 ;
        RECT 1000.125 1328.960 1000.415 1329.005 ;
        RECT 1048.885 1328.960 1049.175 1329.005 ;
        RECT 1000.125 1328.820 1049.175 1328.960 ;
        RECT 1000.125 1328.775 1000.415 1328.820 ;
        RECT 1048.885 1328.775 1049.175 1328.820 ;
        RECT 1100.405 1328.960 1100.695 1329.005 ;
        RECT 1145.485 1328.960 1145.775 1329.005 ;
        RECT 1100.405 1328.820 1145.775 1328.960 ;
        RECT 1100.405 1328.775 1100.695 1328.820 ;
        RECT 1145.485 1328.775 1145.775 1328.820 ;
        RECT 1193.325 1328.960 1193.615 1329.005 ;
        RECT 1242.085 1328.960 1242.375 1329.005 ;
        RECT 1193.325 1328.820 1242.375 1328.960 ;
        RECT 1193.325 1328.775 1193.615 1328.820 ;
        RECT 1242.085 1328.775 1242.375 1328.820 ;
        RECT 1289.925 1328.960 1290.215 1329.005 ;
        RECT 1338.685 1328.960 1338.975 1329.005 ;
        RECT 1289.925 1328.820 1338.975 1328.960 ;
        RECT 1289.925 1328.775 1290.215 1328.820 ;
        RECT 1338.685 1328.775 1338.975 1328.820 ;
        RECT 1386.525 1328.960 1386.815 1329.005 ;
        RECT 1435.285 1328.960 1435.575 1329.005 ;
        RECT 1386.525 1328.820 1435.575 1328.960 ;
        RECT 1386.525 1328.775 1386.815 1328.820 ;
        RECT 1435.285 1328.775 1435.575 1328.820 ;
        RECT 1507.505 1328.960 1507.795 1329.005 ;
        RECT 1535.105 1328.960 1535.395 1329.005 ;
        RECT 1507.505 1328.820 1535.395 1328.960 ;
        RECT 1507.505 1328.775 1507.795 1328.820 ;
        RECT 1535.105 1328.775 1535.395 1328.820 ;
        RECT 1579.725 1328.960 1580.015 1329.005 ;
        RECT 1628.485 1328.960 1628.775 1329.005 ;
        RECT 1579.725 1328.820 1628.775 1328.960 ;
        RECT 1579.725 1328.775 1580.015 1328.820 ;
        RECT 1628.485 1328.775 1628.775 1328.820 ;
        RECT 1680.465 1328.960 1680.755 1329.005 ;
        RECT 1727.845 1328.960 1728.135 1329.005 ;
        RECT 1680.465 1328.820 1728.135 1328.960 ;
        RECT 1680.465 1328.775 1680.755 1328.820 ;
        RECT 1727.845 1328.775 1728.135 1328.820 ;
        RECT 944.005 1327.940 944.295 1327.985 ;
        RECT 1000.125 1327.940 1000.415 1327.985 ;
        RECT 944.005 1327.800 1000.415 1327.940 ;
        RECT 944.005 1327.755 944.295 1327.800 ;
        RECT 1000.125 1327.755 1000.415 1327.800 ;
        RECT 1048.885 1327.940 1049.175 1327.985 ;
        RECT 1100.405 1327.940 1100.695 1327.985 ;
        RECT 1048.885 1327.800 1100.695 1327.940 ;
        RECT 1048.885 1327.755 1049.175 1327.800 ;
        RECT 1100.405 1327.755 1100.695 1327.800 ;
        RECT 1145.485 1327.940 1145.775 1327.985 ;
        RECT 1193.325 1327.940 1193.615 1327.985 ;
        RECT 1145.485 1327.800 1193.615 1327.940 ;
        RECT 1145.485 1327.755 1145.775 1327.800 ;
        RECT 1193.325 1327.755 1193.615 1327.800 ;
        RECT 1242.085 1327.940 1242.375 1327.985 ;
        RECT 1289.925 1327.940 1290.215 1327.985 ;
        RECT 1242.085 1327.800 1290.215 1327.940 ;
        RECT 1242.085 1327.755 1242.375 1327.800 ;
        RECT 1289.925 1327.755 1290.215 1327.800 ;
        RECT 1338.685 1327.940 1338.975 1327.985 ;
        RECT 1386.525 1327.940 1386.815 1327.985 ;
        RECT 1338.685 1327.800 1386.815 1327.940 ;
        RECT 1338.685 1327.755 1338.975 1327.800 ;
        RECT 1386.525 1327.755 1386.815 1327.800 ;
        RECT 1435.285 1327.940 1435.575 1327.985 ;
        RECT 1507.505 1327.940 1507.795 1327.985 ;
        RECT 1435.285 1327.800 1507.795 1327.940 ;
        RECT 1435.285 1327.755 1435.575 1327.800 ;
        RECT 1507.505 1327.755 1507.795 1327.800 ;
        RECT 1728.765 1327.940 1729.055 1327.985 ;
        RECT 1751.765 1327.940 1752.055 1327.985 ;
        RECT 1728.765 1327.800 1752.055 1327.940 ;
        RECT 1728.765 1327.755 1729.055 1327.800 ;
        RECT 1751.765 1327.755 1752.055 1327.800 ;
        RECT 1535.105 1327.260 1535.395 1327.305 ;
        RECT 1579.265 1327.260 1579.555 1327.305 ;
        RECT 1535.105 1327.120 1579.555 1327.260 ;
        RECT 1535.105 1327.075 1535.395 1327.120 ;
        RECT 1579.265 1327.075 1579.555 1327.120 ;
        RECT 765.510 1326.240 765.830 1326.300 ;
        RECT 765.315 1326.100 765.830 1326.240 ;
        RECT 765.510 1326.040 765.830 1326.100 ;
        RECT 855.685 1326.240 855.975 1326.285 ;
        RECT 903.525 1326.240 903.815 1326.285 ;
        RECT 855.685 1326.100 903.815 1326.240 ;
        RECT 855.685 1326.055 855.975 1326.100 ;
        RECT 903.525 1326.055 903.815 1326.100 ;
        RECT 1628.485 1326.240 1628.775 1326.285 ;
        RECT 1680.465 1326.240 1680.755 1326.285 ;
        RECT 1628.485 1326.100 1680.755 1326.240 ;
        RECT 1628.485 1326.055 1628.775 1326.100 ;
        RECT 1680.465 1326.055 1680.755 1326.100 ;
      LAYER via ;
        RECT 1768.340 1566.420 1768.600 1566.680 ;
        RECT 1778.920 1566.420 1779.180 1566.680 ;
        RECT 1778.920 1329.100 1779.180 1329.360 ;
        RECT 765.540 1326.040 765.800 1326.300 ;
      LAYER met2 ;
        RECT 1768.330 1569.595 1768.610 1569.965 ;
        RECT 1768.400 1566.710 1768.540 1569.595 ;
        RECT 1768.340 1566.390 1768.600 1566.710 ;
        RECT 1778.920 1566.390 1779.180 1566.710 ;
        RECT 1778.980 1329.390 1779.120 1566.390 ;
        RECT 1778.920 1329.070 1779.180 1329.390 ;
        RECT 765.540 1326.010 765.800 1326.330 ;
        RECT 765.600 6.530 765.740 1326.010 ;
        RECT 763.760 6.390 765.740 6.530 ;
        RECT 763.760 2.400 763.900 6.390 ;
        RECT 763.550 -4.800 764.110 2.400 ;
      LAYER via2 ;
        RECT 1768.330 1569.640 1768.610 1569.920 ;
      LAYER met3 ;
        RECT 1755.835 1569.930 1759.835 1569.935 ;
        RECT 1768.305 1569.930 1768.635 1569.945 ;
        RECT 1755.835 1569.630 1768.635 1569.930 ;
        RECT 1755.835 1569.335 1759.835 1569.630 ;
        RECT 1768.305 1569.615 1768.635 1569.630 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 720.045 1307.385 720.215 1340.195 ;
      LAYER mcon ;
        RECT 720.045 1340.025 720.215 1340.195 ;
      LAYER met1 ;
        RECT 717.210 1432.320 717.530 1432.380 ;
        RECT 719.970 1432.320 720.290 1432.380 ;
        RECT 717.210 1432.180 720.290 1432.320 ;
        RECT 717.210 1432.120 717.530 1432.180 ;
        RECT 719.970 1432.120 720.290 1432.180 ;
        RECT 719.970 1340.180 720.290 1340.240 ;
        RECT 719.775 1340.040 720.290 1340.180 ;
        RECT 719.970 1339.980 720.290 1340.040 ;
        RECT 719.970 1307.540 720.290 1307.600 ;
        RECT 719.775 1307.400 720.290 1307.540 ;
        RECT 719.970 1307.340 720.290 1307.400 ;
        RECT 719.970 60.760 720.290 60.820 ;
        RECT 2065.930 60.760 2066.250 60.820 ;
        RECT 719.970 60.620 2066.250 60.760 ;
        RECT 719.970 60.560 720.290 60.620 ;
        RECT 2065.930 60.560 2066.250 60.620 ;
      LAYER via ;
        RECT 717.240 1432.120 717.500 1432.380 ;
        RECT 720.000 1432.120 720.260 1432.380 ;
        RECT 720.000 1339.980 720.260 1340.240 ;
        RECT 720.000 1307.340 720.260 1307.600 ;
        RECT 720.000 60.560 720.260 60.820 ;
        RECT 2065.960 60.560 2066.220 60.820 ;
      LAYER met2 ;
        RECT 717.230 1468.955 717.510 1469.325 ;
        RECT 717.300 1432.410 717.440 1468.955 ;
        RECT 717.240 1432.090 717.500 1432.410 ;
        RECT 720.000 1432.090 720.260 1432.410 ;
        RECT 720.060 1340.270 720.200 1432.090 ;
        RECT 720.000 1339.950 720.260 1340.270 ;
        RECT 720.000 1307.310 720.260 1307.630 ;
        RECT 720.060 60.850 720.200 1307.310 ;
        RECT 720.000 60.530 720.260 60.850 ;
        RECT 2065.960 60.530 2066.220 60.850 ;
        RECT 2066.020 20.130 2066.160 60.530 ;
        RECT 2066.020 19.990 2066.620 20.130 ;
        RECT 2066.480 2.400 2066.620 19.990 ;
        RECT 2066.270 -4.800 2066.830 2.400 ;
      LAYER via2 ;
        RECT 717.230 1469.000 717.510 1469.280 ;
      LAYER met3 ;
        RECT 715.810 1471.415 719.810 1472.015 ;
        RECT 716.990 1469.305 717.290 1471.415 ;
        RECT 716.990 1468.990 717.535 1469.305 ;
        RECT 717.205 1468.975 717.535 1468.990 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1058.990 1315.700 1059.310 1315.760 ;
        RECT 2066.390 1315.700 2066.710 1315.760 ;
        RECT 1058.990 1315.560 2066.710 1315.700 ;
        RECT 1058.990 1315.500 1059.310 1315.560 ;
        RECT 2066.390 1315.500 2066.710 1315.560 ;
        RECT 2066.390 20.640 2066.710 20.700 ;
        RECT 2084.330 20.640 2084.650 20.700 ;
        RECT 2066.390 20.500 2084.650 20.640 ;
        RECT 2066.390 20.440 2066.710 20.500 ;
        RECT 2084.330 20.440 2084.650 20.500 ;
      LAYER via ;
        RECT 1059.020 1315.500 1059.280 1315.760 ;
        RECT 2066.420 1315.500 2066.680 1315.760 ;
        RECT 2066.420 20.440 2066.680 20.700 ;
        RECT 2084.360 20.440 2084.620 20.700 ;
      LAYER met2 ;
        RECT 1059.060 1323.135 1059.340 1327.135 ;
        RECT 1059.080 1315.790 1059.220 1323.135 ;
        RECT 1059.020 1315.470 1059.280 1315.790 ;
        RECT 2066.420 1315.470 2066.680 1315.790 ;
        RECT 2066.480 20.730 2066.620 1315.470 ;
        RECT 2066.420 20.410 2066.680 20.730 ;
        RECT 2084.360 20.410 2084.620 20.730 ;
        RECT 2084.420 2.400 2084.560 20.410 ;
        RECT 2084.210 -4.800 2084.770 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1354.310 1316.040 1354.630 1316.100 ;
        RECT 2087.550 1316.040 2087.870 1316.100 ;
        RECT 1354.310 1315.900 2087.870 1316.040 ;
        RECT 1354.310 1315.840 1354.630 1315.900 ;
        RECT 2087.550 1315.840 2087.870 1315.900 ;
        RECT 2087.550 15.880 2087.870 15.940 ;
        RECT 2101.810 15.880 2102.130 15.940 ;
        RECT 2087.550 15.740 2102.130 15.880 ;
        RECT 2087.550 15.680 2087.870 15.740 ;
        RECT 2101.810 15.680 2102.130 15.740 ;
      LAYER via ;
        RECT 1354.340 1315.840 1354.600 1316.100 ;
        RECT 2087.580 1315.840 2087.840 1316.100 ;
        RECT 2087.580 15.680 2087.840 15.940 ;
        RECT 2101.840 15.680 2102.100 15.940 ;
      LAYER met2 ;
        RECT 1354.380 1323.135 1354.660 1327.135 ;
        RECT 1354.400 1316.130 1354.540 1323.135 ;
        RECT 1354.340 1315.810 1354.600 1316.130 ;
        RECT 2087.580 1315.810 2087.840 1316.130 ;
        RECT 2087.640 15.970 2087.780 1315.810 ;
        RECT 2087.580 15.650 2087.840 15.970 ;
        RECT 2101.840 15.650 2102.100 15.970 ;
        RECT 2101.900 2.400 2102.040 15.650 ;
        RECT 2101.690 -4.800 2102.250 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1542.910 2390.100 1543.230 2390.160 ;
        RECT 2100.890 2390.100 2101.210 2390.160 ;
        RECT 1542.910 2389.960 2101.210 2390.100 ;
        RECT 1542.910 2389.900 1543.230 2389.960 ;
        RECT 2100.890 2389.900 2101.210 2389.960 ;
        RECT 2100.890 20.640 2101.210 20.700 ;
        RECT 2119.750 20.640 2120.070 20.700 ;
        RECT 2100.890 20.500 2120.070 20.640 ;
        RECT 2100.890 20.440 2101.210 20.500 ;
        RECT 2119.750 20.440 2120.070 20.500 ;
      LAYER via ;
        RECT 1542.940 2389.900 1543.200 2390.160 ;
        RECT 2100.920 2389.900 2101.180 2390.160 ;
        RECT 2100.920 20.440 2101.180 20.700 ;
        RECT 2119.780 20.440 2120.040 20.700 ;
      LAYER met2 ;
        RECT 1542.940 2389.870 1543.200 2390.190 ;
        RECT 2100.920 2389.870 2101.180 2390.190 ;
        RECT 1543.000 2377.880 1543.140 2389.870 ;
        RECT 1542.980 2373.880 1543.260 2377.880 ;
        RECT 2100.980 20.730 2101.120 2389.870 ;
        RECT 2100.920 20.410 2101.180 20.730 ;
        RECT 2119.780 20.410 2120.040 20.730 ;
        RECT 2119.840 2.400 2119.980 20.410 ;
        RECT 2119.630 -4.800 2120.190 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2132.190 1300.995 2132.470 1301.365 ;
        RECT 2132.260 16.730 2132.400 1300.995 ;
        RECT 2132.260 16.590 2137.920 16.730 ;
        RECT 2137.780 2.400 2137.920 16.590 ;
        RECT 2137.570 -4.800 2138.130 2.400 ;
      LAYER via2 ;
        RECT 2132.190 1301.040 2132.470 1301.320 ;
      LAYER met3 ;
        RECT 705.910 1874.570 706.290 1874.580 ;
        RECT 715.810 1874.570 719.810 1874.575 ;
        RECT 705.910 1874.270 719.810 1874.570 ;
        RECT 705.910 1874.260 706.290 1874.270 ;
        RECT 715.810 1873.975 719.810 1874.270 ;
        RECT 705.910 1301.330 706.290 1301.340 ;
        RECT 2132.165 1301.330 2132.495 1301.345 ;
        RECT 705.910 1301.030 2132.495 1301.330 ;
        RECT 705.910 1301.020 706.290 1301.030 ;
        RECT 2132.165 1301.015 2132.495 1301.030 ;
      LAYER via3 ;
        RECT 705.940 1874.260 706.260 1874.580 ;
        RECT 705.940 1301.020 706.260 1301.340 ;
      LAYER met4 ;
        RECT 705.935 1874.255 706.265 1874.585 ;
        RECT 705.950 1301.345 706.250 1874.255 ;
        RECT 705.935 1301.015 706.265 1301.345 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1772.910 1870.240 1773.230 1870.300 ;
        RECT 2135.390 1870.240 2135.710 1870.300 ;
        RECT 1772.910 1870.100 2135.710 1870.240 ;
        RECT 1772.910 1870.040 1773.230 1870.100 ;
        RECT 2135.390 1870.040 2135.710 1870.100 ;
        RECT 2135.390 19.960 2135.710 20.020 ;
        RECT 2155.630 19.960 2155.950 20.020 ;
        RECT 2135.390 19.820 2155.950 19.960 ;
        RECT 2135.390 19.760 2135.710 19.820 ;
        RECT 2155.630 19.760 2155.950 19.820 ;
      LAYER via ;
        RECT 1772.940 1870.040 1773.200 1870.300 ;
        RECT 2135.420 1870.040 2135.680 1870.300 ;
        RECT 2135.420 19.760 2135.680 20.020 ;
        RECT 2155.660 19.760 2155.920 20.020 ;
      LAYER met2 ;
        RECT 1772.930 1870.155 1773.210 1870.525 ;
        RECT 1772.940 1870.010 1773.200 1870.155 ;
        RECT 2135.420 1870.010 2135.680 1870.330 ;
        RECT 2135.480 20.050 2135.620 1870.010 ;
        RECT 2135.420 19.730 2135.680 20.050 ;
        RECT 2155.660 19.730 2155.920 20.050 ;
        RECT 2155.720 2.400 2155.860 19.730 ;
        RECT 2155.510 -4.800 2156.070 2.400 ;
      LAYER via2 ;
        RECT 1772.930 1870.200 1773.210 1870.480 ;
      LAYER met3 ;
        RECT 1755.835 1870.490 1759.835 1870.495 ;
        RECT 1772.905 1870.490 1773.235 1870.505 ;
        RECT 1755.835 1870.190 1773.235 1870.490 ;
        RECT 1755.835 1869.895 1759.835 1870.190 ;
        RECT 1772.905 1870.175 1773.235 1870.190 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1366.270 1315.360 1366.590 1315.420 ;
        RECT 2156.090 1315.360 2156.410 1315.420 ;
        RECT 1366.270 1315.220 2156.410 1315.360 ;
        RECT 1366.270 1315.160 1366.590 1315.220 ;
        RECT 2156.090 1315.160 2156.410 1315.220 ;
        RECT 2156.090 20.640 2156.410 20.700 ;
        RECT 2173.110 20.640 2173.430 20.700 ;
        RECT 2156.090 20.500 2173.430 20.640 ;
        RECT 2156.090 20.440 2156.410 20.500 ;
        RECT 2173.110 20.440 2173.430 20.500 ;
      LAYER via ;
        RECT 1366.300 1315.160 1366.560 1315.420 ;
        RECT 2156.120 1315.160 2156.380 1315.420 ;
        RECT 2156.120 20.440 2156.380 20.700 ;
        RECT 2173.140 20.440 2173.400 20.700 ;
      LAYER met2 ;
        RECT 1366.340 1323.135 1366.620 1327.135 ;
        RECT 1366.360 1315.450 1366.500 1323.135 ;
        RECT 1366.300 1315.130 1366.560 1315.450 ;
        RECT 2156.120 1315.130 2156.380 1315.450 ;
        RECT 2156.180 20.730 2156.320 1315.130 ;
        RECT 2156.120 20.410 2156.380 20.730 ;
        RECT 2173.140 20.410 2173.400 20.730 ;
        RECT 2173.200 2.400 2173.340 20.410 ;
        RECT 2172.990 -4.800 2173.550 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2187.390 72.235 2187.670 72.605 ;
        RECT 2187.460 24.210 2187.600 72.235 ;
        RECT 2187.460 24.070 2191.280 24.210 ;
        RECT 2191.140 2.400 2191.280 24.070 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
      LAYER via2 ;
        RECT 2187.390 72.280 2187.670 72.560 ;
      LAYER met3 ;
        RECT 701.310 2165.610 701.690 2165.620 ;
        RECT 715.810 2165.610 719.810 2165.615 ;
        RECT 701.310 2165.310 719.810 2165.610 ;
        RECT 701.310 2165.300 701.690 2165.310 ;
        RECT 715.810 2165.015 719.810 2165.310 ;
        RECT 701.310 72.570 701.690 72.580 ;
        RECT 2187.365 72.570 2187.695 72.585 ;
        RECT 701.310 72.270 2187.695 72.570 ;
        RECT 701.310 72.260 701.690 72.270 ;
        RECT 2187.365 72.255 2187.695 72.270 ;
      LAYER via3 ;
        RECT 701.340 2165.300 701.660 2165.620 ;
        RECT 701.340 72.260 701.660 72.580 ;
      LAYER met4 ;
        RECT 701.335 2165.295 701.665 2165.625 ;
        RECT 701.350 72.585 701.650 2165.295 ;
        RECT 701.335 72.255 701.665 72.585 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1441.710 73.340 1442.030 73.400 ;
        RECT 2208.070 73.340 2208.390 73.400 ;
        RECT 1441.710 73.200 2208.390 73.340 ;
        RECT 1441.710 73.140 1442.030 73.200 ;
        RECT 2208.070 73.140 2208.390 73.200 ;
      LAYER via ;
        RECT 1441.740 73.140 1442.000 73.400 ;
        RECT 2208.100 73.140 2208.360 73.400 ;
      LAYER met2 ;
        RECT 1441.780 1323.135 1442.060 1327.135 ;
        RECT 1441.800 73.430 1441.940 1323.135 ;
        RECT 1441.740 73.110 1442.000 73.430 ;
        RECT 2208.100 73.110 2208.360 73.430 ;
        RECT 2208.160 16.730 2208.300 73.110 ;
        RECT 2208.160 16.590 2209.220 16.730 ;
        RECT 2209.080 2.400 2209.220 16.590 ;
        RECT 2208.870 -4.800 2209.430 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2221.890 80.395 2222.170 80.765 ;
        RECT 2221.960 16.730 2222.100 80.395 ;
        RECT 2221.960 16.590 2227.160 16.730 ;
        RECT 2227.020 2.400 2227.160 16.590 ;
        RECT 2226.810 -4.800 2227.370 2.400 ;
      LAYER via2 ;
        RECT 2221.890 80.440 2222.170 80.720 ;
      LAYER met3 ;
        RECT 700.390 2020.090 700.770 2020.100 ;
        RECT 715.810 2020.090 719.810 2020.095 ;
        RECT 700.390 2019.790 719.810 2020.090 ;
        RECT 700.390 2019.780 700.770 2019.790 ;
        RECT 715.810 2019.495 719.810 2019.790 ;
        RECT 700.390 80.730 700.770 80.740 ;
        RECT 2221.865 80.730 2222.195 80.745 ;
        RECT 700.390 80.430 2222.195 80.730 ;
        RECT 700.390 80.420 700.770 80.430 ;
        RECT 2221.865 80.415 2222.195 80.430 ;
      LAYER via3 ;
        RECT 700.420 2019.780 700.740 2020.100 ;
        RECT 700.420 80.420 700.740 80.740 ;
      LAYER met4 ;
        RECT 700.415 2019.775 700.745 2020.105 ;
        RECT 700.430 80.745 700.730 2019.775 ;
        RECT 700.415 80.415 700.745 80.745 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 714.450 1322.500 714.770 1322.560 ;
        RECT 780.230 1322.500 780.550 1322.560 ;
        RECT 714.450 1322.360 780.550 1322.500 ;
        RECT 714.450 1322.300 714.770 1322.360 ;
        RECT 780.230 1322.300 780.550 1322.360 ;
      LAYER via ;
        RECT 714.480 1322.300 714.740 1322.560 ;
        RECT 780.260 1322.300 780.520 1322.560 ;
      LAYER met2 ;
        RECT 714.470 2327.115 714.750 2327.485 ;
        RECT 714.540 1322.590 714.680 2327.115 ;
        RECT 714.480 1322.270 714.740 1322.590 ;
        RECT 780.260 1322.270 780.520 1322.590 ;
        RECT 780.320 7.210 780.460 1322.270 ;
        RECT 780.320 7.070 781.840 7.210 ;
        RECT 781.700 2.400 781.840 7.070 ;
        RECT 781.490 -4.800 782.050 2.400 ;
      LAYER via2 ;
        RECT 714.470 2327.160 714.750 2327.440 ;
      LAYER met3 ;
        RECT 714.445 2327.450 714.775 2327.465 ;
        RECT 715.810 2327.450 719.810 2327.455 ;
        RECT 714.445 2327.150 719.810 2327.450 ;
        RECT 714.445 2327.135 714.775 2327.150 ;
        RECT 715.810 2326.855 719.810 2327.150 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 721.420 2374.970 721.700 2377.880 ;
        RECT 722.750 2374.970 723.030 2375.085 ;
        RECT 721.420 2374.830 723.030 2374.970 ;
        RECT 721.420 2373.880 721.700 2374.830 ;
        RECT 722.750 2374.715 723.030 2374.830 ;
        RECT 2244.890 17.835 2245.170 18.205 ;
        RECT 2244.960 2.400 2245.100 17.835 ;
        RECT 2244.750 -4.800 2245.310 2.400 ;
      LAYER via2 ;
        RECT 722.750 2374.760 723.030 2375.040 ;
        RECT 2244.890 17.880 2245.170 18.160 ;
      LAYER met3 ;
        RECT 722.725 2375.050 723.055 2375.065 ;
        RECT 736.270 2375.050 736.650 2375.060 ;
        RECT 722.725 2374.750 736.650 2375.050 ;
        RECT 722.725 2374.735 723.055 2374.750 ;
        RECT 736.270 2374.740 736.650 2374.750 ;
        RECT 1776.790 2222.420 1777.170 2222.740 ;
        RECT 1776.830 2221.380 1777.130 2222.420 ;
        RECT 1776.790 2221.060 1777.170 2221.380 ;
        RECT 1776.790 959.660 1777.170 959.980 ;
        RECT 1776.830 958.620 1777.130 959.660 ;
        RECT 1776.790 958.300 1777.170 958.620 ;
        RECT 1776.790 18.170 1777.170 18.180 ;
        RECT 2244.865 18.170 2245.195 18.185 ;
        RECT 1776.790 17.870 2245.195 18.170 ;
        RECT 1776.790 17.860 1777.170 17.870 ;
        RECT 2244.865 17.855 2245.195 17.870 ;
      LAYER via3 ;
        RECT 736.300 2374.740 736.620 2375.060 ;
        RECT 1776.820 2222.420 1777.140 2222.740 ;
        RECT 1776.820 2221.060 1777.140 2221.380 ;
        RECT 1776.820 959.660 1777.140 959.980 ;
        RECT 1776.820 958.300 1777.140 958.620 ;
        RECT 1776.820 17.860 1777.140 18.180 ;
      LAYER met4 ;
        RECT 735.870 2374.310 737.050 2375.490 ;
        RECT 1776.390 2374.310 1777.570 2375.490 ;
        RECT 1776.830 2222.745 1777.130 2374.310 ;
        RECT 1776.815 2222.415 1777.145 2222.745 ;
        RECT 1776.815 2221.055 1777.145 2221.385 ;
        RECT 1776.830 959.985 1777.130 2221.055 ;
        RECT 1776.815 959.655 1777.145 959.985 ;
        RECT 1776.815 958.295 1777.145 958.625 ;
        RECT 1776.830 18.185 1777.130 958.295 ;
        RECT 1776.815 17.855 1777.145 18.185 ;
      LAYER met5 ;
        RECT 735.660 2374.100 1777.780 2375.700 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 712.685 1423.665 712.855 1430.295 ;
        RECT 719.585 1339.345 719.755 1401.735 ;
      LAYER mcon ;
        RECT 712.685 1430.125 712.855 1430.295 ;
        RECT 719.585 1401.565 719.755 1401.735 ;
      LAYER met1 ;
        RECT 712.610 1430.280 712.930 1430.340 ;
        RECT 712.415 1430.140 712.930 1430.280 ;
        RECT 712.610 1430.080 712.930 1430.140 ;
        RECT 712.610 1423.820 712.930 1423.880 ;
        RECT 712.415 1423.680 712.930 1423.820 ;
        RECT 712.610 1423.620 712.930 1423.680 ;
        RECT 712.610 1401.720 712.930 1401.780 ;
        RECT 719.525 1401.720 719.815 1401.765 ;
        RECT 712.610 1401.580 719.815 1401.720 ;
        RECT 712.610 1401.520 712.930 1401.580 ;
        RECT 719.525 1401.535 719.815 1401.580 ;
        RECT 719.050 1339.500 719.370 1339.560 ;
        RECT 719.525 1339.500 719.815 1339.545 ;
        RECT 719.050 1339.360 719.815 1339.500 ;
        RECT 719.050 1339.300 719.370 1339.360 ;
        RECT 719.525 1339.315 719.815 1339.360 ;
      LAYER via ;
        RECT 712.640 1430.080 712.900 1430.340 ;
        RECT 712.640 1423.620 712.900 1423.880 ;
        RECT 712.640 1401.520 712.900 1401.780 ;
        RECT 719.080 1339.300 719.340 1339.560 ;
      LAYER met2 ;
        RECT 712.630 1451.275 712.910 1451.645 ;
        RECT 712.700 1430.370 712.840 1451.275 ;
        RECT 712.640 1430.050 712.900 1430.370 ;
        RECT 712.640 1423.590 712.900 1423.910 ;
        RECT 712.700 1401.810 712.840 1423.590 ;
        RECT 712.640 1401.490 712.900 1401.810 ;
        RECT 719.080 1339.445 719.340 1339.590 ;
        RECT 719.070 1339.075 719.350 1339.445 ;
        RECT 2256.850 58.635 2257.130 59.005 ;
        RECT 2256.920 5.850 2257.060 58.635 ;
        RECT 2256.920 5.710 2262.580 5.850 ;
        RECT 2262.440 2.400 2262.580 5.710 ;
        RECT 2262.230 -4.800 2262.790 2.400 ;
      LAYER via2 ;
        RECT 712.630 1451.320 712.910 1451.600 ;
        RECT 719.070 1339.120 719.350 1339.400 ;
        RECT 2256.850 58.680 2257.130 58.960 ;
      LAYER met3 ;
        RECT 715.810 1455.095 719.810 1455.695 ;
        RECT 712.605 1451.610 712.935 1451.625 ;
        RECT 717.910 1451.610 718.210 1455.095 ;
        RECT 712.605 1451.310 718.210 1451.610 ;
        RECT 712.605 1451.295 712.935 1451.310 ;
        RECT 717.870 1339.410 718.250 1339.420 ;
        RECT 719.045 1339.410 719.375 1339.425 ;
        RECT 717.870 1339.110 719.375 1339.410 ;
        RECT 717.870 1339.100 718.250 1339.110 ;
        RECT 719.045 1339.095 719.375 1339.110 ;
        RECT 719.710 546.220 720.090 546.540 ;
        RECT 719.750 545.180 720.050 546.220 ;
        RECT 719.710 544.860 720.090 545.180 ;
        RECT 719.710 58.970 720.090 58.980 ;
        RECT 2256.825 58.970 2257.155 58.985 ;
        RECT 719.710 58.670 2257.155 58.970 ;
        RECT 719.710 58.660 720.090 58.670 ;
        RECT 2256.825 58.655 2257.155 58.670 ;
      LAYER via3 ;
        RECT 717.900 1339.100 718.220 1339.420 ;
        RECT 719.740 546.220 720.060 546.540 ;
        RECT 719.740 544.860 720.060 545.180 ;
        RECT 719.740 58.660 720.060 58.980 ;
      LAYER met4 ;
        RECT 717.910 1341.150 720.050 1341.450 ;
        RECT 717.910 1339.425 718.210 1341.150 ;
        RECT 717.895 1339.095 718.225 1339.425 ;
        RECT 719.750 546.545 720.050 1341.150 ;
        RECT 719.735 546.215 720.065 546.545 ;
        RECT 719.735 544.855 720.065 545.185 ;
        RECT 719.750 158.930 720.050 544.855 ;
        RECT 718.830 158.630 720.050 158.930 ;
        RECT 718.830 154.850 719.130 158.630 ;
        RECT 718.830 154.550 720.050 154.850 ;
        RECT 719.750 58.985 720.050 154.550 ;
        RECT 719.735 58.655 720.065 58.985 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1772.910 1787.280 1773.230 1787.340 ;
        RECT 2259.590 1787.280 2259.910 1787.340 ;
        RECT 1772.910 1787.140 2259.910 1787.280 ;
        RECT 1772.910 1787.080 1773.230 1787.140 ;
        RECT 2259.590 1787.080 2259.910 1787.140 ;
        RECT 2259.590 18.260 2259.910 18.320 ;
        RECT 2280.290 18.260 2280.610 18.320 ;
        RECT 2259.590 18.120 2280.610 18.260 ;
        RECT 2259.590 18.060 2259.910 18.120 ;
        RECT 2280.290 18.060 2280.610 18.120 ;
      LAYER via ;
        RECT 1772.940 1787.080 1773.200 1787.340 ;
        RECT 2259.620 1787.080 2259.880 1787.340 ;
        RECT 2259.620 18.060 2259.880 18.320 ;
        RECT 2280.320 18.060 2280.580 18.320 ;
      LAYER met2 ;
        RECT 1772.930 1792.635 1773.210 1793.005 ;
        RECT 1773.000 1787.370 1773.140 1792.635 ;
        RECT 1772.940 1787.050 1773.200 1787.370 ;
        RECT 2259.620 1787.050 2259.880 1787.370 ;
        RECT 2259.680 18.350 2259.820 1787.050 ;
        RECT 2259.620 18.030 2259.880 18.350 ;
        RECT 2280.320 18.030 2280.580 18.350 ;
        RECT 2280.380 2.400 2280.520 18.030 ;
        RECT 2280.170 -4.800 2280.730 2.400 ;
      LAYER via2 ;
        RECT 1772.930 1792.680 1773.210 1792.960 ;
      LAYER met3 ;
        RECT 1755.835 1792.970 1759.835 1792.975 ;
        RECT 1772.905 1792.970 1773.235 1792.985 ;
        RECT 1755.835 1792.670 1773.235 1792.970 ;
        RECT 1755.835 1792.375 1759.835 1792.670 ;
        RECT 1772.905 1792.655 1773.235 1792.670 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1121.165 2390.625 1121.335 2392.155 ;
      LAYER mcon ;
        RECT 1121.165 2391.985 1121.335 2392.155 ;
      LAYER met1 ;
        RECT 1097.630 2392.140 1097.950 2392.200 ;
        RECT 1121.105 2392.140 1121.395 2392.185 ;
        RECT 1097.630 2392.000 1121.395 2392.140 ;
        RECT 1097.630 2391.940 1097.950 2392.000 ;
        RECT 1121.105 2391.955 1121.395 2392.000 ;
        RECT 1121.105 2390.780 1121.395 2390.825 ;
        RECT 1704.370 2390.780 1704.690 2390.840 ;
        RECT 1121.105 2390.640 1704.690 2390.780 ;
        RECT 1121.105 2390.595 1121.395 2390.640 ;
        RECT 1704.370 2390.580 1704.690 2390.640 ;
        RECT 1704.370 2386.020 1704.690 2386.080 ;
        RECT 2297.770 2386.020 2298.090 2386.080 ;
        RECT 1704.370 2385.880 2298.090 2386.020 ;
        RECT 1704.370 2385.820 1704.690 2385.880 ;
        RECT 2297.770 2385.820 2298.090 2385.880 ;
      LAYER via ;
        RECT 1097.660 2391.940 1097.920 2392.200 ;
        RECT 1704.400 2390.580 1704.660 2390.840 ;
        RECT 1704.400 2385.820 1704.660 2386.080 ;
        RECT 2297.800 2385.820 2298.060 2386.080 ;
      LAYER met2 ;
        RECT 1097.660 2391.910 1097.920 2392.230 ;
        RECT 1097.720 2377.880 1097.860 2391.910 ;
        RECT 1704.400 2390.550 1704.660 2390.870 ;
        RECT 1704.460 2386.110 1704.600 2390.550 ;
        RECT 1704.400 2385.790 1704.660 2386.110 ;
        RECT 2297.800 2385.790 2298.060 2386.110 ;
        RECT 1097.700 2373.880 1097.980 2377.880 ;
        RECT 2297.860 24.210 2298.000 2385.790 ;
        RECT 2297.860 24.070 2298.460 24.210 ;
        RECT 2298.320 2.400 2298.460 24.070 ;
        RECT 2298.110 -4.800 2298.670 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1772.910 1773.680 1773.230 1773.740 ;
        RECT 2300.990 1773.680 2301.310 1773.740 ;
        RECT 1772.910 1773.540 2301.310 1773.680 ;
        RECT 1772.910 1773.480 1773.230 1773.540 ;
        RECT 2300.990 1773.480 2301.310 1773.540 ;
        RECT 2300.990 19.620 2301.310 19.680 ;
        RECT 2316.170 19.620 2316.490 19.680 ;
        RECT 2300.990 19.480 2316.490 19.620 ;
        RECT 2300.990 19.420 2301.310 19.480 ;
        RECT 2316.170 19.420 2316.490 19.480 ;
      LAYER via ;
        RECT 1772.940 1773.480 1773.200 1773.740 ;
        RECT 2301.020 1773.480 2301.280 1773.740 ;
        RECT 2301.020 19.420 2301.280 19.680 ;
        RECT 2316.200 19.420 2316.460 19.680 ;
      LAYER met2 ;
        RECT 1772.930 1774.955 1773.210 1775.325 ;
        RECT 1773.000 1773.770 1773.140 1774.955 ;
        RECT 1772.940 1773.450 1773.200 1773.770 ;
        RECT 2301.020 1773.450 2301.280 1773.770 ;
        RECT 2301.080 19.710 2301.220 1773.450 ;
        RECT 2301.020 19.390 2301.280 19.710 ;
        RECT 2316.200 19.390 2316.460 19.710 ;
        RECT 2316.260 2.400 2316.400 19.390 ;
        RECT 2316.050 -4.800 2316.610 2.400 ;
      LAYER via2 ;
        RECT 1772.930 1775.000 1773.210 1775.280 ;
      LAYER met3 ;
        RECT 1755.835 1775.290 1759.835 1775.295 ;
        RECT 1772.905 1775.290 1773.235 1775.305 ;
        RECT 1755.835 1774.990 1773.235 1775.290 ;
        RECT 1755.835 1774.695 1759.835 1774.990 ;
        RECT 1772.905 1774.975 1773.235 1774.990 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1684.590 1311.280 1684.910 1311.340 ;
        RECT 1690.110 1311.280 1690.430 1311.340 ;
        RECT 1684.590 1311.140 1690.430 1311.280 ;
        RECT 1684.590 1311.080 1684.910 1311.140 ;
        RECT 1690.110 1311.080 1690.430 1311.140 ;
        RECT 1690.110 554.240 1690.430 554.500 ;
        RECT 1690.200 553.480 1690.340 554.240 ;
        RECT 1690.110 553.220 1690.430 553.480 ;
        RECT 1690.110 53.280 1690.430 53.340 ;
        RECT 2334.110 53.280 2334.430 53.340 ;
        RECT 1690.110 53.140 2334.430 53.280 ;
        RECT 1690.110 53.080 1690.430 53.140 ;
        RECT 2334.110 53.080 2334.430 53.140 ;
      LAYER via ;
        RECT 1684.620 1311.080 1684.880 1311.340 ;
        RECT 1690.140 1311.080 1690.400 1311.340 ;
        RECT 1690.140 554.240 1690.400 554.500 ;
        RECT 1690.140 553.220 1690.400 553.480 ;
        RECT 1690.140 53.080 1690.400 53.340 ;
        RECT 2334.140 53.080 2334.400 53.340 ;
      LAYER met2 ;
        RECT 1684.660 1323.135 1684.940 1327.135 ;
        RECT 1684.680 1311.370 1684.820 1323.135 ;
        RECT 1684.620 1311.050 1684.880 1311.370 ;
        RECT 1690.140 1311.050 1690.400 1311.370 ;
        RECT 1690.200 554.530 1690.340 1311.050 ;
        RECT 1690.140 554.210 1690.400 554.530 ;
        RECT 1690.140 553.190 1690.400 553.510 ;
        RECT 1690.200 53.370 1690.340 553.190 ;
        RECT 1690.140 53.050 1690.400 53.370 ;
        RECT 2334.140 53.050 2334.400 53.370 ;
        RECT 2334.200 2.400 2334.340 53.050 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1755.505 2318.545 1755.675 2366.655 ;
      LAYER mcon ;
        RECT 1755.505 2366.485 1755.675 2366.655 ;
      LAYER met1 ;
        RECT 888.790 2389.760 889.110 2389.820 ;
        RECT 1538.310 2389.760 1538.630 2389.820 ;
        RECT 888.790 2389.620 1538.630 2389.760 ;
        RECT 888.790 2389.560 889.110 2389.620 ;
        RECT 1538.310 2389.560 1538.630 2389.620 ;
        RECT 1755.430 2366.640 1755.750 2366.700 ;
        RECT 1755.235 2366.500 1755.750 2366.640 ;
        RECT 1755.430 2366.440 1755.750 2366.500 ;
        RECT 1755.445 2318.700 1755.735 2318.745 ;
        RECT 1755.890 2318.700 1756.210 2318.760 ;
        RECT 1755.445 2318.560 1756.210 2318.700 ;
        RECT 1755.445 2318.515 1755.735 2318.560 ;
        RECT 1755.890 2318.500 1756.210 2318.560 ;
        RECT 1755.890 2294.220 1756.210 2294.280 ;
        RECT 2346.070 2294.220 2346.390 2294.280 ;
        RECT 1755.890 2294.080 2346.390 2294.220 ;
        RECT 1755.890 2294.020 1756.210 2294.080 ;
        RECT 2346.070 2294.020 2346.390 2294.080 ;
        RECT 2346.070 62.120 2346.390 62.180 ;
        RECT 2351.590 62.120 2351.910 62.180 ;
        RECT 2346.070 61.980 2351.910 62.120 ;
        RECT 2346.070 61.920 2346.390 61.980 ;
        RECT 2351.590 61.920 2351.910 61.980 ;
      LAYER via ;
        RECT 888.820 2389.560 889.080 2389.820 ;
        RECT 1538.340 2389.560 1538.600 2389.820 ;
        RECT 1755.460 2366.440 1755.720 2366.700 ;
        RECT 1755.920 2318.500 1756.180 2318.760 ;
        RECT 1755.920 2294.020 1756.180 2294.280 ;
        RECT 2346.100 2294.020 2346.360 2294.280 ;
        RECT 2346.100 61.920 2346.360 62.180 ;
        RECT 2351.620 61.920 2351.880 62.180 ;
      LAYER met2 ;
        RECT 1538.330 2391.035 1538.610 2391.405 ;
        RECT 1754.990 2391.035 1755.270 2391.405 ;
        RECT 1538.400 2389.850 1538.540 2391.035 ;
        RECT 888.820 2389.530 889.080 2389.850 ;
        RECT 1538.340 2389.530 1538.600 2389.850 ;
        RECT 888.880 2377.880 889.020 2389.530 ;
        RECT 1755.060 2378.370 1755.200 2391.035 ;
        RECT 1755.060 2378.230 1755.660 2378.370 ;
        RECT 888.860 2373.880 889.140 2377.880 ;
        RECT 1755.520 2366.730 1755.660 2378.230 ;
        RECT 1755.460 2366.410 1755.720 2366.730 ;
        RECT 1755.920 2318.470 1756.180 2318.790 ;
        RECT 1755.980 2294.310 1756.120 2318.470 ;
        RECT 1755.920 2293.990 1756.180 2294.310 ;
        RECT 2346.100 2293.990 2346.360 2294.310 ;
        RECT 2346.160 62.210 2346.300 2293.990 ;
        RECT 2346.100 61.890 2346.360 62.210 ;
        RECT 2351.620 61.890 2351.880 62.210 ;
        RECT 2351.680 2.400 2351.820 61.890 ;
        RECT 2351.470 -4.800 2352.030 2.400 ;
      LAYER via2 ;
        RECT 1538.330 2391.080 1538.610 2391.360 ;
        RECT 1754.990 2391.080 1755.270 2391.360 ;
      LAYER met3 ;
        RECT 1538.305 2391.370 1538.635 2391.385 ;
        RECT 1754.965 2391.370 1755.295 2391.385 ;
        RECT 1538.305 2391.070 1755.295 2391.370 ;
        RECT 1538.305 2391.055 1538.635 2391.070 ;
        RECT 1754.965 2391.055 1755.295 2391.070 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2366.845 2.805 2367.015 48.195 ;
      LAYER mcon ;
        RECT 2366.845 48.025 2367.015 48.195 ;
      LAYER met1 ;
        RECT 747.110 1303.460 747.430 1303.520 ;
        RECT 751.710 1303.460 752.030 1303.520 ;
        RECT 747.110 1303.320 752.030 1303.460 ;
        RECT 747.110 1303.260 747.430 1303.320 ;
        RECT 751.710 1303.260 752.030 1303.320 ;
        RECT 751.710 79.800 752.030 79.860 ;
        RECT 2366.770 79.800 2367.090 79.860 ;
        RECT 751.710 79.660 2367.090 79.800 ;
        RECT 751.710 79.600 752.030 79.660 ;
        RECT 2366.770 79.600 2367.090 79.660 ;
        RECT 2366.770 48.180 2367.090 48.240 ;
        RECT 2366.770 48.040 2367.285 48.180 ;
        RECT 2366.770 47.980 2367.090 48.040 ;
        RECT 2366.785 2.960 2367.075 3.005 ;
        RECT 2369.530 2.960 2369.850 3.020 ;
        RECT 2366.785 2.820 2369.850 2.960 ;
        RECT 2366.785 2.775 2367.075 2.820 ;
        RECT 2369.530 2.760 2369.850 2.820 ;
      LAYER via ;
        RECT 747.140 1303.260 747.400 1303.520 ;
        RECT 751.740 1303.260 752.000 1303.520 ;
        RECT 751.740 79.600 752.000 79.860 ;
        RECT 2366.800 79.600 2367.060 79.860 ;
        RECT 2366.800 47.980 2367.060 48.240 ;
        RECT 2369.560 2.760 2369.820 3.020 ;
      LAYER met2 ;
        RECT 747.180 1323.135 747.460 1327.135 ;
        RECT 747.200 1303.550 747.340 1323.135 ;
        RECT 747.140 1303.230 747.400 1303.550 ;
        RECT 751.740 1303.230 752.000 1303.550 ;
        RECT 751.800 79.890 751.940 1303.230 ;
        RECT 751.740 79.570 752.000 79.890 ;
        RECT 2366.800 79.570 2367.060 79.890 ;
        RECT 2366.860 48.270 2367.000 79.570 ;
        RECT 2366.800 47.950 2367.060 48.270 ;
        RECT 2369.560 2.730 2369.820 3.050 ;
        RECT 2369.620 2.400 2369.760 2.730 ;
        RECT 2369.410 -4.800 2369.970 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1671.250 2389.760 1671.570 2389.820 ;
        RECT 2349.290 2389.760 2349.610 2389.820 ;
        RECT 1671.250 2389.620 2349.610 2389.760 ;
        RECT 1671.250 2389.560 1671.570 2389.620 ;
        RECT 2349.290 2389.560 2349.610 2389.620 ;
        RECT 2349.290 19.620 2349.610 19.680 ;
        RECT 2387.470 19.620 2387.790 19.680 ;
        RECT 2349.290 19.480 2387.790 19.620 ;
        RECT 2349.290 19.420 2349.610 19.480 ;
        RECT 2387.470 19.420 2387.790 19.480 ;
      LAYER via ;
        RECT 1671.280 2389.560 1671.540 2389.820 ;
        RECT 2349.320 2389.560 2349.580 2389.820 ;
        RECT 2349.320 19.420 2349.580 19.680 ;
        RECT 2387.500 19.420 2387.760 19.680 ;
      LAYER met2 ;
        RECT 1671.280 2389.530 1671.540 2389.850 ;
        RECT 2349.320 2389.530 2349.580 2389.850 ;
        RECT 1669.940 2377.690 1670.220 2377.880 ;
        RECT 1671.340 2377.690 1671.480 2389.530 ;
        RECT 1669.940 2377.550 1671.480 2377.690 ;
        RECT 1669.940 2373.880 1670.220 2377.550 ;
        RECT 2349.380 19.710 2349.520 2389.530 ;
        RECT 2349.320 19.390 2349.580 19.710 ;
        RECT 2387.500 19.390 2387.760 19.710 ;
        RECT 2387.560 2.400 2387.700 19.390 ;
        RECT 2387.350 -4.800 2387.910 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1652.005 2391.305 1653.555 2391.475 ;
        RECT 1652.005 2390.965 1652.175 2391.305 ;
        RECT 1653.385 2389.265 1653.555 2391.305 ;
      LAYER met1 ;
        RECT 1634.450 2391.120 1634.770 2391.180 ;
        RECT 1651.945 2391.120 1652.235 2391.165 ;
        RECT 1634.450 2390.980 1652.235 2391.120 ;
        RECT 1634.450 2390.920 1634.770 2390.980 ;
        RECT 1651.945 2390.935 1652.235 2390.980 ;
        RECT 1653.325 2389.420 1653.615 2389.465 ;
        RECT 2369.990 2389.420 2370.310 2389.480 ;
        RECT 1653.325 2389.280 2370.310 2389.420 ;
        RECT 1653.325 2389.235 1653.615 2389.280 ;
        RECT 2369.990 2389.220 2370.310 2389.280 ;
        RECT 2369.990 15.200 2370.310 15.260 ;
        RECT 2405.410 15.200 2405.730 15.260 ;
        RECT 2369.990 15.060 2405.730 15.200 ;
        RECT 2369.990 15.000 2370.310 15.060 ;
        RECT 2405.410 15.000 2405.730 15.060 ;
      LAYER via ;
        RECT 1634.480 2390.920 1634.740 2391.180 ;
        RECT 2370.020 2389.220 2370.280 2389.480 ;
        RECT 2370.020 15.000 2370.280 15.260 ;
        RECT 2405.440 15.000 2405.700 15.260 ;
      LAYER met2 ;
        RECT 1634.480 2390.890 1634.740 2391.210 ;
        RECT 1634.540 2377.690 1634.680 2390.890 ;
        RECT 2370.020 2389.190 2370.280 2389.510 ;
        RECT 1634.980 2377.690 1635.260 2377.880 ;
        RECT 1634.540 2377.550 1635.260 2377.690 ;
        RECT 1634.980 2373.880 1635.260 2377.550 ;
        RECT 2370.080 15.290 2370.220 2389.190 ;
        RECT 2370.020 14.970 2370.280 15.290 ;
        RECT 2405.440 14.970 2405.700 15.290 ;
        RECT 2405.500 2.400 2405.640 14.970 ;
        RECT 2405.290 -4.800 2405.850 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 703.410 2376.500 703.730 2376.560 ;
        RECT 765.970 2376.500 766.290 2376.560 ;
        RECT 703.410 2376.360 766.290 2376.500 ;
        RECT 703.410 2376.300 703.730 2376.360 ;
        RECT 765.970 2376.300 766.290 2376.360 ;
        RECT 703.410 14.520 703.730 14.580 ;
        RECT 799.550 14.520 799.870 14.580 ;
        RECT 703.410 14.380 799.870 14.520 ;
        RECT 703.410 14.320 703.730 14.380 ;
        RECT 799.550 14.320 799.870 14.380 ;
      LAYER via ;
        RECT 703.440 2376.300 703.700 2376.560 ;
        RECT 766.000 2376.300 766.260 2376.560 ;
        RECT 703.440 14.320 703.700 14.580 ;
        RECT 799.580 14.320 799.840 14.580 ;
      LAYER met2 ;
        RECT 703.440 2376.270 703.700 2376.590 ;
        RECT 766.000 2376.330 766.260 2376.590 ;
        RECT 767.420 2376.330 767.700 2377.880 ;
        RECT 766.000 2376.270 767.700 2376.330 ;
        RECT 703.500 1393.845 703.640 2376.270 ;
        RECT 766.060 2376.190 767.700 2376.270 ;
        RECT 767.420 2373.880 767.700 2376.190 ;
        RECT 703.430 1393.475 703.710 1393.845 ;
        RECT 703.430 1391.435 703.710 1391.805 ;
        RECT 703.500 14.610 703.640 1391.435 ;
        RECT 703.440 14.290 703.700 14.610 ;
        RECT 799.580 14.290 799.840 14.610 ;
        RECT 799.640 2.400 799.780 14.290 ;
        RECT 799.430 -4.800 799.990 2.400 ;
      LAYER via2 ;
        RECT 703.430 1393.520 703.710 1393.800 ;
        RECT 703.430 1391.480 703.710 1391.760 ;
      LAYER met3 ;
        RECT 703.405 1393.810 703.735 1393.825 ;
        RECT 703.190 1393.495 703.735 1393.810 ;
        RECT 703.190 1391.785 703.490 1393.495 ;
        RECT 703.190 1391.470 703.735 1391.785 ;
        RECT 703.405 1391.455 703.735 1391.470 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 648.210 2145.980 648.530 2146.040 ;
        RECT 704.330 2145.980 704.650 2146.040 ;
        RECT 648.210 2145.840 704.650 2145.980 ;
        RECT 648.210 2145.780 648.530 2145.840 ;
        RECT 704.330 2145.780 704.650 2145.840 ;
        RECT 644.990 17.240 645.310 17.300 ;
        RECT 648.210 17.240 648.530 17.300 ;
        RECT 644.990 17.100 648.530 17.240 ;
        RECT 644.990 17.040 645.310 17.100 ;
        RECT 648.210 17.040 648.530 17.100 ;
      LAYER via ;
        RECT 648.240 2145.780 648.500 2146.040 ;
        RECT 704.360 2145.780 704.620 2146.040 ;
        RECT 645.020 17.040 645.280 17.300 ;
        RECT 648.240 17.040 648.500 17.300 ;
      LAYER met2 ;
        RECT 704.350 2147.595 704.630 2147.965 ;
        RECT 704.420 2146.070 704.560 2147.595 ;
        RECT 648.240 2145.750 648.500 2146.070 ;
        RECT 704.360 2145.750 704.620 2146.070 ;
        RECT 648.300 17.330 648.440 2145.750 ;
        RECT 645.020 17.010 645.280 17.330 ;
        RECT 648.240 17.010 648.500 17.330 ;
        RECT 645.080 2.400 645.220 17.010 ;
        RECT 644.870 -4.800 645.430 2.400 ;
      LAYER via2 ;
        RECT 704.350 2147.640 704.630 2147.920 ;
      LAYER met3 ;
        RECT 704.325 2147.930 704.655 2147.945 ;
        RECT 715.810 2147.930 719.810 2147.935 ;
        RECT 704.325 2147.630 719.810 2147.930 ;
        RECT 704.325 2147.615 704.655 2147.630 ;
        RECT 715.810 2147.335 719.810 2147.630 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1771.070 2104.840 1771.390 2104.900 ;
        RECT 2391.150 2104.840 2391.470 2104.900 ;
        RECT 1771.070 2104.700 2391.470 2104.840 ;
        RECT 1771.070 2104.640 1771.390 2104.700 ;
        RECT 2391.150 2104.640 2391.470 2104.700 ;
        RECT 2391.150 19.280 2391.470 19.340 ;
        RECT 2428.870 19.280 2429.190 19.340 ;
        RECT 2391.150 19.140 2429.190 19.280 ;
        RECT 2391.150 19.080 2391.470 19.140 ;
        RECT 2428.870 19.080 2429.190 19.140 ;
      LAYER via ;
        RECT 1771.100 2104.640 1771.360 2104.900 ;
        RECT 2391.180 2104.640 2391.440 2104.900 ;
        RECT 2391.180 19.080 2391.440 19.340 ;
        RECT 2428.900 19.080 2429.160 19.340 ;
      LAYER met2 ;
        RECT 1771.090 2109.515 1771.370 2109.885 ;
        RECT 1771.160 2104.930 1771.300 2109.515 ;
        RECT 1771.100 2104.610 1771.360 2104.930 ;
        RECT 2391.180 2104.610 2391.440 2104.930 ;
        RECT 2391.240 19.370 2391.380 2104.610 ;
        RECT 2391.180 19.050 2391.440 19.370 ;
        RECT 2428.900 19.050 2429.160 19.370 ;
        RECT 2428.960 2.400 2429.100 19.050 ;
        RECT 2428.750 -4.800 2429.310 2.400 ;
      LAYER via2 ;
        RECT 1771.090 2109.560 1771.370 2109.840 ;
      LAYER met3 ;
        RECT 1755.835 2109.850 1759.835 2109.855 ;
        RECT 1771.065 2109.850 1771.395 2109.865 ;
        RECT 1755.835 2109.550 1771.395 2109.850 ;
        RECT 1755.835 2109.255 1759.835 2109.550 ;
        RECT 1771.065 2109.535 1771.395 2109.550 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1236.550 2393.160 1236.870 2393.220 ;
        RECT 2390.690 2393.160 2391.010 2393.220 ;
        RECT 1236.550 2393.020 2391.010 2393.160 ;
        RECT 1236.550 2392.960 1236.870 2393.020 ;
        RECT 2390.690 2392.960 2391.010 2393.020 ;
        RECT 2390.690 20.640 2391.010 20.700 ;
        RECT 2393.910 20.640 2394.230 20.700 ;
        RECT 2390.690 20.500 2394.230 20.640 ;
        RECT 2390.690 20.440 2391.010 20.500 ;
        RECT 2393.910 20.440 2394.230 20.500 ;
        RECT 2393.910 18.940 2394.230 19.000 ;
        RECT 2446.810 18.940 2447.130 19.000 ;
        RECT 2393.910 18.800 2447.130 18.940 ;
        RECT 2393.910 18.740 2394.230 18.800 ;
        RECT 2446.810 18.740 2447.130 18.800 ;
      LAYER via ;
        RECT 1236.580 2392.960 1236.840 2393.220 ;
        RECT 2390.720 2392.960 2390.980 2393.220 ;
        RECT 2390.720 20.440 2390.980 20.700 ;
        RECT 2393.940 20.440 2394.200 20.700 ;
        RECT 2393.940 18.740 2394.200 19.000 ;
        RECT 2446.840 18.740 2447.100 19.000 ;
      LAYER met2 ;
        RECT 1236.580 2392.930 1236.840 2393.250 ;
        RECT 2390.720 2392.930 2390.980 2393.250 ;
        RECT 1236.640 2377.880 1236.780 2392.930 ;
        RECT 1236.620 2373.880 1236.900 2377.880 ;
        RECT 2390.780 20.730 2390.920 2392.930 ;
        RECT 2390.720 20.410 2390.980 20.730 ;
        RECT 2393.940 20.410 2394.200 20.730 ;
        RECT 2394.000 19.030 2394.140 20.410 ;
        RECT 2393.940 18.710 2394.200 19.030 ;
        RECT 2446.840 18.710 2447.100 19.030 ;
        RECT 2446.900 2.400 2447.040 18.710 ;
        RECT 2446.690 -4.800 2447.250 2.400 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2404.490 1314.680 2404.810 1314.740 ;
        RECT 1083.460 1314.540 2404.810 1314.680 ;
        RECT 1076.470 1314.340 1076.790 1314.400 ;
        RECT 1083.460 1314.340 1083.600 1314.540 ;
        RECT 2404.490 1314.480 2404.810 1314.540 ;
        RECT 1076.470 1314.200 1083.600 1314.340 ;
        RECT 1076.470 1314.140 1076.790 1314.200 ;
        RECT 2404.490 17.920 2404.810 17.980 ;
        RECT 2464.750 17.920 2465.070 17.980 ;
        RECT 2404.490 17.780 2465.070 17.920 ;
        RECT 2404.490 17.720 2404.810 17.780 ;
        RECT 2464.750 17.720 2465.070 17.780 ;
      LAYER via ;
        RECT 1076.500 1314.140 1076.760 1314.400 ;
        RECT 2404.520 1314.480 2404.780 1314.740 ;
        RECT 2404.520 17.720 2404.780 17.980 ;
        RECT 2464.780 17.720 2465.040 17.980 ;
      LAYER met2 ;
        RECT 1076.540 1323.135 1076.820 1327.135 ;
        RECT 1076.560 1314.430 1076.700 1323.135 ;
        RECT 2404.520 1314.450 2404.780 1314.770 ;
        RECT 1076.500 1314.110 1076.760 1314.430 ;
        RECT 2404.580 18.010 2404.720 1314.450 ;
        RECT 2404.520 17.690 2404.780 18.010 ;
        RECT 2464.780 17.690 2465.040 18.010 ;
        RECT 2464.840 2.400 2464.980 17.690 ;
        RECT 2464.630 -4.800 2465.190 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1105.910 1314.340 1106.230 1314.400 ;
        RECT 2432.090 1314.340 2432.410 1314.400 ;
        RECT 1105.910 1314.200 2432.410 1314.340 ;
        RECT 1105.910 1314.140 1106.230 1314.200 ;
        RECT 2432.090 1314.140 2432.410 1314.200 ;
        RECT 2432.090 19.620 2432.410 19.680 ;
        RECT 2432.090 19.480 2447.960 19.620 ;
        RECT 2432.090 19.420 2432.410 19.480 ;
        RECT 2447.820 19.280 2447.960 19.480 ;
        RECT 2482.690 19.280 2483.010 19.340 ;
        RECT 2447.820 19.140 2483.010 19.280 ;
        RECT 2482.690 19.080 2483.010 19.140 ;
      LAYER via ;
        RECT 1105.940 1314.140 1106.200 1314.400 ;
        RECT 2432.120 1314.140 2432.380 1314.400 ;
        RECT 2432.120 19.420 2432.380 19.680 ;
        RECT 2482.720 19.080 2482.980 19.340 ;
      LAYER met2 ;
        RECT 1105.980 1323.135 1106.260 1327.135 ;
        RECT 1106.000 1314.430 1106.140 1323.135 ;
        RECT 1105.940 1314.110 1106.200 1314.430 ;
        RECT 2432.120 1314.110 2432.380 1314.430 ;
        RECT 2432.180 19.710 2432.320 1314.110 ;
        RECT 2432.120 19.390 2432.380 19.710 ;
        RECT 2482.720 19.050 2482.980 19.370 ;
        RECT 2482.780 2.400 2482.920 19.050 ;
        RECT 2482.570 -4.800 2483.130 2.400 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1768.310 1890.980 1768.630 1891.040 ;
        RECT 2438.990 1890.980 2439.310 1891.040 ;
        RECT 1768.310 1890.840 2439.310 1890.980 ;
        RECT 1768.310 1890.780 1768.630 1890.840 ;
        RECT 2438.990 1890.780 2439.310 1890.840 ;
        RECT 2438.990 19.960 2439.310 20.020 ;
        RECT 2500.630 19.960 2500.950 20.020 ;
        RECT 2438.990 19.820 2500.950 19.960 ;
        RECT 2438.990 19.760 2439.310 19.820 ;
        RECT 2500.630 19.760 2500.950 19.820 ;
      LAYER via ;
        RECT 1768.340 1890.780 1768.600 1891.040 ;
        RECT 2439.020 1890.780 2439.280 1891.040 ;
        RECT 2439.020 19.760 2439.280 20.020 ;
        RECT 2500.660 19.760 2500.920 20.020 ;
      LAYER met2 ;
        RECT 1768.330 1894.635 1768.610 1895.005 ;
        RECT 1768.400 1891.070 1768.540 1894.635 ;
        RECT 1768.340 1890.750 1768.600 1891.070 ;
        RECT 2439.020 1890.750 2439.280 1891.070 ;
        RECT 2439.080 20.050 2439.220 1890.750 ;
        RECT 2439.020 19.730 2439.280 20.050 ;
        RECT 2500.660 19.730 2500.920 20.050 ;
        RECT 2500.720 2.400 2500.860 19.730 ;
        RECT 2500.510 -4.800 2501.070 2.400 ;
      LAYER via2 ;
        RECT 1768.330 1894.680 1768.610 1894.960 ;
      LAYER met3 ;
        RECT 1755.835 1894.970 1759.835 1894.975 ;
        RECT 1768.305 1894.970 1768.635 1894.985 ;
        RECT 1755.835 1894.670 1768.635 1894.970 ;
        RECT 1755.835 1894.375 1759.835 1894.670 ;
        RECT 1768.305 1894.655 1768.635 1894.670 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1772.910 1732.200 1773.230 1732.260 ;
        RECT 2445.890 1732.200 2446.210 1732.260 ;
        RECT 1772.910 1732.060 2446.210 1732.200 ;
        RECT 1772.910 1732.000 1773.230 1732.060 ;
        RECT 2445.890 1732.000 2446.210 1732.060 ;
        RECT 2445.890 19.280 2446.210 19.340 ;
        RECT 2445.890 19.140 2447.500 19.280 ;
        RECT 2445.890 19.080 2446.210 19.140 ;
        RECT 2447.360 18.940 2447.500 19.140 ;
        RECT 2518.110 18.940 2518.430 19.000 ;
        RECT 2447.360 18.800 2518.430 18.940 ;
        RECT 2518.110 18.740 2518.430 18.800 ;
      LAYER via ;
        RECT 1772.940 1732.000 1773.200 1732.260 ;
        RECT 2445.920 1732.000 2446.180 1732.260 ;
        RECT 2445.920 19.080 2446.180 19.340 ;
        RECT 2518.140 18.740 2518.400 19.000 ;
      LAYER met2 ;
        RECT 1772.930 1732.795 1773.210 1733.165 ;
        RECT 1773.000 1732.290 1773.140 1732.795 ;
        RECT 1772.940 1731.970 1773.200 1732.290 ;
        RECT 2445.920 1731.970 2446.180 1732.290 ;
        RECT 2445.980 19.370 2446.120 1731.970 ;
        RECT 2445.920 19.050 2446.180 19.370 ;
        RECT 2518.140 18.710 2518.400 19.030 ;
        RECT 2518.200 2.400 2518.340 18.710 ;
        RECT 2517.990 -4.800 2518.550 2.400 ;
      LAYER via2 ;
        RECT 1772.930 1732.840 1773.210 1733.120 ;
      LAYER met3 ;
        RECT 1755.835 1733.130 1759.835 1733.135 ;
        RECT 1772.905 1733.130 1773.235 1733.145 ;
        RECT 1755.835 1732.830 1773.235 1733.130 ;
        RECT 1755.835 1732.535 1759.835 1732.830 ;
        RECT 1772.905 1732.815 1773.235 1732.830 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 752.630 1311.620 752.950 1311.680 ;
        RECT 758.150 1311.620 758.470 1311.680 ;
        RECT 752.630 1311.480 758.470 1311.620 ;
        RECT 752.630 1311.420 752.950 1311.480 ;
        RECT 758.150 1311.420 758.470 1311.480 ;
        RECT 758.150 79.460 758.470 79.520 ;
        RECT 2532.370 79.460 2532.690 79.520 ;
        RECT 758.150 79.320 2532.690 79.460 ;
        RECT 758.150 79.260 758.470 79.320 ;
        RECT 2532.370 79.260 2532.690 79.320 ;
        RECT 2532.370 62.120 2532.690 62.180 ;
        RECT 2536.050 62.120 2536.370 62.180 ;
        RECT 2532.370 61.980 2536.370 62.120 ;
        RECT 2532.370 61.920 2532.690 61.980 ;
        RECT 2536.050 61.920 2536.370 61.980 ;
      LAYER via ;
        RECT 752.660 1311.420 752.920 1311.680 ;
        RECT 758.180 1311.420 758.440 1311.680 ;
        RECT 758.180 79.260 758.440 79.520 ;
        RECT 2532.400 79.260 2532.660 79.520 ;
        RECT 2532.400 61.920 2532.660 62.180 ;
        RECT 2536.080 61.920 2536.340 62.180 ;
      LAYER met2 ;
        RECT 752.700 1323.135 752.980 1327.135 ;
        RECT 752.720 1311.710 752.860 1323.135 ;
        RECT 752.660 1311.390 752.920 1311.710 ;
        RECT 758.180 1311.390 758.440 1311.710 ;
        RECT 758.240 821.965 758.380 1311.390 ;
        RECT 758.170 821.595 758.450 821.965 ;
        RECT 758.170 820.915 758.450 821.285 ;
        RECT 758.240 79.550 758.380 820.915 ;
        RECT 758.180 79.230 758.440 79.550 ;
        RECT 2532.400 79.230 2532.660 79.550 ;
        RECT 2532.460 62.210 2532.600 79.230 ;
        RECT 2532.400 61.890 2532.660 62.210 ;
        RECT 2536.080 61.890 2536.340 62.210 ;
        RECT 2536.140 2.400 2536.280 61.890 ;
        RECT 2535.930 -4.800 2536.490 2.400 ;
      LAYER via2 ;
        RECT 758.170 821.640 758.450 821.920 ;
        RECT 758.170 820.960 758.450 821.240 ;
      LAYER met3 ;
        RECT 758.145 821.930 758.475 821.945 ;
        RECT 758.145 821.615 758.690 821.930 ;
        RECT 758.390 821.265 758.690 821.615 ;
        RECT 758.145 820.950 758.690 821.265 ;
        RECT 758.145 820.935 758.475 820.950 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1163.870 1315.020 1164.190 1315.080 ;
        RECT 2480.390 1315.020 2480.710 1315.080 ;
        RECT 1163.870 1314.880 2480.710 1315.020 ;
        RECT 1163.870 1314.820 1164.190 1314.880 ;
        RECT 2480.390 1314.820 2480.710 1314.880 ;
        RECT 2480.390 19.620 2480.710 19.680 ;
        RECT 2480.390 19.480 2483.380 19.620 ;
        RECT 2480.390 19.420 2480.710 19.480 ;
        RECT 2483.240 19.280 2483.380 19.480 ;
        RECT 2553.990 19.280 2554.310 19.340 ;
        RECT 2483.240 19.140 2554.310 19.280 ;
        RECT 2553.990 19.080 2554.310 19.140 ;
      LAYER via ;
        RECT 1163.900 1314.820 1164.160 1315.080 ;
        RECT 2480.420 1314.820 2480.680 1315.080 ;
        RECT 2480.420 19.420 2480.680 19.680 ;
        RECT 2554.020 19.080 2554.280 19.340 ;
      LAYER met2 ;
        RECT 1163.940 1323.135 1164.220 1327.135 ;
        RECT 1163.960 1315.110 1164.100 1323.135 ;
        RECT 1163.900 1314.790 1164.160 1315.110 ;
        RECT 2480.420 1314.790 2480.680 1315.110 ;
        RECT 2480.480 19.710 2480.620 1314.790 ;
        RECT 2480.420 19.390 2480.680 19.710 ;
        RECT 2554.020 19.050 2554.280 19.370 ;
        RECT 2554.080 2.400 2554.220 19.050 ;
        RECT 2553.870 -4.800 2554.430 2.400 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1772.910 2159.920 1773.230 2159.980 ;
        RECT 2494.190 2159.920 2494.510 2159.980 ;
        RECT 1772.910 2159.780 2494.510 2159.920 ;
        RECT 1772.910 2159.720 1773.230 2159.780 ;
        RECT 2494.190 2159.720 2494.510 2159.780 ;
        RECT 2495.110 19.620 2495.430 19.680 ;
        RECT 2571.930 19.620 2572.250 19.680 ;
        RECT 2495.110 19.480 2572.250 19.620 ;
        RECT 2495.110 19.420 2495.430 19.480 ;
        RECT 2571.930 19.420 2572.250 19.480 ;
      LAYER via ;
        RECT 1772.940 2159.720 1773.200 2159.980 ;
        RECT 2494.220 2159.720 2494.480 2159.980 ;
        RECT 2495.140 19.420 2495.400 19.680 ;
        RECT 2571.960 19.420 2572.220 19.680 ;
      LAYER met2 ;
        RECT 1772.930 2159.835 1773.210 2160.205 ;
        RECT 1772.940 2159.690 1773.200 2159.835 ;
        RECT 2494.220 2159.690 2494.480 2160.010 ;
        RECT 2494.280 33.730 2494.420 2159.690 ;
        RECT 2494.280 33.590 2495.340 33.730 ;
        RECT 2495.200 19.710 2495.340 33.590 ;
        RECT 2495.140 19.390 2495.400 19.710 ;
        RECT 2571.960 19.390 2572.220 19.710 ;
        RECT 2572.020 2.400 2572.160 19.390 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
      LAYER via2 ;
        RECT 1772.930 2159.880 1773.210 2160.160 ;
      LAYER met3 ;
        RECT 1755.835 2160.170 1759.835 2160.175 ;
        RECT 1772.905 2160.170 1773.235 2160.185 ;
        RECT 1755.835 2159.870 1773.235 2160.170 ;
        RECT 1755.835 2159.575 1759.835 2159.870 ;
        RECT 1772.905 2159.855 1773.235 2159.870 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2501.090 17.920 2501.410 17.980 ;
        RECT 2589.410 17.920 2589.730 17.980 ;
        RECT 2501.090 17.780 2589.730 17.920 ;
        RECT 2501.090 17.720 2501.410 17.780 ;
        RECT 2589.410 17.720 2589.730 17.780 ;
      LAYER via ;
        RECT 2501.120 17.720 2501.380 17.980 ;
        RECT 2589.440 17.720 2589.700 17.980 ;
      LAYER met2 ;
        RECT 1184.130 2388.315 1184.410 2388.685 ;
        RECT 2501.110 2388.315 2501.390 2388.685 ;
        RECT 1184.200 2377.880 1184.340 2388.315 ;
        RECT 1184.180 2373.880 1184.460 2377.880 ;
        RECT 2501.180 18.010 2501.320 2388.315 ;
        RECT 2501.120 17.690 2501.380 18.010 ;
        RECT 2589.440 17.690 2589.700 18.010 ;
        RECT 2589.500 2.400 2589.640 17.690 ;
        RECT 2589.290 -4.800 2589.850 2.400 ;
      LAYER via2 ;
        RECT 1184.130 2388.360 1184.410 2388.640 ;
        RECT 2501.110 2388.360 2501.390 2388.640 ;
      LAYER met3 ;
        RECT 1184.105 2388.650 1184.435 2388.665 ;
        RECT 2501.085 2388.650 2501.415 2388.665 ;
        RECT 1184.105 2388.350 2501.415 2388.650 ;
        RECT 1184.105 2388.335 1184.435 2388.350 ;
        RECT 2501.085 2388.335 2501.415 2388.350 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 823.490 59.315 823.770 59.685 ;
        RECT 823.560 2.400 823.700 59.315 ;
        RECT 823.350 -4.800 823.910 2.400 ;
      LAYER via2 ;
        RECT 823.490 59.360 823.770 59.640 ;
      LAYER met3 ;
        RECT 1755.835 1990.170 1759.835 1990.175 ;
        RECT 1767.590 1990.170 1767.970 1990.180 ;
        RECT 1755.835 1989.870 1767.970 1990.170 ;
        RECT 1755.835 1989.575 1759.835 1989.870 ;
        RECT 1767.590 1989.860 1767.970 1989.870 ;
        RECT 823.465 59.650 823.795 59.665 ;
        RECT 1767.590 59.650 1767.970 59.660 ;
        RECT 823.465 59.350 1767.970 59.650 ;
        RECT 823.465 59.335 823.795 59.350 ;
        RECT 1767.590 59.340 1767.970 59.350 ;
      LAYER via3 ;
        RECT 1767.620 1989.860 1767.940 1990.180 ;
        RECT 1767.620 59.340 1767.940 59.660 ;
      LAYER met4 ;
        RECT 1767.615 1989.855 1767.945 1990.185 ;
        RECT 1767.630 59.665 1767.930 1989.855 ;
        RECT 1767.615 59.335 1767.945 59.665 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2518.645 18.785 2518.815 19.975 ;
      LAYER mcon ;
        RECT 2518.645 19.805 2518.815 19.975 ;
      LAYER met1 ;
        RECT 2515.350 19.960 2515.670 20.020 ;
        RECT 2518.585 19.960 2518.875 20.005 ;
        RECT 2515.350 19.820 2518.875 19.960 ;
        RECT 2515.350 19.760 2515.670 19.820 ;
        RECT 2518.585 19.775 2518.875 19.820 ;
        RECT 2518.585 18.940 2518.875 18.985 ;
        RECT 2607.350 18.940 2607.670 19.000 ;
        RECT 2518.585 18.800 2607.670 18.940 ;
        RECT 2518.585 18.755 2518.875 18.800 ;
        RECT 2607.350 18.740 2607.670 18.800 ;
      LAYER via ;
        RECT 2515.380 19.760 2515.640 20.020 ;
        RECT 2607.380 18.740 2607.640 19.000 ;
      LAYER met2 ;
        RECT 1189.650 2387.635 1189.930 2388.005 ;
        RECT 2515.370 2387.635 2515.650 2388.005 ;
        RECT 1189.720 2377.880 1189.860 2387.635 ;
        RECT 1189.700 2373.880 1189.980 2377.880 ;
        RECT 2515.440 20.050 2515.580 2387.635 ;
        RECT 2515.380 19.730 2515.640 20.050 ;
        RECT 2607.380 18.710 2607.640 19.030 ;
        RECT 2607.440 2.400 2607.580 18.710 ;
        RECT 2607.230 -4.800 2607.790 2.400 ;
      LAYER via2 ;
        RECT 1189.650 2387.680 1189.930 2387.960 ;
        RECT 2515.370 2387.680 2515.650 2387.960 ;
      LAYER met3 ;
        RECT 1189.625 2387.970 1189.955 2387.985 ;
        RECT 2515.345 2387.970 2515.675 2387.985 ;
        RECT 1189.625 2387.670 2515.675 2387.970 ;
        RECT 1189.625 2387.655 1189.955 2387.670 ;
        RECT 2515.345 2387.655 2515.675 2387.670 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1444.470 2393.500 1444.790 2393.560 ;
        RECT 2514.890 2393.500 2515.210 2393.560 ;
        RECT 1444.470 2393.360 2515.210 2393.500 ;
        RECT 1444.470 2393.300 1444.790 2393.360 ;
        RECT 2514.890 2393.300 2515.210 2393.360 ;
        RECT 2514.890 20.640 2515.210 20.700 ;
        RECT 2625.290 20.640 2625.610 20.700 ;
        RECT 2514.890 20.500 2625.610 20.640 ;
        RECT 2514.890 20.440 2515.210 20.500 ;
        RECT 2625.290 20.440 2625.610 20.500 ;
      LAYER via ;
        RECT 1444.500 2393.300 1444.760 2393.560 ;
        RECT 2514.920 2393.300 2515.180 2393.560 ;
        RECT 2514.920 20.440 2515.180 20.700 ;
        RECT 2625.320 20.440 2625.580 20.700 ;
      LAYER met2 ;
        RECT 1444.500 2393.270 1444.760 2393.590 ;
        RECT 2514.920 2393.270 2515.180 2393.590 ;
        RECT 1444.560 2377.880 1444.700 2393.270 ;
        RECT 1444.540 2373.880 1444.820 2377.880 ;
        RECT 2514.980 20.730 2515.120 2393.270 ;
        RECT 2514.920 20.410 2515.180 20.730 ;
        RECT 2625.320 20.410 2625.580 20.730 ;
        RECT 2625.380 2.400 2625.520 20.410 ;
        RECT 2625.170 -4.800 2625.730 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1400.310 31.860 1400.630 31.920 ;
        RECT 2643.230 31.860 2643.550 31.920 ;
        RECT 1400.310 31.720 2643.550 31.860 ;
        RECT 1400.310 31.660 1400.630 31.720 ;
        RECT 2643.230 31.660 2643.550 31.720 ;
      LAYER via ;
        RECT 1400.340 31.660 1400.600 31.920 ;
        RECT 2643.260 31.660 2643.520 31.920 ;
      LAYER met2 ;
        RECT 1400.380 1323.135 1400.660 1327.135 ;
        RECT 1400.400 31.950 1400.540 1323.135 ;
        RECT 1400.340 31.630 1400.600 31.950 ;
        RECT 2643.260 31.630 2643.520 31.950 ;
        RECT 2643.320 2.400 2643.460 31.630 ;
        RECT 2643.110 -4.800 2643.670 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1186.870 1311.280 1187.190 1311.340 ;
        RECT 1193.310 1311.280 1193.630 1311.340 ;
        RECT 1186.870 1311.140 1193.630 1311.280 ;
        RECT 1186.870 1311.080 1187.190 1311.140 ;
        RECT 1193.310 1311.080 1193.630 1311.140 ;
        RECT 1193.310 31.180 1193.630 31.240 ;
        RECT 2661.170 31.180 2661.490 31.240 ;
        RECT 1193.310 31.040 2661.490 31.180 ;
        RECT 1193.310 30.980 1193.630 31.040 ;
        RECT 2661.170 30.980 2661.490 31.040 ;
      LAYER via ;
        RECT 1186.900 1311.080 1187.160 1311.340 ;
        RECT 1193.340 1311.080 1193.600 1311.340 ;
        RECT 1193.340 30.980 1193.600 31.240 ;
        RECT 2661.200 30.980 2661.460 31.240 ;
      LAYER met2 ;
        RECT 1186.940 1323.135 1187.220 1327.135 ;
        RECT 1186.960 1311.370 1187.100 1323.135 ;
        RECT 1186.900 1311.050 1187.160 1311.370 ;
        RECT 1193.340 1311.050 1193.600 1311.370 ;
        RECT 1193.400 31.270 1193.540 1311.050 ;
        RECT 1193.340 30.950 1193.600 31.270 ;
        RECT 2661.200 30.950 2661.460 31.270 ;
        RECT 2661.260 2.400 2661.400 30.950 ;
        RECT 2661.050 -4.800 2661.610 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 717.285 1504.585 717.455 1562.215 ;
        RECT 711.765 1431.485 711.935 1498.975 ;
      LAYER mcon ;
        RECT 717.285 1562.045 717.455 1562.215 ;
        RECT 711.765 1498.805 711.935 1498.975 ;
      LAYER met1 ;
        RECT 717.670 2192.220 717.990 2192.280 ;
        RECT 719.510 2192.220 719.830 2192.280 ;
        RECT 717.670 2192.080 719.830 2192.220 ;
        RECT 717.670 2192.020 717.990 2192.080 ;
        RECT 719.510 2192.020 719.830 2192.080 ;
        RECT 717.670 2152.780 717.990 2152.840 ;
        RECT 719.510 2152.780 719.830 2152.840 ;
        RECT 717.670 2152.640 719.830 2152.780 ;
        RECT 717.670 2152.580 717.990 2152.640 ;
        RECT 719.510 2152.580 719.830 2152.640 ;
        RECT 717.210 1562.200 717.530 1562.260 ;
        RECT 717.015 1562.060 717.530 1562.200 ;
        RECT 717.210 1562.000 717.530 1562.060 ;
        RECT 717.210 1504.740 717.530 1504.800 ;
        RECT 717.015 1504.600 717.530 1504.740 ;
        RECT 717.210 1504.540 717.530 1504.600 ;
        RECT 711.690 1498.960 712.010 1499.020 ;
        RECT 711.495 1498.820 712.010 1498.960 ;
        RECT 711.690 1498.760 712.010 1498.820 ;
        RECT 711.705 1431.640 711.995 1431.685 ;
        RECT 717.210 1431.640 717.530 1431.700 ;
        RECT 711.705 1431.500 717.530 1431.640 ;
        RECT 711.705 1431.455 711.995 1431.500 ;
        RECT 717.210 1431.440 717.530 1431.500 ;
      LAYER via ;
        RECT 717.700 2192.020 717.960 2192.280 ;
        RECT 719.540 2192.020 719.800 2192.280 ;
        RECT 717.700 2152.580 717.960 2152.840 ;
        RECT 719.540 2152.580 719.800 2152.840 ;
        RECT 717.240 1562.000 717.500 1562.260 ;
        RECT 717.240 1504.540 717.500 1504.800 ;
        RECT 711.720 1498.760 711.980 1499.020 ;
        RECT 717.240 1431.440 717.500 1431.700 ;
      LAYER met2 ;
        RECT 718.150 2308.075 718.430 2308.445 ;
        RECT 718.220 2245.885 718.360 2308.075 ;
        RECT 718.150 2245.515 718.430 2245.885 ;
        RECT 717.690 2211.515 717.970 2211.885 ;
        RECT 717.760 2192.310 717.900 2211.515 ;
        RECT 717.700 2191.990 717.960 2192.310 ;
        RECT 719.540 2191.990 719.800 2192.310 ;
        RECT 719.600 2152.870 719.740 2191.990 ;
        RECT 717.700 2152.550 717.960 2152.870 ;
        RECT 719.540 2152.550 719.800 2152.870 ;
        RECT 717.760 2127.450 717.900 2152.550 ;
        RECT 717.760 2127.310 718.360 2127.450 ;
        RECT 718.220 2086.085 718.360 2127.310 ;
        RECT 718.150 2085.715 718.430 2086.085 ;
        RECT 718.610 2052.395 718.890 2052.765 ;
        RECT 718.680 2005.845 718.820 2052.395 ;
        RECT 718.610 2005.475 718.890 2005.845 ;
        RECT 713.550 1963.315 713.830 1963.685 ;
        RECT 713.620 1938.525 713.760 1963.315 ;
        RECT 713.550 1938.155 713.830 1938.525 ;
        RECT 718.610 1579.115 718.890 1579.485 ;
        RECT 718.680 1573.365 718.820 1579.115 ;
        RECT 718.610 1572.995 718.890 1573.365 ;
        RECT 717.230 1562.115 717.510 1562.485 ;
        RECT 717.240 1561.970 717.500 1562.115 ;
        RECT 717.240 1504.685 717.500 1504.830 ;
        RECT 717.230 1504.315 717.510 1504.685 ;
        RECT 711.710 1498.875 711.990 1499.245 ;
        RECT 711.720 1498.730 711.980 1498.875 ;
        RECT 717.240 1431.410 717.500 1431.730 ;
        RECT 717.300 1431.245 717.440 1431.410 ;
        RECT 717.230 1430.875 717.510 1431.245 ;
        RECT 717.690 516.955 717.970 517.325 ;
        RECT 717.760 475.845 717.900 516.955 ;
        RECT 717.690 475.475 717.970 475.845 ;
        RECT 2678.670 57.955 2678.950 58.325 ;
        RECT 2678.740 2.400 2678.880 57.955 ;
        RECT 2678.530 -4.800 2679.090 2.400 ;
      LAYER via2 ;
        RECT 718.150 2308.120 718.430 2308.400 ;
        RECT 718.150 2245.560 718.430 2245.840 ;
        RECT 717.690 2211.560 717.970 2211.840 ;
        RECT 718.150 2085.760 718.430 2086.040 ;
        RECT 718.610 2052.440 718.890 2052.720 ;
        RECT 718.610 2005.520 718.890 2005.800 ;
        RECT 713.550 1963.360 713.830 1963.640 ;
        RECT 713.550 1938.200 713.830 1938.480 ;
        RECT 718.610 1579.160 718.890 1579.440 ;
        RECT 718.610 1573.040 718.890 1573.320 ;
        RECT 717.230 1562.160 717.510 1562.440 ;
        RECT 717.230 1504.360 717.510 1504.640 ;
        RECT 711.710 1498.920 711.990 1499.200 ;
        RECT 717.230 1430.920 717.510 1431.200 ;
        RECT 717.690 517.000 717.970 517.280 ;
        RECT 717.690 475.520 717.970 475.800 ;
        RECT 2678.670 58.000 2678.950 58.280 ;
      LAYER met3 ;
        RECT 715.810 2310.535 719.810 2311.135 ;
        RECT 717.910 2308.425 718.210 2310.535 ;
        RECT 717.910 2308.110 718.455 2308.425 ;
        RECT 718.125 2308.095 718.455 2308.110 ;
        RECT 718.125 2245.860 718.455 2245.865 ;
        RECT 717.870 2245.850 718.455 2245.860 ;
        RECT 717.670 2245.550 718.455 2245.850 ;
        RECT 717.870 2245.540 718.455 2245.550 ;
        RECT 718.125 2245.535 718.455 2245.540 ;
        RECT 717.665 2211.860 717.995 2211.865 ;
        RECT 717.665 2211.850 718.250 2211.860 ;
        RECT 717.665 2211.550 718.450 2211.850 ;
        RECT 717.665 2211.540 718.250 2211.550 ;
        RECT 717.665 2211.535 717.995 2211.540 ;
        RECT 718.125 2086.050 718.455 2086.065 ;
        RECT 718.790 2086.050 719.170 2086.060 ;
        RECT 718.125 2085.750 719.170 2086.050 ;
        RECT 718.125 2085.735 718.455 2085.750 ;
        RECT 718.790 2085.740 719.170 2085.750 ;
        RECT 718.585 2052.740 718.915 2052.745 ;
        RECT 718.585 2052.730 719.170 2052.740 ;
        RECT 718.360 2052.430 719.170 2052.730 ;
        RECT 718.585 2052.420 719.170 2052.430 ;
        RECT 718.585 2052.415 718.915 2052.420 ;
        RECT 716.030 2005.810 716.410 2005.820 ;
        RECT 718.585 2005.810 718.915 2005.825 ;
        RECT 716.030 2005.510 718.915 2005.810 ;
        RECT 716.030 2005.500 716.410 2005.510 ;
        RECT 718.585 2005.495 718.915 2005.510 ;
        RECT 713.525 1963.650 713.855 1963.665 ;
        RECT 716.030 1963.650 716.410 1963.660 ;
        RECT 713.525 1963.350 716.410 1963.650 ;
        RECT 713.525 1963.335 713.855 1963.350 ;
        RECT 716.030 1963.340 716.410 1963.350 ;
        RECT 713.525 1938.490 713.855 1938.505 ;
        RECT 717.870 1938.490 718.250 1938.500 ;
        RECT 713.525 1938.190 718.250 1938.490 ;
        RECT 713.525 1938.175 713.855 1938.190 ;
        RECT 717.870 1938.180 718.250 1938.190 ;
        RECT 717.870 1917.780 718.250 1918.100 ;
        RECT 717.910 1917.420 718.210 1917.780 ;
        RECT 717.640 1917.110 718.210 1917.420 ;
        RECT 717.640 1917.100 718.020 1917.110 ;
        RECT 716.030 1816.770 716.410 1816.780 ;
        RECT 716.030 1816.470 718.210 1816.770 ;
        RECT 716.030 1816.460 716.410 1816.470 ;
        RECT 717.910 1815.410 718.210 1816.470 ;
        RECT 718.790 1815.410 719.170 1815.420 ;
        RECT 717.910 1815.110 719.170 1815.410 ;
        RECT 718.790 1815.100 719.170 1815.110 ;
        RECT 716.030 1811.330 716.410 1811.340 ;
        RECT 718.790 1811.330 719.170 1811.340 ;
        RECT 716.030 1811.030 719.170 1811.330 ;
        RECT 716.030 1811.020 716.410 1811.030 ;
        RECT 718.790 1811.020 719.170 1811.030 ;
        RECT 716.030 1625.690 716.410 1625.700 ;
        RECT 718.790 1625.690 719.170 1625.700 ;
        RECT 716.030 1625.390 719.170 1625.690 ;
        RECT 716.030 1625.380 716.410 1625.390 ;
        RECT 718.790 1625.380 719.170 1625.390 ;
        RECT 718.585 1579.460 718.915 1579.465 ;
        RECT 718.585 1579.450 719.170 1579.460 ;
        RECT 718.585 1579.150 719.370 1579.450 ;
        RECT 718.585 1579.140 719.170 1579.150 ;
        RECT 718.585 1579.135 718.915 1579.140 ;
        RECT 718.585 1573.330 718.915 1573.345 ;
        RECT 717.910 1573.030 718.915 1573.330 ;
        RECT 717.910 1571.970 718.210 1573.030 ;
        RECT 718.585 1573.015 718.915 1573.030 ;
        RECT 718.790 1571.970 719.170 1571.980 ;
        RECT 717.910 1571.670 719.170 1571.970 ;
        RECT 718.790 1571.660 719.170 1571.670 ;
        RECT 717.205 1562.450 717.535 1562.465 ;
        RECT 718.790 1562.450 719.170 1562.460 ;
        RECT 717.205 1562.150 719.170 1562.450 ;
        RECT 717.205 1562.135 717.535 1562.150 ;
        RECT 718.790 1562.140 719.170 1562.150 ;
        RECT 717.205 1504.650 717.535 1504.665 ;
        RECT 718.790 1504.650 719.170 1504.660 ;
        RECT 717.205 1504.350 719.170 1504.650 ;
        RECT 717.205 1504.335 717.535 1504.350 ;
        RECT 718.790 1504.340 719.170 1504.350 ;
        RECT 711.685 1499.210 712.015 1499.225 ;
        RECT 718.790 1499.210 719.170 1499.220 ;
        RECT 711.685 1498.910 719.170 1499.210 ;
        RECT 711.685 1498.895 712.015 1498.910 ;
        RECT 718.790 1498.900 719.170 1498.910 ;
        RECT 715.110 1431.210 715.490 1431.220 ;
        RECT 717.205 1431.210 717.535 1431.225 ;
        RECT 715.110 1430.910 717.535 1431.210 ;
        RECT 715.110 1430.900 715.490 1430.910 ;
        RECT 717.205 1430.895 717.535 1430.910 ;
        RECT 715.110 1403.330 715.490 1403.340 ;
        RECT 714.230 1403.030 715.490 1403.330 ;
        RECT 714.230 1401.970 714.530 1403.030 ;
        RECT 715.110 1403.020 715.490 1403.030 ;
        RECT 716.950 1401.970 717.330 1401.980 ;
        RECT 714.230 1401.670 717.330 1401.970 ;
        RECT 716.950 1401.660 717.330 1401.670 ;
        RECT 716.950 1355.730 717.330 1355.740 ;
        RECT 715.150 1355.430 717.330 1355.730 ;
        RECT 715.150 1350.290 715.450 1355.430 ;
        RECT 716.950 1355.420 717.330 1355.430 ;
        RECT 715.150 1349.990 716.370 1350.290 ;
        RECT 716.070 1347.570 716.370 1349.990 ;
        RECT 718.790 1347.570 719.170 1347.580 ;
        RECT 716.070 1347.270 719.170 1347.570 ;
        RECT 718.790 1347.260 719.170 1347.270 ;
        RECT 717.870 1321.730 718.250 1321.740 ;
        RECT 720.630 1321.730 721.010 1321.740 ;
        RECT 717.870 1321.430 721.010 1321.730 ;
        RECT 717.870 1321.420 718.250 1321.430 ;
        RECT 720.630 1321.420 721.010 1321.430 ;
        RECT 717.870 1210.890 718.250 1210.900 ;
        RECT 720.630 1210.890 721.010 1210.900 ;
        RECT 717.870 1210.590 721.010 1210.890 ;
        RECT 717.870 1210.580 718.250 1210.590 ;
        RECT 720.630 1210.580 721.010 1210.590 ;
        RECT 717.870 1052.450 718.250 1052.460 ;
        RECT 720.630 1052.450 721.010 1052.460 ;
        RECT 717.870 1052.150 721.010 1052.450 ;
        RECT 717.870 1052.140 718.250 1052.150 ;
        RECT 720.630 1052.140 721.010 1052.150 ;
        RECT 717.870 1017.770 718.250 1017.780 ;
        RECT 720.630 1017.770 721.010 1017.780 ;
        RECT 717.870 1017.470 721.010 1017.770 ;
        RECT 717.870 1017.460 718.250 1017.470 ;
        RECT 720.630 1017.460 721.010 1017.470 ;
        RECT 717.870 955.890 718.250 955.900 ;
        RECT 720.630 955.890 721.010 955.900 ;
        RECT 717.870 955.590 721.010 955.890 ;
        RECT 717.870 955.580 718.250 955.590 ;
        RECT 720.630 955.580 721.010 955.590 ;
        RECT 717.870 921.210 718.250 921.220 ;
        RECT 720.630 921.210 721.010 921.220 ;
        RECT 717.870 920.910 721.010 921.210 ;
        RECT 717.870 920.900 718.250 920.910 ;
        RECT 720.630 920.900 721.010 920.910 ;
        RECT 720.630 525.450 721.010 525.460 ;
        RECT 717.910 525.150 721.010 525.450 ;
        RECT 717.910 524.780 718.210 525.150 ;
        RECT 720.630 525.140 721.010 525.150 ;
        RECT 717.870 524.460 718.250 524.780 ;
        RECT 717.665 517.300 717.995 517.305 ;
        RECT 717.665 517.290 718.250 517.300 ;
        RECT 717.440 516.990 718.250 517.290 ;
        RECT 717.665 516.980 718.250 516.990 ;
        RECT 717.665 516.975 717.995 516.980 ;
        RECT 717.665 475.820 717.995 475.825 ;
        RECT 717.665 475.810 718.250 475.820 ;
        RECT 717.665 475.510 718.450 475.810 ;
        RECT 717.665 475.500 718.250 475.510 ;
        RECT 717.665 475.495 717.995 475.500 ;
        RECT 717.870 438.410 718.250 438.420 ;
        RECT 720.630 438.410 721.010 438.420 ;
        RECT 717.870 438.110 721.010 438.410 ;
        RECT 717.870 438.100 718.250 438.110 ;
        RECT 720.630 438.100 721.010 438.110 ;
        RECT 720.630 58.290 721.010 58.300 ;
        RECT 2678.645 58.290 2678.975 58.305 ;
        RECT 720.630 57.990 2678.975 58.290 ;
        RECT 720.630 57.980 721.010 57.990 ;
        RECT 2678.645 57.975 2678.975 57.990 ;
      LAYER via3 ;
        RECT 717.900 2245.540 718.220 2245.860 ;
        RECT 717.900 2211.540 718.220 2211.860 ;
        RECT 718.820 2085.740 719.140 2086.060 ;
        RECT 718.820 2052.420 719.140 2052.740 ;
        RECT 716.060 2005.500 716.380 2005.820 ;
        RECT 716.060 1963.340 716.380 1963.660 ;
        RECT 717.900 1938.180 718.220 1938.500 ;
        RECT 717.900 1917.780 718.220 1918.100 ;
        RECT 717.670 1917.100 717.990 1917.420 ;
        RECT 716.060 1816.460 716.380 1816.780 ;
        RECT 718.820 1815.100 719.140 1815.420 ;
        RECT 716.060 1811.020 716.380 1811.340 ;
        RECT 718.820 1811.020 719.140 1811.340 ;
        RECT 716.060 1625.380 716.380 1625.700 ;
        RECT 718.820 1625.380 719.140 1625.700 ;
        RECT 718.820 1579.140 719.140 1579.460 ;
        RECT 718.820 1571.660 719.140 1571.980 ;
        RECT 718.820 1562.140 719.140 1562.460 ;
        RECT 718.820 1504.340 719.140 1504.660 ;
        RECT 718.820 1498.900 719.140 1499.220 ;
        RECT 715.140 1430.900 715.460 1431.220 ;
        RECT 715.140 1403.020 715.460 1403.340 ;
        RECT 716.980 1401.660 717.300 1401.980 ;
        RECT 716.980 1355.420 717.300 1355.740 ;
        RECT 718.820 1347.260 719.140 1347.580 ;
        RECT 717.900 1321.420 718.220 1321.740 ;
        RECT 720.660 1321.420 720.980 1321.740 ;
        RECT 717.900 1210.580 718.220 1210.900 ;
        RECT 720.660 1210.580 720.980 1210.900 ;
        RECT 717.900 1052.140 718.220 1052.460 ;
        RECT 720.660 1052.140 720.980 1052.460 ;
        RECT 717.900 1017.460 718.220 1017.780 ;
        RECT 720.660 1017.460 720.980 1017.780 ;
        RECT 717.900 955.580 718.220 955.900 ;
        RECT 720.660 955.580 720.980 955.900 ;
        RECT 717.900 920.900 718.220 921.220 ;
        RECT 720.660 920.900 720.980 921.220 ;
        RECT 720.660 525.140 720.980 525.460 ;
        RECT 717.900 524.460 718.220 524.780 ;
        RECT 717.900 516.980 718.220 517.300 ;
        RECT 717.900 475.500 718.220 475.820 ;
        RECT 717.900 438.100 718.220 438.420 ;
        RECT 720.660 438.100 720.980 438.420 ;
        RECT 720.660 57.980 720.980 58.300 ;
      LAYER met4 ;
        RECT 717.895 2245.535 718.225 2245.865 ;
        RECT 717.910 2211.865 718.210 2245.535 ;
        RECT 717.895 2211.535 718.225 2211.865 ;
        RECT 718.815 2086.050 719.145 2086.065 ;
        RECT 718.815 2085.750 720.050 2086.050 ;
        RECT 718.815 2085.735 719.145 2085.750 ;
        RECT 719.750 2072.450 720.050 2085.750 ;
        RECT 718.830 2072.150 720.050 2072.450 ;
        RECT 718.830 2052.745 719.130 2072.150 ;
        RECT 718.815 2052.415 719.145 2052.745 ;
        RECT 716.055 2005.495 716.385 2005.825 ;
        RECT 716.070 1963.665 716.370 2005.495 ;
        RECT 716.055 1963.335 716.385 1963.665 ;
        RECT 717.895 1938.175 718.225 1938.505 ;
        RECT 717.910 1918.105 718.210 1938.175 ;
        RECT 717.895 1917.775 718.225 1918.105 ;
        RECT 717.665 1917.095 717.995 1917.425 ;
        RECT 717.680 1916.050 717.980 1917.095 ;
        RECT 717.680 1915.750 718.210 1916.050 ;
        RECT 717.910 1909.250 718.210 1915.750 ;
        RECT 716.070 1908.950 718.210 1909.250 ;
        RECT 716.070 1816.785 716.370 1908.950 ;
        RECT 716.055 1816.455 716.385 1816.785 ;
        RECT 718.815 1815.095 719.145 1815.425 ;
        RECT 718.830 1811.345 719.130 1815.095 ;
        RECT 716.055 1811.015 716.385 1811.345 ;
        RECT 718.815 1811.015 719.145 1811.345 ;
        RECT 716.070 1625.705 716.370 1811.015 ;
        RECT 716.055 1625.375 716.385 1625.705 ;
        RECT 718.815 1625.690 719.145 1625.705 ;
        RECT 718.815 1625.390 720.970 1625.690 ;
        RECT 718.815 1625.375 719.145 1625.390 ;
        RECT 718.815 1579.450 719.145 1579.465 ;
        RECT 720.670 1579.450 720.970 1625.390 ;
        RECT 718.815 1579.150 720.970 1579.450 ;
        RECT 718.815 1579.135 719.145 1579.150 ;
        RECT 718.815 1571.655 719.145 1571.985 ;
        RECT 718.830 1569.250 719.130 1571.655 ;
        RECT 718.830 1568.950 722.810 1569.250 ;
        RECT 718.815 1562.450 719.145 1562.465 ;
        RECT 722.510 1562.450 722.810 1568.950 ;
        RECT 718.815 1562.150 722.810 1562.450 ;
        RECT 718.815 1562.135 719.145 1562.150 ;
        RECT 718.815 1504.650 719.145 1504.665 ;
        RECT 718.815 1504.350 720.050 1504.650 ;
        RECT 718.815 1504.335 719.145 1504.350 ;
        RECT 719.750 1501.250 720.050 1504.350 ;
        RECT 718.830 1500.950 720.050 1501.250 ;
        RECT 718.830 1499.225 719.130 1500.950 ;
        RECT 718.815 1498.895 719.145 1499.225 ;
        RECT 715.135 1430.895 715.465 1431.225 ;
        RECT 715.150 1403.345 715.450 1430.895 ;
        RECT 715.135 1403.015 715.465 1403.345 ;
        RECT 716.975 1401.655 717.305 1401.985 ;
        RECT 716.990 1355.745 717.290 1401.655 ;
        RECT 716.975 1355.415 717.305 1355.745 ;
        RECT 718.815 1347.255 719.145 1347.585 ;
        RECT 718.830 1344.850 719.130 1347.255 ;
        RECT 718.830 1344.550 720.970 1344.850 ;
        RECT 720.670 1321.745 720.970 1344.550 ;
        RECT 717.895 1321.415 718.225 1321.745 ;
        RECT 720.655 1321.415 720.985 1321.745 ;
        RECT 717.910 1210.905 718.210 1321.415 ;
        RECT 717.895 1210.575 718.225 1210.905 ;
        RECT 720.655 1210.575 720.985 1210.905 ;
        RECT 720.670 1052.465 720.970 1210.575 ;
        RECT 717.895 1052.135 718.225 1052.465 ;
        RECT 720.655 1052.135 720.985 1052.465 ;
        RECT 717.910 1017.785 718.210 1052.135 ;
        RECT 717.895 1017.455 718.225 1017.785 ;
        RECT 720.655 1017.455 720.985 1017.785 ;
        RECT 720.670 955.905 720.970 1017.455 ;
        RECT 717.895 955.575 718.225 955.905 ;
        RECT 720.655 955.575 720.985 955.905 ;
        RECT 717.910 921.225 718.210 955.575 ;
        RECT 717.895 920.895 718.225 921.225 ;
        RECT 720.655 920.895 720.985 921.225 ;
        RECT 720.670 525.465 720.970 920.895 ;
        RECT 720.655 525.135 720.985 525.465 ;
        RECT 717.895 524.455 718.225 524.785 ;
        RECT 717.910 517.305 718.210 524.455 ;
        RECT 717.895 516.975 718.225 517.305 ;
        RECT 717.895 475.495 718.225 475.825 ;
        RECT 717.910 438.425 718.210 475.495 ;
        RECT 717.895 438.095 718.225 438.425 ;
        RECT 720.655 438.095 720.985 438.425 ;
        RECT 720.670 58.305 720.970 438.095 ;
        RECT 720.655 57.975 720.985 58.305 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 712.610 1328.280 712.930 1328.340 ;
        RECT 2691.070 1328.280 2691.390 1328.340 ;
        RECT 712.610 1328.140 2691.390 1328.280 ;
        RECT 712.610 1328.080 712.930 1328.140 ;
        RECT 2691.070 1328.080 2691.390 1328.140 ;
        RECT 2691.070 2.960 2691.390 3.020 ;
        RECT 2696.590 2.960 2696.910 3.020 ;
        RECT 2691.070 2.820 2696.910 2.960 ;
        RECT 2691.070 2.760 2691.390 2.820 ;
        RECT 2696.590 2.760 2696.910 2.820 ;
      LAYER via ;
        RECT 712.640 1328.080 712.900 1328.340 ;
        RECT 2691.100 1328.080 2691.360 1328.340 ;
        RECT 2691.100 2.760 2691.360 3.020 ;
        RECT 2696.620 2.760 2696.880 3.020 ;
      LAYER met2 ;
        RECT 712.630 1395.515 712.910 1395.885 ;
        RECT 712.700 1328.370 712.840 1395.515 ;
        RECT 712.640 1328.050 712.900 1328.370 ;
        RECT 2691.100 1328.050 2691.360 1328.370 ;
        RECT 2691.160 3.050 2691.300 1328.050 ;
        RECT 2691.100 2.730 2691.360 3.050 ;
        RECT 2696.620 2.730 2696.880 3.050 ;
        RECT 2696.680 2.400 2696.820 2.730 ;
        RECT 2696.470 -4.800 2697.030 2.400 ;
      LAYER via2 ;
        RECT 712.630 1395.560 712.910 1395.840 ;
      LAYER met3 ;
        RECT 712.605 1395.850 712.935 1395.865 ;
        RECT 715.810 1395.850 719.810 1395.855 ;
        RECT 712.605 1395.550 719.810 1395.850 ;
        RECT 712.605 1395.535 712.935 1395.550 ;
        RECT 715.810 1395.255 719.810 1395.550 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2711.770 2.960 2712.090 3.020 ;
        RECT 2714.530 2.960 2714.850 3.020 ;
        RECT 2711.770 2.820 2714.850 2.960 ;
        RECT 2711.770 2.760 2712.090 2.820 ;
        RECT 2714.530 2.760 2714.850 2.820 ;
      LAYER via ;
        RECT 2711.800 2.760 2712.060 3.020 ;
        RECT 2714.560 2.760 2714.820 3.020 ;
      LAYER met2 ;
        RECT 1062.690 2383.555 1062.970 2383.925 ;
        RECT 1062.760 2377.880 1062.900 2383.555 ;
        RECT 1062.740 2373.880 1063.020 2377.880 ;
        RECT 1758.210 2293.795 1758.490 2294.165 ;
        RECT 1758.280 2270.365 1758.420 2293.795 ;
        RECT 1758.210 2269.995 1758.490 2270.365 ;
        RECT 2711.790 2204.035 2712.070 2204.405 ;
        RECT 2711.860 3.050 2712.000 2204.035 ;
        RECT 2711.800 2.730 2712.060 3.050 ;
        RECT 2714.560 2.730 2714.820 3.050 ;
        RECT 2714.620 2.400 2714.760 2.730 ;
        RECT 2714.410 -4.800 2714.970 2.400 ;
      LAYER via2 ;
        RECT 1062.690 2383.600 1062.970 2383.880 ;
        RECT 1758.210 2293.840 1758.490 2294.120 ;
        RECT 1758.210 2270.040 1758.490 2270.320 ;
        RECT 2711.790 2204.080 2712.070 2204.360 ;
      LAYER met3 ;
        RECT 1739.070 2385.250 1739.450 2385.260 ;
        RECT 1754.710 2385.250 1755.090 2385.260 ;
        RECT 1739.070 2384.950 1755.090 2385.250 ;
        RECT 1739.070 2384.940 1739.450 2384.950 ;
        RECT 1754.710 2384.940 1755.090 2384.950 ;
        RECT 1062.665 2383.890 1062.995 2383.905 ;
        RECT 1084.030 2383.890 1084.410 2383.900 ;
        RECT 1062.665 2383.590 1084.410 2383.890 ;
        RECT 1062.665 2383.575 1062.995 2383.590 ;
        RECT 1084.030 2383.580 1084.410 2383.590 ;
        RECT 1758.185 2294.140 1758.515 2294.145 ;
        RECT 1758.185 2294.130 1758.770 2294.140 ;
        RECT 1758.185 2293.830 1758.970 2294.130 ;
        RECT 1758.185 2293.820 1758.770 2293.830 ;
        RECT 1758.185 2293.815 1758.515 2293.820 ;
        RECT 1757.470 2270.330 1757.850 2270.340 ;
        RECT 1758.185 2270.330 1758.515 2270.345 ;
        RECT 1757.470 2270.030 1758.515 2270.330 ;
        RECT 1757.470 2270.020 1757.850 2270.030 ;
        RECT 1758.185 2270.015 1758.515 2270.030 ;
        RECT 1758.390 2206.780 1758.770 2207.100 ;
        RECT 1758.430 2204.370 1758.730 2206.780 ;
        RECT 2711.765 2204.370 2712.095 2204.385 ;
        RECT 1758.430 2204.070 2712.095 2204.370 ;
        RECT 2711.765 2204.055 2712.095 2204.070 ;
      LAYER via3 ;
        RECT 1739.100 2384.940 1739.420 2385.260 ;
        RECT 1754.740 2384.940 1755.060 2385.260 ;
        RECT 1084.060 2383.580 1084.380 2383.900 ;
        RECT 1758.420 2293.820 1758.740 2294.140 ;
        RECT 1757.500 2270.020 1757.820 2270.340 ;
        RECT 1758.420 2206.780 1758.740 2207.100 ;
      LAYER met4 ;
        RECT 1083.630 2387.910 1084.810 2389.090 ;
        RECT 1738.670 2387.910 1739.850 2389.090 ;
        RECT 1084.070 2383.905 1084.370 2387.910 ;
        RECT 1739.110 2385.265 1739.410 2387.910 ;
        RECT 1739.095 2384.935 1739.425 2385.265 ;
        RECT 1754.735 2384.935 1755.065 2385.265 ;
        RECT 1084.055 2383.575 1084.385 2383.905 ;
        RECT 1754.750 2304.330 1755.050 2384.935 ;
        RECT 1754.750 2304.030 1758.730 2304.330 ;
        RECT 1758.430 2294.145 1758.730 2304.030 ;
        RECT 1758.415 2293.815 1758.745 2294.145 ;
        RECT 1757.495 2270.015 1757.825 2270.345 ;
        RECT 1757.510 2259.450 1757.810 2270.015 ;
        RECT 1757.510 2259.150 1758.730 2259.450 ;
        RECT 1758.430 2207.105 1758.730 2259.150 ;
        RECT 1758.415 2206.775 1758.745 2207.105 ;
      LAYER met5 ;
        RECT 1083.420 2387.700 1740.060 2389.300 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2542.490 20.300 2542.810 20.360 ;
        RECT 2732.470 20.300 2732.790 20.360 ;
        RECT 2542.490 20.160 2732.790 20.300 ;
        RECT 2542.490 20.100 2542.810 20.160 ;
        RECT 2732.470 20.100 2732.790 20.160 ;
      LAYER via ;
        RECT 2542.520 20.100 2542.780 20.360 ;
        RECT 2732.500 20.100 2732.760 20.360 ;
      LAYER met2 ;
        RECT 1282.570 2388.995 1282.850 2389.365 ;
        RECT 2542.510 2388.995 2542.790 2389.365 ;
        RECT 1282.640 2377.880 1282.780 2388.995 ;
        RECT 1282.620 2373.880 1282.900 2377.880 ;
        RECT 2542.580 20.390 2542.720 2388.995 ;
        RECT 2542.520 20.070 2542.780 20.390 ;
        RECT 2732.500 20.070 2732.760 20.390 ;
        RECT 2732.560 2.400 2732.700 20.070 ;
        RECT 2732.350 -4.800 2732.910 2.400 ;
      LAYER via2 ;
        RECT 1282.570 2389.040 1282.850 2389.320 ;
        RECT 2542.510 2389.040 2542.790 2389.320 ;
      LAYER met3 ;
        RECT 1282.545 2389.330 1282.875 2389.345 ;
        RECT 2542.485 2389.330 2542.815 2389.345 ;
        RECT 1282.545 2389.030 2542.815 2389.330 ;
        RECT 1282.545 2389.015 1282.875 2389.030 ;
        RECT 2542.485 2389.015 2542.815 2389.030 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1772.910 1573.420 1773.230 1573.480 ;
        RECT 2549.390 1573.420 2549.710 1573.480 ;
        RECT 1772.910 1573.280 2549.710 1573.420 ;
        RECT 1772.910 1573.220 1773.230 1573.280 ;
        RECT 2549.390 1573.220 2549.710 1573.280 ;
        RECT 2549.390 19.960 2549.710 20.020 ;
        RECT 2750.410 19.960 2750.730 20.020 ;
        RECT 2549.390 19.820 2750.730 19.960 ;
        RECT 2549.390 19.760 2549.710 19.820 ;
        RECT 2750.410 19.760 2750.730 19.820 ;
      LAYER via ;
        RECT 1772.940 1573.220 1773.200 1573.480 ;
        RECT 2549.420 1573.220 2549.680 1573.480 ;
        RECT 2549.420 19.760 2549.680 20.020 ;
        RECT 2750.440 19.760 2750.700 20.020 ;
      LAYER met2 ;
        RECT 1772.930 1579.115 1773.210 1579.485 ;
        RECT 1773.000 1573.510 1773.140 1579.115 ;
        RECT 1772.940 1573.190 1773.200 1573.510 ;
        RECT 2549.420 1573.190 2549.680 1573.510 ;
        RECT 2549.480 20.050 2549.620 1573.190 ;
        RECT 2549.420 19.730 2549.680 20.050 ;
        RECT 2750.440 19.730 2750.700 20.050 ;
        RECT 2750.500 2.400 2750.640 19.730 ;
        RECT 2750.290 -4.800 2750.850 2.400 ;
      LAYER via2 ;
        RECT 1772.930 1579.160 1773.210 1579.440 ;
      LAYER met3 ;
        RECT 1755.835 1579.450 1759.835 1579.455 ;
        RECT 1772.905 1579.450 1773.235 1579.465 ;
        RECT 1755.835 1579.150 1773.235 1579.450 ;
        RECT 1755.835 1578.855 1759.835 1579.150 ;
        RECT 1772.905 1579.135 1773.235 1579.150 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2766.990 79.035 2767.270 79.405 ;
        RECT 2767.060 17.410 2767.200 79.035 ;
        RECT 2767.060 17.270 2768.120 17.410 ;
        RECT 2767.980 2.400 2768.120 17.270 ;
        RECT 2767.770 -4.800 2768.330 2.400 ;
      LAYER via2 ;
        RECT 2766.990 79.080 2767.270 79.360 ;
      LAYER met3 ;
        RECT 698.550 1686.890 698.930 1686.900 ;
        RECT 715.810 1686.890 719.810 1686.895 ;
        RECT 698.550 1686.590 719.810 1686.890 ;
        RECT 698.550 1686.580 698.930 1686.590 ;
        RECT 715.810 1686.295 719.810 1686.590 ;
        RECT 698.550 79.370 698.930 79.380 ;
        RECT 2766.965 79.370 2767.295 79.385 ;
        RECT 698.550 79.070 2767.295 79.370 ;
        RECT 698.550 79.060 698.930 79.070 ;
        RECT 2766.965 79.055 2767.295 79.070 ;
      LAYER via3 ;
        RECT 698.580 1686.580 698.900 1686.900 ;
        RECT 698.580 79.060 698.900 79.380 ;
      LAYER met4 ;
        RECT 698.575 1686.575 698.905 1686.905 ;
        RECT 698.590 79.385 698.890 1686.575 ;
        RECT 698.575 79.055 698.905 79.385 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 728.325 1327.105 728.495 1333.055 ;
      LAYER mcon ;
        RECT 728.325 1332.885 728.495 1333.055 ;
      LAYER met1 ;
        RECT 690.990 2392.820 691.310 2392.880 ;
        RECT 1004.710 2392.820 1005.030 2392.880 ;
        RECT 690.990 2392.680 1005.030 2392.820 ;
        RECT 690.990 2392.620 691.310 2392.680 ;
        RECT 1004.710 2392.620 1005.030 2392.680 ;
        RECT 690.990 1333.040 691.310 1333.100 ;
        RECT 728.265 1333.040 728.555 1333.085 ;
        RECT 690.990 1332.900 728.555 1333.040 ;
        RECT 690.990 1332.840 691.310 1332.900 ;
        RECT 728.265 1332.855 728.555 1332.900 ;
        RECT 728.265 1327.260 728.555 1327.305 ;
        RECT 728.265 1327.120 759.300 1327.260 ;
        RECT 728.265 1327.075 728.555 1327.120 ;
        RECT 759.160 1326.580 759.300 1327.120 ;
        RECT 835.430 1326.580 835.750 1326.640 ;
        RECT 759.160 1326.440 835.750 1326.580 ;
        RECT 835.430 1326.380 835.750 1326.440 ;
        RECT 835.430 15.540 835.750 15.600 ;
        RECT 840.950 15.540 841.270 15.600 ;
        RECT 835.430 15.400 841.270 15.540 ;
        RECT 835.430 15.340 835.750 15.400 ;
        RECT 840.950 15.340 841.270 15.400 ;
      LAYER via ;
        RECT 691.020 2392.620 691.280 2392.880 ;
        RECT 1004.740 2392.620 1005.000 2392.880 ;
        RECT 691.020 1332.840 691.280 1333.100 ;
        RECT 835.460 1326.380 835.720 1326.640 ;
        RECT 835.460 15.340 835.720 15.600 ;
        RECT 840.980 15.340 841.240 15.600 ;
      LAYER met2 ;
        RECT 691.020 2392.590 691.280 2392.910 ;
        RECT 1004.740 2392.590 1005.000 2392.910 ;
        RECT 691.080 1393.845 691.220 2392.590 ;
        RECT 1004.800 2377.880 1004.940 2392.590 ;
        RECT 1004.780 2373.880 1005.060 2377.880 ;
        RECT 691.010 1393.475 691.290 1393.845 ;
        RECT 691.010 1392.115 691.290 1392.485 ;
        RECT 691.080 1333.130 691.220 1392.115 ;
        RECT 691.020 1332.810 691.280 1333.130 ;
        RECT 835.460 1326.350 835.720 1326.670 ;
        RECT 835.520 15.630 835.660 1326.350 ;
        RECT 835.460 15.310 835.720 15.630 ;
        RECT 840.980 15.310 841.240 15.630 ;
        RECT 841.040 2.400 841.180 15.310 ;
        RECT 840.830 -4.800 841.390 2.400 ;
      LAYER via2 ;
        RECT 691.010 1393.520 691.290 1393.800 ;
        RECT 691.010 1392.160 691.290 1392.440 ;
      LAYER met3 ;
        RECT 690.985 1393.810 691.315 1393.825 ;
        RECT 690.985 1393.495 691.530 1393.810 ;
        RECT 691.230 1392.465 691.530 1393.495 ;
        RECT 690.985 1392.150 691.530 1392.465 ;
        RECT 690.985 1392.135 691.315 1392.150 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2597.765 17.425 2597.935 19.635 ;
      LAYER mcon ;
        RECT 2597.765 19.465 2597.935 19.635 ;
      LAYER met1 ;
        RECT 2597.705 19.620 2597.995 19.665 ;
        RECT 2785.830 19.620 2786.150 19.680 ;
        RECT 2597.705 19.480 2786.150 19.620 ;
        RECT 2597.705 19.435 2597.995 19.480 ;
        RECT 2785.830 19.420 2786.150 19.480 ;
        RECT 2570.090 17.580 2570.410 17.640 ;
        RECT 2597.705 17.580 2597.995 17.625 ;
        RECT 2570.090 17.440 2597.995 17.580 ;
        RECT 2570.090 17.380 2570.410 17.440 ;
        RECT 2597.705 17.395 2597.995 17.440 ;
      LAYER via ;
        RECT 2785.860 19.420 2786.120 19.680 ;
        RECT 2570.120 17.380 2570.380 17.640 ;
      LAYER met2 ;
        RECT 1415.970 2390.355 1416.250 2390.725 ;
        RECT 2570.110 2390.355 2570.390 2390.725 ;
        RECT 1416.040 2377.880 1416.180 2390.355 ;
        RECT 1416.020 2373.880 1416.300 2377.880 ;
        RECT 2570.180 17.670 2570.320 2390.355 ;
        RECT 2785.860 19.390 2786.120 19.710 ;
        RECT 2570.120 17.350 2570.380 17.670 ;
        RECT 2785.920 2.400 2786.060 19.390 ;
        RECT 2785.710 -4.800 2786.270 2.400 ;
      LAYER via2 ;
        RECT 1415.970 2390.400 1416.250 2390.680 ;
        RECT 2570.110 2390.400 2570.390 2390.680 ;
      LAYER met3 ;
        RECT 1415.945 2390.690 1416.275 2390.705 ;
        RECT 2570.085 2390.690 2570.415 2390.705 ;
        RECT 1415.945 2390.390 2570.415 2390.690 ;
        RECT 1415.945 2390.375 1416.275 2390.390 ;
        RECT 2570.085 2390.375 2570.415 2390.390 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 711.690 58.720 712.010 58.780 ;
        RECT 2801.470 58.720 2801.790 58.780 ;
        RECT 711.690 58.580 2801.790 58.720 ;
        RECT 711.690 58.520 712.010 58.580 ;
        RECT 2801.470 58.520 2801.790 58.580 ;
      LAYER via ;
        RECT 711.720 58.520 711.980 58.780 ;
        RECT 2801.500 58.520 2801.760 58.780 ;
      LAYER met2 ;
        RECT 711.710 1463.515 711.990 1463.885 ;
        RECT 711.780 58.810 711.920 1463.515 ;
        RECT 711.720 58.490 711.980 58.810 ;
        RECT 2801.500 58.490 2801.760 58.810 ;
        RECT 2801.560 17.410 2801.700 58.490 ;
        RECT 2801.560 17.270 2804.000 17.410 ;
        RECT 2803.860 2.400 2804.000 17.270 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
      LAYER via2 ;
        RECT 711.710 1463.560 711.990 1463.840 ;
      LAYER met3 ;
        RECT 711.685 1463.850 712.015 1463.865 ;
        RECT 715.810 1463.850 719.810 1463.855 ;
        RECT 711.685 1463.550 719.810 1463.850 ;
        RECT 711.685 1463.535 712.015 1463.550 ;
        RECT 715.810 1463.255 719.810 1463.550 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2608.345 17.765 2608.515 19.295 ;
      LAYER mcon ;
        RECT 2608.345 19.125 2608.515 19.295 ;
      LAYER met1 ;
        RECT 1772.450 1352.760 1772.770 1352.820 ;
        RECT 2590.790 1352.760 2591.110 1352.820 ;
        RECT 1772.450 1352.620 2591.110 1352.760 ;
        RECT 1772.450 1352.560 1772.770 1352.620 ;
        RECT 2590.790 1352.560 2591.110 1352.620 ;
        RECT 2608.285 19.280 2608.575 19.325 ;
        RECT 2821.710 19.280 2822.030 19.340 ;
        RECT 2608.285 19.140 2822.030 19.280 ;
        RECT 2608.285 19.095 2608.575 19.140 ;
        RECT 2821.710 19.080 2822.030 19.140 ;
        RECT 2590.790 17.920 2591.110 17.980 ;
        RECT 2608.285 17.920 2608.575 17.965 ;
        RECT 2590.790 17.780 2608.575 17.920 ;
        RECT 2590.790 17.720 2591.110 17.780 ;
        RECT 2608.285 17.735 2608.575 17.780 ;
      LAYER via ;
        RECT 1772.480 1352.560 1772.740 1352.820 ;
        RECT 2590.820 1352.560 2591.080 1352.820 ;
        RECT 2821.740 19.080 2822.000 19.340 ;
        RECT 2590.820 17.720 2591.080 17.980 ;
      LAYER met2 ;
        RECT 1772.470 1356.075 1772.750 1356.445 ;
        RECT 1772.540 1352.850 1772.680 1356.075 ;
        RECT 1772.480 1352.530 1772.740 1352.850 ;
        RECT 2590.820 1352.530 2591.080 1352.850 ;
        RECT 2590.880 18.010 2591.020 1352.530 ;
        RECT 2821.740 19.050 2822.000 19.370 ;
        RECT 2590.820 17.690 2591.080 18.010 ;
        RECT 2821.800 2.400 2821.940 19.050 ;
        RECT 2821.590 -4.800 2822.150 2.400 ;
      LAYER via2 ;
        RECT 1772.470 1356.120 1772.750 1356.400 ;
      LAYER met3 ;
        RECT 1755.835 1356.410 1759.835 1356.415 ;
        RECT 1772.445 1356.410 1772.775 1356.425 ;
        RECT 1755.835 1356.110 1772.775 1356.410 ;
        RECT 1755.835 1355.815 1759.835 1356.110 ;
        RECT 1772.445 1356.095 1772.775 1356.110 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1270.590 2391.800 1270.910 2391.860 ;
        RECT 1711.270 2391.800 1711.590 2391.860 ;
        RECT 1270.590 2391.660 1711.590 2391.800 ;
        RECT 1270.590 2391.600 1270.910 2391.660 ;
        RECT 1711.270 2391.600 1711.590 2391.660 ;
        RECT 2604.590 19.280 2604.910 19.340 ;
        RECT 2604.590 19.140 2608.040 19.280 ;
        RECT 2604.590 19.080 2604.910 19.140 ;
        RECT 2607.900 18.940 2608.040 19.140 ;
        RECT 2839.190 18.940 2839.510 19.000 ;
        RECT 2607.900 18.800 2839.510 18.940 ;
        RECT 2839.190 18.740 2839.510 18.800 ;
      LAYER via ;
        RECT 1270.620 2391.600 1270.880 2391.860 ;
        RECT 1711.300 2391.600 1711.560 2391.860 ;
        RECT 2604.620 19.080 2604.880 19.340 ;
        RECT 2839.220 18.740 2839.480 19.000 ;
      LAYER met2 ;
        RECT 1270.620 2391.570 1270.880 2391.890 ;
        RECT 1711.300 2391.570 1711.560 2391.890 ;
        RECT 1270.680 2377.880 1270.820 2391.570 ;
        RECT 1711.360 2390.045 1711.500 2391.570 ;
        RECT 1711.290 2389.675 1711.570 2390.045 ;
        RECT 2604.610 2389.675 2604.890 2390.045 ;
        RECT 1270.660 2373.880 1270.940 2377.880 ;
        RECT 2604.680 19.370 2604.820 2389.675 ;
        RECT 2604.620 19.050 2604.880 19.370 ;
        RECT 2839.220 18.710 2839.480 19.030 ;
        RECT 2839.280 2.400 2839.420 18.710 ;
        RECT 2839.070 -4.800 2839.630 2.400 ;
      LAYER via2 ;
        RECT 1711.290 2389.720 1711.570 2390.000 ;
        RECT 2604.610 2389.720 2604.890 2390.000 ;
      LAYER met3 ;
        RECT 1711.265 2390.010 1711.595 2390.025 ;
        RECT 2604.585 2390.010 2604.915 2390.025 ;
        RECT 1711.265 2389.710 2604.915 2390.010 ;
        RECT 1711.265 2389.695 1711.595 2389.710 ;
        RECT 2604.585 2389.695 2604.915 2389.710 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1702.990 31.520 1703.310 31.580 ;
        RECT 2857.130 31.520 2857.450 31.580 ;
        RECT 1702.990 31.380 2857.450 31.520 ;
        RECT 1702.990 31.320 1703.310 31.380 ;
        RECT 2857.130 31.320 2857.450 31.380 ;
      LAYER via ;
        RECT 1703.020 31.320 1703.280 31.580 ;
        RECT 2857.160 31.320 2857.420 31.580 ;
      LAYER met2 ;
        RECT 1701.220 1323.690 1701.500 1327.135 ;
        RECT 1701.220 1323.550 1703.680 1323.690 ;
        RECT 1701.220 1323.135 1701.500 1323.550 ;
        RECT 1703.540 46.650 1703.680 1323.550 ;
        RECT 1703.080 46.510 1703.680 46.650 ;
        RECT 1703.080 31.610 1703.220 46.510 ;
        RECT 1703.020 31.290 1703.280 31.610 ;
        RECT 2857.160 31.290 2857.420 31.610 ;
        RECT 2857.220 2.400 2857.360 31.290 ;
        RECT 2857.010 -4.800 2857.570 2.400 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2608.805 16.745 2608.975 17.935 ;
      LAYER mcon ;
        RECT 2608.805 17.765 2608.975 17.935 ;
      LAYER met1 ;
        RECT 1771.070 2360.180 1771.390 2360.240 ;
        RECT 2605.050 2360.180 2605.370 2360.240 ;
        RECT 1771.070 2360.040 2605.370 2360.180 ;
        RECT 1771.070 2359.980 1771.390 2360.040 ;
        RECT 2605.050 2359.980 2605.370 2360.040 ;
        RECT 2608.745 17.920 2609.035 17.965 ;
        RECT 2875.070 17.920 2875.390 17.980 ;
        RECT 2608.745 17.780 2875.390 17.920 ;
        RECT 2608.745 17.735 2609.035 17.780 ;
        RECT 2875.070 17.720 2875.390 17.780 ;
        RECT 2605.050 16.900 2605.370 16.960 ;
        RECT 2608.745 16.900 2609.035 16.945 ;
        RECT 2605.050 16.760 2609.035 16.900 ;
        RECT 2605.050 16.700 2605.370 16.760 ;
        RECT 2608.745 16.715 2609.035 16.760 ;
      LAYER via ;
        RECT 1771.100 2359.980 1771.360 2360.240 ;
        RECT 2605.080 2359.980 2605.340 2360.240 ;
        RECT 2875.100 17.720 2875.360 17.980 ;
        RECT 2605.080 16.700 2605.340 16.960 ;
      LAYER met2 ;
        RECT 1771.090 2365.195 1771.370 2365.565 ;
        RECT 1771.160 2360.270 1771.300 2365.195 ;
        RECT 1771.100 2359.950 1771.360 2360.270 ;
        RECT 2605.080 2359.950 2605.340 2360.270 ;
        RECT 2605.140 16.990 2605.280 2359.950 ;
        RECT 2875.100 17.690 2875.360 18.010 ;
        RECT 2605.080 16.670 2605.340 16.990 ;
        RECT 2875.160 2.400 2875.300 17.690 ;
        RECT 2874.950 -4.800 2875.510 2.400 ;
      LAYER via2 ;
        RECT 1771.090 2365.240 1771.370 2365.520 ;
      LAYER met3 ;
        RECT 1755.835 2365.530 1759.835 2365.535 ;
        RECT 1771.065 2365.530 1771.395 2365.545 ;
        RECT 1755.835 2365.230 1771.395 2365.530 ;
        RECT 1755.835 2364.935 1759.835 2365.230 ;
        RECT 1771.065 2365.215 1771.395 2365.230 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1772.910 1435.380 1773.230 1435.440 ;
        RECT 2625.290 1435.380 2625.610 1435.440 ;
        RECT 1772.910 1435.240 2625.610 1435.380 ;
        RECT 1772.910 1435.180 1773.230 1435.240 ;
        RECT 2625.290 1435.180 2625.610 1435.240 ;
        RECT 2624.830 17.580 2625.150 17.640 ;
        RECT 2893.010 17.580 2893.330 17.640 ;
        RECT 2624.830 17.440 2893.330 17.580 ;
        RECT 2624.830 17.380 2625.150 17.440 ;
        RECT 2893.010 17.380 2893.330 17.440 ;
      LAYER via ;
        RECT 1772.940 1435.180 1773.200 1435.440 ;
        RECT 2625.320 1435.180 2625.580 1435.440 ;
        RECT 2624.860 17.380 2625.120 17.640 ;
        RECT 2893.040 17.380 2893.300 17.640 ;
      LAYER met2 ;
        RECT 1772.930 1441.755 1773.210 1442.125 ;
        RECT 1773.000 1435.470 1773.140 1441.755 ;
        RECT 1772.940 1435.150 1773.200 1435.470 ;
        RECT 2625.320 1435.150 2625.580 1435.470 ;
        RECT 2625.380 39.850 2625.520 1435.150 ;
        RECT 2624.920 39.710 2625.520 39.850 ;
        RECT 2624.920 17.670 2625.060 39.710 ;
        RECT 2624.860 17.350 2625.120 17.670 ;
        RECT 2893.040 17.350 2893.300 17.670 ;
        RECT 2893.100 2.400 2893.240 17.350 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
      LAYER via2 ;
        RECT 1772.930 1441.800 1773.210 1442.080 ;
      LAYER met3 ;
        RECT 1755.835 1442.090 1759.835 1442.095 ;
        RECT 1772.905 1442.090 1773.235 1442.105 ;
        RECT 1755.835 1441.790 1773.235 1442.090 ;
        RECT 1755.835 1441.495 1759.835 1441.790 ;
        RECT 1772.905 1441.775 1773.235 1441.790 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 863.030 1311.620 863.350 1311.680 ;
        RECT 869.010 1311.620 869.330 1311.680 ;
        RECT 863.030 1311.480 869.330 1311.620 ;
        RECT 863.030 1311.420 863.350 1311.480 ;
        RECT 869.010 1311.420 869.330 1311.480 ;
        RECT 869.010 30.840 869.330 30.900 ;
        RECT 2910.950 30.840 2911.270 30.900 ;
        RECT 869.010 30.700 2911.270 30.840 ;
        RECT 869.010 30.640 869.330 30.700 ;
        RECT 2910.950 30.640 2911.270 30.700 ;
      LAYER via ;
        RECT 863.060 1311.420 863.320 1311.680 ;
        RECT 869.040 1311.420 869.300 1311.680 ;
        RECT 869.040 30.640 869.300 30.900 ;
        RECT 2910.980 30.640 2911.240 30.900 ;
      LAYER met2 ;
        RECT 863.100 1323.135 863.380 1327.135 ;
        RECT 863.120 1311.710 863.260 1323.135 ;
        RECT 863.060 1311.390 863.320 1311.710 ;
        RECT 869.040 1311.390 869.300 1311.710 ;
        RECT 869.100 30.930 869.240 1311.390 ;
        RECT 869.040 30.610 869.300 30.930 ;
        RECT 2910.980 30.610 2911.240 30.930 ;
        RECT 2911.040 2.400 2911.180 30.610 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 724.570 655.420 724.890 655.480 ;
        RECT 725.490 655.420 725.810 655.480 ;
        RECT 724.570 655.280 725.810 655.420 ;
        RECT 724.570 655.220 724.890 655.280 ;
        RECT 725.490 655.220 725.810 655.280 ;
      LAYER via ;
        RECT 724.600 655.220 724.860 655.480 ;
        RECT 725.520 655.220 725.780 655.480 ;
      LAYER met2 ;
        RECT 724.590 1277.875 724.870 1278.245 ;
        RECT 724.660 1210.925 724.800 1277.875 ;
        RECT 724.590 1210.555 724.870 1210.925 ;
        RECT 725.050 1162.275 725.330 1162.645 ;
        RECT 725.120 1055.885 725.260 1162.275 ;
        RECT 725.050 1055.515 725.330 1055.885 ;
        RECT 725.050 965.075 725.330 965.445 ;
        RECT 725.120 921.245 725.260 965.075 ;
        RECT 725.050 920.875 725.330 921.245 ;
        RECT 725.970 885.515 726.250 885.885 ;
        RECT 726.040 824.685 726.180 885.515 ;
        RECT 725.970 824.315 726.250 824.685 ;
        RECT 724.590 679.475 724.870 679.845 ;
        RECT 724.660 655.510 724.800 679.475 ;
        RECT 724.600 655.190 724.860 655.510 ;
        RECT 725.520 655.190 725.780 655.510 ;
        RECT 725.580 572.405 725.720 655.190 ;
        RECT 725.510 572.035 725.790 572.405 ;
        RECT 725.510 548.235 725.790 548.605 ;
        RECT 725.580 524.805 725.720 548.235 ;
        RECT 725.510 524.435 725.790 524.805 ;
        RECT 727.350 396.595 727.630 396.965 ;
        RECT 727.420 341.885 727.560 396.595 ;
        RECT 727.350 341.515 727.630 341.885 ;
        RECT 724.590 306.835 724.870 307.205 ;
        RECT 724.660 269.125 724.800 306.835 ;
        RECT 724.590 268.755 724.870 269.125 ;
        RECT 725.510 268.755 725.790 269.125 ;
        RECT 725.580 187.525 725.720 268.755 ;
        RECT 725.510 187.155 725.790 187.525 ;
        RECT 725.510 51.835 725.790 52.205 ;
        RECT 725.580 14.805 725.720 51.835 ;
        RECT 725.510 14.435 725.790 14.805 ;
        RECT 858.910 14.435 859.190 14.805 ;
        RECT 858.980 2.400 859.120 14.435 ;
        RECT 858.770 -4.800 859.330 2.400 ;
      LAYER via2 ;
        RECT 724.590 1277.920 724.870 1278.200 ;
        RECT 724.590 1210.600 724.870 1210.880 ;
        RECT 725.050 1162.320 725.330 1162.600 ;
        RECT 725.050 1055.560 725.330 1055.840 ;
        RECT 725.050 965.120 725.330 965.400 ;
        RECT 725.050 920.920 725.330 921.200 ;
        RECT 725.970 885.560 726.250 885.840 ;
        RECT 725.970 824.360 726.250 824.640 ;
        RECT 724.590 679.520 724.870 679.800 ;
        RECT 725.510 572.080 725.790 572.360 ;
        RECT 725.510 548.280 725.790 548.560 ;
        RECT 725.510 524.480 725.790 524.760 ;
        RECT 727.350 396.640 727.630 396.920 ;
        RECT 727.350 341.560 727.630 341.840 ;
        RECT 724.590 306.880 724.870 307.160 ;
        RECT 724.590 268.800 724.870 269.080 ;
        RECT 725.510 268.800 725.790 269.080 ;
        RECT 725.510 187.200 725.790 187.480 ;
        RECT 725.510 51.880 725.790 52.160 ;
        RECT 725.510 14.480 725.790 14.760 ;
        RECT 858.910 14.480 859.190 14.760 ;
      LAYER met3 ;
        RECT 704.990 1720.890 705.370 1720.900 ;
        RECT 715.810 1720.890 719.810 1720.895 ;
        RECT 704.990 1720.590 719.810 1720.890 ;
        RECT 704.990 1720.580 705.370 1720.590 ;
        RECT 715.810 1720.295 719.810 1720.590 ;
        RECT 704.990 1306.770 705.370 1306.780 ;
        RECT 725.230 1306.770 725.610 1306.780 ;
        RECT 704.990 1306.470 725.610 1306.770 ;
        RECT 704.990 1306.460 705.370 1306.470 ;
        RECT 725.230 1306.460 725.610 1306.470 ;
        RECT 724.565 1278.210 724.895 1278.225 ;
        RECT 725.230 1278.210 725.610 1278.220 ;
        RECT 724.565 1277.910 725.610 1278.210 ;
        RECT 724.565 1277.895 724.895 1277.910 ;
        RECT 725.230 1277.900 725.610 1277.910 ;
        RECT 724.565 1210.900 724.895 1210.905 ;
        RECT 724.310 1210.890 724.895 1210.900 ;
        RECT 724.110 1210.590 724.895 1210.890 ;
        RECT 724.310 1210.580 724.895 1210.590 ;
        RECT 724.565 1210.575 724.895 1210.580 ;
        RECT 724.310 1162.610 724.690 1162.620 ;
        RECT 725.025 1162.610 725.355 1162.625 ;
        RECT 724.310 1162.310 725.355 1162.610 ;
        RECT 724.310 1162.300 724.690 1162.310 ;
        RECT 725.025 1162.295 725.355 1162.310 ;
        RECT 725.025 1055.860 725.355 1055.865 ;
        RECT 725.025 1055.850 725.610 1055.860 ;
        RECT 724.800 1055.550 725.610 1055.850 ;
        RECT 725.025 1055.540 725.610 1055.550 ;
        RECT 725.025 1055.535 725.355 1055.540 ;
        RECT 725.025 965.420 725.355 965.425 ;
        RECT 725.025 965.410 725.610 965.420 ;
        RECT 724.800 965.110 725.610 965.410 ;
        RECT 725.025 965.100 725.610 965.110 ;
        RECT 725.025 965.095 725.355 965.100 ;
        RECT 725.025 921.220 725.355 921.225 ;
        RECT 725.025 921.210 725.610 921.220 ;
        RECT 724.800 920.910 725.610 921.210 ;
        RECT 725.025 920.900 725.610 920.910 ;
        RECT 725.025 920.895 725.355 920.900 ;
        RECT 725.230 885.850 725.610 885.860 ;
        RECT 725.945 885.850 726.275 885.865 ;
        RECT 725.230 885.550 726.275 885.850 ;
        RECT 725.230 885.540 725.610 885.550 ;
        RECT 725.945 885.535 726.275 885.550 ;
        RECT 725.230 824.650 725.610 824.660 ;
        RECT 725.945 824.650 726.275 824.665 ;
        RECT 725.230 824.350 726.275 824.650 ;
        RECT 725.230 824.340 725.610 824.350 ;
        RECT 725.945 824.335 726.275 824.350 ;
        RECT 725.230 773.650 725.610 773.660 ;
        RECT 724.350 773.350 725.610 773.650 ;
        RECT 724.350 772.300 724.650 773.350 ;
        RECT 725.230 773.340 725.610 773.350 ;
        RECT 724.310 771.980 724.690 772.300 ;
        RECT 724.565 679.810 724.895 679.825 ;
        RECT 725.230 679.810 725.610 679.820 ;
        RECT 724.565 679.510 725.610 679.810 ;
        RECT 724.565 679.495 724.895 679.510 ;
        RECT 725.230 679.500 725.610 679.510 ;
        RECT 725.485 572.380 725.815 572.385 ;
        RECT 725.230 572.370 725.815 572.380 ;
        RECT 725.030 572.070 725.815 572.370 ;
        RECT 725.230 572.060 725.815 572.070 ;
        RECT 725.485 572.055 725.815 572.060 ;
        RECT 725.485 548.580 725.815 548.585 ;
        RECT 725.230 548.570 725.815 548.580 ;
        RECT 725.030 548.270 725.815 548.570 ;
        RECT 725.230 548.260 725.815 548.270 ;
        RECT 725.485 548.255 725.815 548.260 ;
        RECT 725.485 524.770 725.815 524.785 ;
        RECT 726.150 524.770 726.530 524.780 ;
        RECT 725.485 524.470 726.530 524.770 ;
        RECT 725.485 524.455 725.815 524.470 ;
        RECT 726.150 524.460 726.530 524.470 ;
        RECT 725.230 396.930 725.610 396.940 ;
        RECT 727.325 396.930 727.655 396.945 ;
        RECT 725.230 396.630 727.655 396.930 ;
        RECT 725.230 396.620 725.610 396.630 ;
        RECT 727.325 396.615 727.655 396.630 ;
        RECT 727.325 341.850 727.655 341.865 ;
        RECT 727.990 341.850 728.370 341.860 ;
        RECT 727.325 341.550 728.370 341.850 ;
        RECT 727.325 341.535 727.655 341.550 ;
        RECT 727.990 341.540 728.370 341.550 ;
        RECT 724.565 307.170 724.895 307.185 ;
        RECT 727.990 307.170 728.370 307.180 ;
        RECT 724.565 306.870 728.370 307.170 ;
        RECT 724.565 306.855 724.895 306.870 ;
        RECT 727.990 306.860 728.370 306.870 ;
        RECT 724.565 269.090 724.895 269.105 ;
        RECT 725.485 269.090 725.815 269.105 ;
        RECT 724.565 268.790 725.815 269.090 ;
        RECT 724.565 268.775 724.895 268.790 ;
        RECT 725.485 268.775 725.815 268.790 ;
        RECT 725.485 187.490 725.815 187.505 ;
        RECT 725.270 187.175 725.815 187.490 ;
        RECT 725.270 186.820 725.570 187.175 ;
        RECT 725.230 186.500 725.610 186.820 ;
        RECT 725.485 52.180 725.815 52.185 ;
        RECT 725.230 52.170 725.815 52.180 ;
        RECT 725.030 51.870 725.815 52.170 ;
        RECT 725.230 51.860 725.815 51.870 ;
        RECT 725.485 51.855 725.815 51.860 ;
        RECT 725.485 14.770 725.815 14.785 ;
        RECT 858.885 14.770 859.215 14.785 ;
        RECT 725.485 14.470 859.215 14.770 ;
        RECT 725.485 14.455 725.815 14.470 ;
        RECT 858.885 14.455 859.215 14.470 ;
      LAYER via3 ;
        RECT 705.020 1720.580 705.340 1720.900 ;
        RECT 705.020 1306.460 705.340 1306.780 ;
        RECT 725.260 1306.460 725.580 1306.780 ;
        RECT 725.260 1277.900 725.580 1278.220 ;
        RECT 724.340 1210.580 724.660 1210.900 ;
        RECT 724.340 1162.300 724.660 1162.620 ;
        RECT 725.260 1055.540 725.580 1055.860 ;
        RECT 725.260 965.100 725.580 965.420 ;
        RECT 725.260 920.900 725.580 921.220 ;
        RECT 725.260 885.540 725.580 885.860 ;
        RECT 725.260 824.340 725.580 824.660 ;
        RECT 725.260 773.340 725.580 773.660 ;
        RECT 724.340 771.980 724.660 772.300 ;
        RECT 725.260 679.500 725.580 679.820 ;
        RECT 725.260 572.060 725.580 572.380 ;
        RECT 725.260 548.260 725.580 548.580 ;
        RECT 726.180 524.460 726.500 524.780 ;
        RECT 725.260 396.620 725.580 396.940 ;
        RECT 728.020 341.540 728.340 341.860 ;
        RECT 728.020 306.860 728.340 307.180 ;
        RECT 725.260 186.500 725.580 186.820 ;
        RECT 725.260 51.860 725.580 52.180 ;
      LAYER met4 ;
        RECT 705.015 1720.575 705.345 1720.905 ;
        RECT 705.030 1306.785 705.330 1720.575 ;
        RECT 705.015 1306.455 705.345 1306.785 ;
        RECT 725.255 1306.455 725.585 1306.785 ;
        RECT 725.270 1278.225 725.570 1306.455 ;
        RECT 725.255 1277.895 725.585 1278.225 ;
        RECT 724.335 1210.575 724.665 1210.905 ;
        RECT 724.350 1162.625 724.650 1210.575 ;
        RECT 724.335 1162.295 724.665 1162.625 ;
        RECT 725.255 1055.535 725.585 1055.865 ;
        RECT 725.270 965.425 725.570 1055.535 ;
        RECT 725.255 965.095 725.585 965.425 ;
        RECT 725.255 920.895 725.585 921.225 ;
        RECT 725.270 885.865 725.570 920.895 ;
        RECT 725.255 885.535 725.585 885.865 ;
        RECT 725.255 824.335 725.585 824.665 ;
        RECT 725.270 773.665 725.570 824.335 ;
        RECT 725.255 773.335 725.585 773.665 ;
        RECT 724.335 771.975 724.665 772.305 ;
        RECT 724.350 729.450 724.650 771.975 ;
        RECT 724.350 729.150 725.570 729.450 ;
        RECT 725.270 679.825 725.570 729.150 ;
        RECT 725.255 679.495 725.585 679.825 ;
        RECT 725.255 572.055 725.585 572.385 ;
        RECT 725.270 548.585 725.570 572.055 ;
        RECT 725.255 548.255 725.585 548.585 ;
        RECT 726.175 524.455 726.505 524.785 ;
        RECT 726.190 484.650 726.490 524.455 ;
        RECT 725.270 484.350 726.490 484.650 ;
        RECT 725.270 396.945 725.570 484.350 ;
        RECT 725.255 396.615 725.585 396.945 ;
        RECT 728.015 341.535 728.345 341.865 ;
        RECT 728.030 307.185 728.330 341.535 ;
        RECT 728.015 306.855 728.345 307.185 ;
        RECT 725.255 186.495 725.585 186.825 ;
        RECT 725.270 137.850 725.570 186.495 ;
        RECT 724.350 137.550 725.570 137.850 ;
        RECT 724.350 114.050 724.650 137.550 ;
        RECT 724.350 113.750 725.570 114.050 ;
        RECT 725.270 52.185 725.570 113.750 ;
        RECT 725.255 51.855 725.585 52.185 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 720.505 1326.425 720.675 1352.775 ;
      LAYER mcon ;
        RECT 720.505 1352.605 720.675 1352.775 ;
      LAYER met1 ;
        RECT 717.210 1352.760 717.530 1352.820 ;
        RECT 720.445 1352.760 720.735 1352.805 ;
        RECT 717.210 1352.620 720.735 1352.760 ;
        RECT 717.210 1352.560 717.530 1352.620 ;
        RECT 720.445 1352.575 720.735 1352.620 ;
        RECT 720.445 1326.580 720.735 1326.625 ;
        RECT 721.350 1326.580 721.670 1326.640 ;
        RECT 720.445 1326.440 721.670 1326.580 ;
        RECT 720.445 1326.395 720.735 1326.440 ;
        RECT 721.350 1326.380 721.670 1326.440 ;
      LAYER via ;
        RECT 717.240 1352.560 717.500 1352.820 ;
        RECT 721.380 1326.380 721.640 1326.640 ;
      LAYER met2 ;
        RECT 1553.970 2392.395 1554.250 2392.765 ;
        RECT 1554.040 2377.880 1554.180 2392.395 ;
        RECT 1554.020 2373.880 1554.300 2377.880 ;
        RECT 715.390 2314.875 715.670 2315.245 ;
        RECT 715.460 2280.565 715.600 2314.875 ;
        RECT 715.390 2280.195 715.670 2280.565 ;
        RECT 713.550 1859.275 713.830 1859.645 ;
        RECT 713.620 1848.085 713.760 1859.275 ;
        RECT 713.550 1847.715 713.830 1848.085 ;
        RECT 717.230 1352.675 717.510 1353.045 ;
        RECT 717.240 1352.530 717.500 1352.675 ;
        RECT 721.380 1326.350 721.640 1326.670 ;
        RECT 721.440 1325.165 721.580 1326.350 ;
        RECT 721.370 1324.795 721.650 1325.165 ;
        RECT 876.850 14.435 877.130 14.805 ;
        RECT 876.920 2.400 877.060 14.435 ;
        RECT 876.710 -4.800 877.270 2.400 ;
      LAYER via2 ;
        RECT 1553.970 2392.440 1554.250 2392.720 ;
        RECT 715.390 2314.920 715.670 2315.200 ;
        RECT 715.390 2280.240 715.670 2280.520 ;
        RECT 713.550 1859.320 713.830 1859.600 ;
        RECT 713.550 1847.760 713.830 1848.040 ;
        RECT 717.230 1352.720 717.510 1353.000 ;
        RECT 721.370 1324.840 721.650 1325.120 ;
        RECT 876.850 14.480 877.130 14.760 ;
      LAYER met3 ;
        RECT 715.110 2392.730 715.490 2392.740 ;
        RECT 1553.945 2392.730 1554.275 2392.745 ;
        RECT 715.110 2392.430 1554.275 2392.730 ;
        RECT 715.110 2392.420 715.490 2392.430 ;
        RECT 1553.945 2392.415 1554.275 2392.430 ;
        RECT 715.365 2315.220 715.695 2315.225 ;
        RECT 715.110 2315.210 715.695 2315.220 ;
        RECT 714.910 2314.910 715.695 2315.210 ;
        RECT 715.110 2314.900 715.695 2314.910 ;
        RECT 715.365 2314.895 715.695 2314.900 ;
        RECT 715.365 2280.540 715.695 2280.545 ;
        RECT 715.110 2280.530 715.695 2280.540 ;
        RECT 714.910 2280.230 715.695 2280.530 ;
        RECT 715.110 2280.220 715.695 2280.230 ;
        RECT 715.365 2280.215 715.695 2280.220 ;
        RECT 713.525 1859.610 713.855 1859.625 ;
        RECT 715.110 1859.610 715.490 1859.620 ;
        RECT 713.525 1859.310 715.490 1859.610 ;
        RECT 713.525 1859.295 713.855 1859.310 ;
        RECT 715.110 1859.300 715.490 1859.310 ;
        RECT 713.525 1848.050 713.855 1848.065 ;
        RECT 715.110 1848.050 715.490 1848.060 ;
        RECT 713.525 1847.750 715.490 1848.050 ;
        RECT 713.525 1847.735 713.855 1847.750 ;
        RECT 715.110 1847.740 715.490 1847.750 ;
        RECT 715.110 1491.050 715.490 1491.060 ;
        RECT 718.790 1491.050 719.170 1491.060 ;
        RECT 715.110 1490.750 719.170 1491.050 ;
        RECT 715.110 1490.740 715.490 1490.750 ;
        RECT 718.790 1490.740 719.170 1490.750 ;
        RECT 717.870 1358.450 718.250 1358.460 ;
        RECT 717.870 1358.150 719.130 1358.450 ;
        RECT 717.870 1358.140 718.250 1358.150 ;
        RECT 718.830 1354.370 719.130 1358.150 ;
        RECT 716.070 1354.070 719.130 1354.370 ;
        RECT 716.070 1353.010 716.370 1354.070 ;
        RECT 717.205 1353.010 717.535 1353.025 ;
        RECT 716.070 1352.710 717.535 1353.010 ;
        RECT 717.205 1352.695 717.535 1352.710 ;
        RECT 721.345 1325.130 721.675 1325.145 ;
        RECT 733.510 1325.130 733.890 1325.140 ;
        RECT 721.345 1324.830 733.890 1325.130 ;
        RECT 721.345 1324.815 721.675 1324.830 ;
        RECT 733.510 1324.820 733.890 1324.830 ;
        RECT 876.110 14.770 876.490 14.780 ;
        RECT 876.825 14.770 877.155 14.785 ;
        RECT 876.110 14.470 877.155 14.770 ;
        RECT 876.110 14.460 876.490 14.470 ;
        RECT 876.825 14.455 877.155 14.470 ;
      LAYER via3 ;
        RECT 715.140 2392.420 715.460 2392.740 ;
        RECT 715.140 2314.900 715.460 2315.220 ;
        RECT 715.140 2280.220 715.460 2280.540 ;
        RECT 715.140 1859.300 715.460 1859.620 ;
        RECT 715.140 1847.740 715.460 1848.060 ;
        RECT 715.140 1490.740 715.460 1491.060 ;
        RECT 718.820 1490.740 719.140 1491.060 ;
        RECT 717.900 1358.140 718.220 1358.460 ;
        RECT 733.540 1324.820 733.860 1325.140 ;
        RECT 876.140 14.460 876.460 14.780 ;
      LAYER met4 ;
        RECT 715.135 2392.415 715.465 2392.745 ;
        RECT 715.150 2315.225 715.450 2392.415 ;
        RECT 715.135 2314.895 715.465 2315.225 ;
        RECT 715.135 2280.215 715.465 2280.545 ;
        RECT 715.150 1859.625 715.450 2280.215 ;
        RECT 715.135 1859.295 715.465 1859.625 ;
        RECT 715.135 1847.735 715.465 1848.065 ;
        RECT 715.150 1491.065 715.450 1847.735 ;
        RECT 715.135 1490.735 715.465 1491.065 ;
        RECT 718.815 1491.050 719.145 1491.065 ;
        RECT 718.815 1490.750 720.050 1491.050 ;
        RECT 718.815 1490.735 719.145 1490.750 ;
        RECT 719.750 1488.090 720.050 1490.750 ;
        RECT 724.350 1489.390 727.410 1489.690 ;
        RECT 724.350 1488.090 724.650 1489.390 ;
        RECT 719.310 1486.910 720.490 1488.090 ;
        RECT 723.910 1486.910 725.090 1488.090 ;
        RECT 727.110 1382.250 727.410 1489.390 ;
        RECT 721.590 1381.950 727.410 1382.250 ;
        RECT 721.590 1372.730 721.890 1381.950 ;
        RECT 717.910 1372.430 721.890 1372.730 ;
        RECT 717.910 1358.465 718.210 1372.430 ;
        RECT 717.895 1358.135 718.225 1358.465 ;
        RECT 733.110 1330.510 734.290 1331.690 ;
        RECT 875.710 1330.510 876.890 1331.690 ;
        RECT 733.550 1325.145 733.850 1330.510 ;
        RECT 733.535 1324.815 733.865 1325.145 ;
        RECT 876.150 14.785 876.450 1330.510 ;
        RECT 876.135 14.455 876.465 14.785 ;
      LAYER met5 ;
        RECT 719.100 1486.700 725.300 1488.300 ;
        RECT 732.900 1330.300 877.100 1331.900 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 896.685 531.505 896.855 579.615 ;
        RECT 896.685 435.285 896.855 483.055 ;
        RECT 896.685 386.325 896.855 434.775 ;
        RECT 896.685 48.365 896.855 96.475 ;
      LAYER mcon ;
        RECT 896.685 579.445 896.855 579.615 ;
        RECT 896.685 482.885 896.855 483.055 ;
        RECT 896.685 434.605 896.855 434.775 ;
        RECT 896.685 96.305 896.855 96.475 ;
      LAYER met1 ;
        RECT 896.610 1314.000 896.930 1314.060 ;
        RECT 1563.150 1314.000 1563.470 1314.060 ;
        RECT 896.610 1313.860 1563.470 1314.000 ;
        RECT 896.610 1313.800 896.930 1313.860 ;
        RECT 1563.150 1313.800 1563.470 1313.860 ;
        RECT 896.610 1256.680 896.930 1256.940 ;
        RECT 896.700 1256.260 896.840 1256.680 ;
        RECT 896.610 1256.000 896.930 1256.260 ;
        RECT 896.610 1207.580 896.930 1207.640 ;
        RECT 897.530 1207.580 897.850 1207.640 ;
        RECT 896.610 1207.440 897.850 1207.580 ;
        RECT 896.610 1207.380 896.930 1207.440 ;
        RECT 897.530 1207.380 897.850 1207.440 ;
        RECT 896.610 1111.020 896.930 1111.080 ;
        RECT 897.530 1111.020 897.850 1111.080 ;
        RECT 896.610 1110.880 897.850 1111.020 ;
        RECT 896.610 1110.820 896.930 1110.880 ;
        RECT 897.530 1110.820 897.850 1110.880 ;
        RECT 896.610 1014.460 896.930 1014.520 ;
        RECT 897.530 1014.460 897.850 1014.520 ;
        RECT 896.610 1014.320 897.850 1014.460 ;
        RECT 896.610 1014.260 896.930 1014.320 ;
        RECT 897.530 1014.260 897.850 1014.320 ;
        RECT 896.610 917.900 896.930 917.960 ;
        RECT 897.530 917.900 897.850 917.960 ;
        RECT 896.610 917.760 897.850 917.900 ;
        RECT 896.610 917.700 896.930 917.760 ;
        RECT 897.530 917.700 897.850 917.760 ;
        RECT 896.610 772.720 896.930 772.780 ;
        RECT 897.530 772.720 897.850 772.780 ;
        RECT 896.610 772.580 897.850 772.720 ;
        RECT 896.610 772.520 896.930 772.580 ;
        RECT 897.530 772.520 897.850 772.580 ;
        RECT 896.610 676.160 896.930 676.220 ;
        RECT 897.530 676.160 897.850 676.220 ;
        RECT 896.610 676.020 897.850 676.160 ;
        RECT 896.610 675.960 896.930 676.020 ;
        RECT 897.530 675.960 897.850 676.020 ;
        RECT 896.610 579.600 896.930 579.660 ;
        RECT 896.415 579.460 896.930 579.600 ;
        RECT 896.610 579.400 896.930 579.460 ;
        RECT 896.610 531.660 896.930 531.720 ;
        RECT 896.415 531.520 896.930 531.660 ;
        RECT 896.610 531.460 896.930 531.520 ;
        RECT 896.610 483.040 896.930 483.100 ;
        RECT 896.415 482.900 896.930 483.040 ;
        RECT 896.610 482.840 896.930 482.900 ;
        RECT 896.610 435.440 896.930 435.500 ;
        RECT 896.415 435.300 896.930 435.440 ;
        RECT 896.610 435.240 896.930 435.300 ;
        RECT 896.610 434.760 896.930 434.820 ;
        RECT 896.415 434.620 896.930 434.760 ;
        RECT 896.610 434.560 896.930 434.620 ;
        RECT 896.610 386.480 896.930 386.540 ;
        RECT 896.415 386.340 896.930 386.480 ;
        RECT 896.610 386.280 896.930 386.340 ;
        RECT 896.610 96.460 896.930 96.520 ;
        RECT 896.415 96.320 896.930 96.460 ;
        RECT 896.610 96.260 896.930 96.320 ;
        RECT 896.610 48.520 896.930 48.580 ;
        RECT 896.415 48.380 896.930 48.520 ;
        RECT 896.610 48.320 896.930 48.380 ;
        RECT 894.770 2.960 895.090 3.020 ;
        RECT 897.530 2.960 897.850 3.020 ;
        RECT 894.770 2.820 897.850 2.960 ;
        RECT 894.770 2.760 895.090 2.820 ;
        RECT 897.530 2.760 897.850 2.820 ;
      LAYER via ;
        RECT 896.640 1313.800 896.900 1314.060 ;
        RECT 1563.180 1313.800 1563.440 1314.060 ;
        RECT 896.640 1256.680 896.900 1256.940 ;
        RECT 896.640 1256.000 896.900 1256.260 ;
        RECT 896.640 1207.380 896.900 1207.640 ;
        RECT 897.560 1207.380 897.820 1207.640 ;
        RECT 896.640 1110.820 896.900 1111.080 ;
        RECT 897.560 1110.820 897.820 1111.080 ;
        RECT 896.640 1014.260 896.900 1014.520 ;
        RECT 897.560 1014.260 897.820 1014.520 ;
        RECT 896.640 917.700 896.900 917.960 ;
        RECT 897.560 917.700 897.820 917.960 ;
        RECT 896.640 772.520 896.900 772.780 ;
        RECT 897.560 772.520 897.820 772.780 ;
        RECT 896.640 675.960 896.900 676.220 ;
        RECT 897.560 675.960 897.820 676.220 ;
        RECT 896.640 579.400 896.900 579.660 ;
        RECT 896.640 531.460 896.900 531.720 ;
        RECT 896.640 482.840 896.900 483.100 ;
        RECT 896.640 435.240 896.900 435.500 ;
        RECT 896.640 434.560 896.900 434.820 ;
        RECT 896.640 386.280 896.900 386.540 ;
        RECT 896.640 96.260 896.900 96.520 ;
        RECT 896.640 48.320 896.900 48.580 ;
        RECT 894.800 2.760 895.060 3.020 ;
        RECT 897.560 2.760 897.820 3.020 ;
      LAYER met2 ;
        RECT 1563.220 1323.135 1563.500 1327.135 ;
        RECT 1563.240 1314.090 1563.380 1323.135 ;
        RECT 896.640 1313.770 896.900 1314.090 ;
        RECT 1563.180 1313.770 1563.440 1314.090 ;
        RECT 896.700 1256.970 896.840 1313.770 ;
        RECT 896.640 1256.650 896.900 1256.970 ;
        RECT 896.640 1255.970 896.900 1256.290 ;
        RECT 896.700 1255.805 896.840 1255.970 ;
        RECT 896.630 1255.435 896.910 1255.805 ;
        RECT 897.550 1255.435 897.830 1255.805 ;
        RECT 897.620 1207.670 897.760 1255.435 ;
        RECT 896.640 1207.350 896.900 1207.670 ;
        RECT 897.560 1207.350 897.820 1207.670 ;
        RECT 896.700 1159.245 896.840 1207.350 ;
        RECT 896.630 1158.875 896.910 1159.245 ;
        RECT 897.550 1158.875 897.830 1159.245 ;
        RECT 897.620 1111.110 897.760 1158.875 ;
        RECT 896.640 1110.790 896.900 1111.110 ;
        RECT 897.560 1110.790 897.820 1111.110 ;
        RECT 896.700 1062.685 896.840 1110.790 ;
        RECT 896.630 1062.315 896.910 1062.685 ;
        RECT 897.550 1062.315 897.830 1062.685 ;
        RECT 897.620 1014.550 897.760 1062.315 ;
        RECT 896.640 1014.230 896.900 1014.550 ;
        RECT 897.560 1014.230 897.820 1014.550 ;
        RECT 896.700 966.125 896.840 1014.230 ;
        RECT 896.630 965.755 896.910 966.125 ;
        RECT 897.550 965.755 897.830 966.125 ;
        RECT 897.620 917.990 897.760 965.755 ;
        RECT 896.640 917.670 896.900 917.990 ;
        RECT 897.560 917.670 897.820 917.990 ;
        RECT 896.700 869.565 896.840 917.670 ;
        RECT 896.630 869.195 896.910 869.565 ;
        RECT 897.550 869.195 897.830 869.565 ;
        RECT 897.620 821.285 897.760 869.195 ;
        RECT 896.630 820.915 896.910 821.285 ;
        RECT 897.550 820.915 897.830 821.285 ;
        RECT 896.700 772.810 896.840 820.915 ;
        RECT 896.640 772.490 896.900 772.810 ;
        RECT 897.560 772.490 897.820 772.810 ;
        RECT 897.620 724.725 897.760 772.490 ;
        RECT 896.630 724.355 896.910 724.725 ;
        RECT 897.550 724.355 897.830 724.725 ;
        RECT 896.700 676.250 896.840 724.355 ;
        RECT 896.640 675.930 896.900 676.250 ;
        RECT 897.560 675.930 897.820 676.250 ;
        RECT 897.620 628.165 897.760 675.930 ;
        RECT 896.630 627.795 896.910 628.165 ;
        RECT 897.550 627.795 897.830 628.165 ;
        RECT 896.700 579.690 896.840 627.795 ;
        RECT 896.640 579.370 896.900 579.690 ;
        RECT 896.640 531.430 896.900 531.750 ;
        RECT 896.700 483.130 896.840 531.430 ;
        RECT 896.640 482.810 896.900 483.130 ;
        RECT 896.640 435.210 896.900 435.530 ;
        RECT 896.700 434.850 896.840 435.210 ;
        RECT 896.640 434.530 896.900 434.850 ;
        RECT 896.640 386.250 896.900 386.570 ;
        RECT 896.700 96.550 896.840 386.250 ;
        RECT 896.640 96.230 896.900 96.550 ;
        RECT 896.640 48.290 896.900 48.610 ;
        RECT 896.700 41.325 896.840 48.290 ;
        RECT 896.630 40.955 896.910 41.325 ;
        RECT 897.550 40.955 897.830 41.325 ;
        RECT 897.620 3.050 897.760 40.955 ;
        RECT 894.800 2.730 895.060 3.050 ;
        RECT 897.560 2.730 897.820 3.050 ;
        RECT 894.860 2.400 895.000 2.730 ;
        RECT 894.650 -4.800 895.210 2.400 ;
      LAYER via2 ;
        RECT 896.630 1255.480 896.910 1255.760 ;
        RECT 897.550 1255.480 897.830 1255.760 ;
        RECT 896.630 1158.920 896.910 1159.200 ;
        RECT 897.550 1158.920 897.830 1159.200 ;
        RECT 896.630 1062.360 896.910 1062.640 ;
        RECT 897.550 1062.360 897.830 1062.640 ;
        RECT 896.630 965.800 896.910 966.080 ;
        RECT 897.550 965.800 897.830 966.080 ;
        RECT 896.630 869.240 896.910 869.520 ;
        RECT 897.550 869.240 897.830 869.520 ;
        RECT 896.630 820.960 896.910 821.240 ;
        RECT 897.550 820.960 897.830 821.240 ;
        RECT 896.630 724.400 896.910 724.680 ;
        RECT 897.550 724.400 897.830 724.680 ;
        RECT 896.630 627.840 896.910 628.120 ;
        RECT 897.550 627.840 897.830 628.120 ;
        RECT 896.630 41.000 896.910 41.280 ;
        RECT 897.550 41.000 897.830 41.280 ;
      LAYER met3 ;
        RECT 896.605 1255.770 896.935 1255.785 ;
        RECT 897.525 1255.770 897.855 1255.785 ;
        RECT 896.605 1255.470 897.855 1255.770 ;
        RECT 896.605 1255.455 896.935 1255.470 ;
        RECT 897.525 1255.455 897.855 1255.470 ;
        RECT 896.605 1159.210 896.935 1159.225 ;
        RECT 897.525 1159.210 897.855 1159.225 ;
        RECT 896.605 1158.910 897.855 1159.210 ;
        RECT 896.605 1158.895 896.935 1158.910 ;
        RECT 897.525 1158.895 897.855 1158.910 ;
        RECT 896.605 1062.650 896.935 1062.665 ;
        RECT 897.525 1062.650 897.855 1062.665 ;
        RECT 896.605 1062.350 897.855 1062.650 ;
        RECT 896.605 1062.335 896.935 1062.350 ;
        RECT 897.525 1062.335 897.855 1062.350 ;
        RECT 896.605 966.090 896.935 966.105 ;
        RECT 897.525 966.090 897.855 966.105 ;
        RECT 896.605 965.790 897.855 966.090 ;
        RECT 896.605 965.775 896.935 965.790 ;
        RECT 897.525 965.775 897.855 965.790 ;
        RECT 896.605 869.530 896.935 869.545 ;
        RECT 897.525 869.530 897.855 869.545 ;
        RECT 896.605 869.230 897.855 869.530 ;
        RECT 896.605 869.215 896.935 869.230 ;
        RECT 897.525 869.215 897.855 869.230 ;
        RECT 896.605 821.250 896.935 821.265 ;
        RECT 897.525 821.250 897.855 821.265 ;
        RECT 896.605 820.950 897.855 821.250 ;
        RECT 896.605 820.935 896.935 820.950 ;
        RECT 897.525 820.935 897.855 820.950 ;
        RECT 896.605 724.690 896.935 724.705 ;
        RECT 897.525 724.690 897.855 724.705 ;
        RECT 896.605 724.390 897.855 724.690 ;
        RECT 896.605 724.375 896.935 724.390 ;
        RECT 897.525 724.375 897.855 724.390 ;
        RECT 896.605 628.130 896.935 628.145 ;
        RECT 897.525 628.130 897.855 628.145 ;
        RECT 896.605 627.830 897.855 628.130 ;
        RECT 896.605 627.815 896.935 627.830 ;
        RECT 897.525 627.815 897.855 627.830 ;
        RECT 896.605 41.290 896.935 41.305 ;
        RECT 897.525 41.290 897.855 41.305 ;
        RECT 896.605 40.990 897.855 41.290 ;
        RECT 896.605 40.975 896.935 40.990 ;
        RECT 897.525 40.975 897.855 40.990 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1754.585 1558.985 1755.215 1559.155 ;
        RECT 1755.045 1472.285 1755.215 1558.985 ;
      LAYER met1 ;
        RECT 1754.510 1587.360 1754.830 1587.420 ;
        RECT 1758.190 1587.360 1758.510 1587.420 ;
        RECT 1754.510 1587.220 1758.510 1587.360 ;
        RECT 1754.510 1587.160 1754.830 1587.220 ;
        RECT 1758.190 1587.160 1758.510 1587.220 ;
        RECT 1754.510 1559.140 1754.830 1559.200 ;
        RECT 1754.315 1559.000 1754.830 1559.140 ;
        RECT 1754.510 1558.940 1754.830 1559.000 ;
        RECT 1754.510 1472.440 1754.830 1472.500 ;
        RECT 1754.985 1472.440 1755.275 1472.485 ;
        RECT 1754.510 1472.300 1755.275 1472.440 ;
        RECT 1754.510 1472.240 1754.830 1472.300 ;
        RECT 1754.985 1472.255 1755.275 1472.300 ;
        RECT 1754.510 1422.460 1754.830 1422.520 ;
        RECT 1754.510 1422.320 1755.200 1422.460 ;
        RECT 1754.510 1422.260 1754.830 1422.320 ;
        RECT 1754.510 1421.100 1754.830 1421.160 ;
        RECT 1755.060 1421.100 1755.200 1422.320 ;
        RECT 1754.510 1420.960 1755.200 1421.100 ;
        RECT 1754.510 1420.900 1754.830 1420.960 ;
        RECT 917.310 67.220 917.630 67.280 ;
        RECT 1754.510 67.220 1754.830 67.280 ;
        RECT 917.310 67.080 1754.830 67.220 ;
        RECT 917.310 67.020 917.630 67.080 ;
        RECT 1754.510 67.020 1754.830 67.080 ;
        RECT 912.710 20.640 913.030 20.700 ;
        RECT 917.310 20.640 917.630 20.700 ;
        RECT 912.710 20.500 917.630 20.640 ;
        RECT 912.710 20.440 913.030 20.500 ;
        RECT 917.310 20.440 917.630 20.500 ;
      LAYER via ;
        RECT 1754.540 1587.160 1754.800 1587.420 ;
        RECT 1758.220 1587.160 1758.480 1587.420 ;
        RECT 1754.540 1558.940 1754.800 1559.200 ;
        RECT 1754.540 1472.240 1754.800 1472.500 ;
        RECT 1754.540 1422.260 1754.800 1422.520 ;
        RECT 1754.540 1420.900 1754.800 1421.160 ;
        RECT 917.340 67.020 917.600 67.280 ;
        RECT 1754.540 67.020 1754.800 67.280 ;
        RECT 912.740 20.440 913.000 20.700 ;
        RECT 917.340 20.440 917.600 20.700 ;
      LAYER met2 ;
        RECT 1758.210 1587.955 1758.490 1588.325 ;
        RECT 1758.280 1587.450 1758.420 1587.955 ;
        RECT 1754.540 1587.130 1754.800 1587.450 ;
        RECT 1758.220 1587.130 1758.480 1587.450 ;
        RECT 1754.600 1559.230 1754.740 1587.130 ;
        RECT 1754.540 1558.910 1754.800 1559.230 ;
        RECT 1754.540 1472.210 1754.800 1472.530 ;
        RECT 1754.600 1422.550 1754.740 1472.210 ;
        RECT 1754.540 1422.230 1754.800 1422.550 ;
        RECT 1754.540 1420.870 1754.800 1421.190 ;
        RECT 1754.600 67.310 1754.740 1420.870 ;
        RECT 917.340 66.990 917.600 67.310 ;
        RECT 1754.540 66.990 1754.800 67.310 ;
        RECT 917.400 20.730 917.540 66.990 ;
        RECT 912.740 20.410 913.000 20.730 ;
        RECT 917.340 20.410 917.600 20.730 ;
        RECT 912.800 2.400 912.940 20.410 ;
        RECT 912.590 -4.800 913.150 2.400 ;
      LAYER via2 ;
        RECT 1758.210 1588.000 1758.490 1588.280 ;
      LAYER met3 ;
        RECT 1758.185 1588.290 1758.515 1588.305 ;
        RECT 1758.185 1587.975 1758.730 1588.290 ;
        RECT 1758.430 1587.615 1758.730 1587.975 ;
        RECT 1755.835 1587.015 1759.835 1587.615 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1754.585 1421.625 1754.755 1545.215 ;
        RECT 1754.125 669.545 1754.295 717.655 ;
        RECT 1754.125 476.085 1754.295 524.195 ;
        RECT 1754.125 379.525 1754.295 427.635 ;
        RECT 1753.665 186.405 1753.835 234.515 ;
        RECT 1753.205 83.045 1753.375 97.155 ;
      LAYER mcon ;
        RECT 1754.585 1545.045 1754.755 1545.215 ;
        RECT 1754.125 717.485 1754.295 717.655 ;
        RECT 1754.125 524.025 1754.295 524.195 ;
        RECT 1754.125 427.465 1754.295 427.635 ;
        RECT 1753.665 234.345 1753.835 234.515 ;
        RECT 1753.205 96.985 1753.375 97.155 ;
      LAYER met1 ;
        RECT 1754.510 1594.160 1754.830 1594.220 ;
        RECT 1759.110 1594.160 1759.430 1594.220 ;
        RECT 1754.510 1594.020 1759.430 1594.160 ;
        RECT 1754.510 1593.960 1754.830 1594.020 ;
        RECT 1759.110 1593.960 1759.430 1594.020 ;
        RECT 1754.510 1545.200 1754.830 1545.260 ;
        RECT 1754.315 1545.060 1754.830 1545.200 ;
        RECT 1754.510 1545.000 1754.830 1545.060 ;
        RECT 1754.510 1421.780 1754.830 1421.840 ;
        RECT 1754.315 1421.640 1754.830 1421.780 ;
        RECT 1754.510 1421.580 1754.830 1421.640 ;
        RECT 1754.050 1307.200 1754.370 1307.260 ;
        RECT 1755.430 1307.200 1755.750 1307.260 ;
        RECT 1754.050 1307.060 1755.750 1307.200 ;
        RECT 1754.050 1307.000 1754.370 1307.060 ;
        RECT 1755.430 1307.000 1755.750 1307.060 ;
        RECT 1754.050 1245.660 1754.370 1245.720 ;
        RECT 1755.430 1245.660 1755.750 1245.720 ;
        RECT 1754.050 1245.520 1755.750 1245.660 ;
        RECT 1754.050 1245.460 1754.370 1245.520 ;
        RECT 1755.430 1245.460 1755.750 1245.520 ;
        RECT 1754.050 909.740 1754.370 909.800 ;
        RECT 1755.430 909.740 1755.750 909.800 ;
        RECT 1754.050 909.600 1755.750 909.740 ;
        RECT 1754.050 909.540 1754.370 909.600 ;
        RECT 1755.430 909.540 1755.750 909.600 ;
        RECT 1754.050 831.200 1754.370 831.260 ;
        RECT 1755.430 831.200 1755.750 831.260 ;
        RECT 1754.050 831.060 1755.750 831.200 ;
        RECT 1754.050 831.000 1754.370 831.060 ;
        RECT 1755.430 831.000 1755.750 831.060 ;
        RECT 1754.050 814.200 1754.370 814.260 ;
        RECT 1755.430 814.200 1755.750 814.260 ;
        RECT 1754.050 814.060 1755.750 814.200 ;
        RECT 1754.050 814.000 1754.370 814.060 ;
        RECT 1755.430 814.000 1755.750 814.060 ;
        RECT 1754.050 717.640 1754.370 717.700 ;
        RECT 1753.855 717.500 1754.370 717.640 ;
        RECT 1754.050 717.440 1754.370 717.500 ;
        RECT 1754.050 669.700 1754.370 669.760 ;
        RECT 1753.855 669.560 1754.370 669.700 ;
        RECT 1754.050 669.500 1754.370 669.560 ;
        RECT 1754.050 524.180 1754.370 524.240 ;
        RECT 1753.855 524.040 1754.370 524.180 ;
        RECT 1754.050 523.980 1754.370 524.040 ;
        RECT 1754.050 476.240 1754.370 476.300 ;
        RECT 1753.855 476.100 1754.370 476.240 ;
        RECT 1754.050 476.040 1754.370 476.100 ;
        RECT 1754.050 427.620 1754.370 427.680 ;
        RECT 1753.855 427.480 1754.370 427.620 ;
        RECT 1754.050 427.420 1754.370 427.480 ;
        RECT 1754.050 379.680 1754.370 379.740 ;
        RECT 1753.855 379.540 1754.370 379.680 ;
        RECT 1754.050 379.480 1754.370 379.540 ;
        RECT 1753.605 234.500 1753.895 234.545 ;
        RECT 1754.050 234.500 1754.370 234.560 ;
        RECT 1753.605 234.360 1754.370 234.500 ;
        RECT 1753.605 234.315 1753.895 234.360 ;
        RECT 1754.050 234.300 1754.370 234.360 ;
        RECT 1753.605 186.560 1753.895 186.605 ;
        RECT 1754.050 186.560 1754.370 186.620 ;
        RECT 1753.605 186.420 1754.370 186.560 ;
        RECT 1753.605 186.375 1753.895 186.420 ;
        RECT 1754.050 186.360 1754.370 186.420 ;
        RECT 1754.050 159.360 1754.370 159.420 ;
        RECT 1753.220 159.220 1754.370 159.360 ;
        RECT 1753.220 158.740 1753.360 159.220 ;
        RECT 1754.050 159.160 1754.370 159.220 ;
        RECT 1753.130 158.480 1753.450 158.740 ;
        RECT 1753.130 97.140 1753.450 97.200 ;
        RECT 1752.935 97.000 1753.450 97.140 ;
        RECT 1753.130 96.940 1753.450 97.000 ;
        RECT 1753.130 83.200 1753.450 83.260 ;
        RECT 1752.935 83.060 1753.450 83.200 ;
        RECT 1753.130 83.000 1753.450 83.060 ;
        RECT 931.110 67.560 931.430 67.620 ;
        RECT 1753.130 67.560 1753.450 67.620 ;
        RECT 931.110 67.420 1753.450 67.560 ;
        RECT 931.110 67.360 931.430 67.420 ;
        RECT 1753.130 67.360 1753.450 67.420 ;
      LAYER via ;
        RECT 1754.540 1593.960 1754.800 1594.220 ;
        RECT 1759.140 1593.960 1759.400 1594.220 ;
        RECT 1754.540 1545.000 1754.800 1545.260 ;
        RECT 1754.540 1421.580 1754.800 1421.840 ;
        RECT 1754.080 1307.000 1754.340 1307.260 ;
        RECT 1755.460 1307.000 1755.720 1307.260 ;
        RECT 1754.080 1245.460 1754.340 1245.720 ;
        RECT 1755.460 1245.460 1755.720 1245.720 ;
        RECT 1754.080 909.540 1754.340 909.800 ;
        RECT 1755.460 909.540 1755.720 909.800 ;
        RECT 1754.080 831.000 1754.340 831.260 ;
        RECT 1755.460 831.000 1755.720 831.260 ;
        RECT 1754.080 814.000 1754.340 814.260 ;
        RECT 1755.460 814.000 1755.720 814.260 ;
        RECT 1754.080 717.440 1754.340 717.700 ;
        RECT 1754.080 669.500 1754.340 669.760 ;
        RECT 1754.080 523.980 1754.340 524.240 ;
        RECT 1754.080 476.040 1754.340 476.300 ;
        RECT 1754.080 427.420 1754.340 427.680 ;
        RECT 1754.080 379.480 1754.340 379.740 ;
        RECT 1754.080 234.300 1754.340 234.560 ;
        RECT 1754.080 186.360 1754.340 186.620 ;
        RECT 1754.080 159.160 1754.340 159.420 ;
        RECT 1753.160 158.480 1753.420 158.740 ;
        RECT 1753.160 96.940 1753.420 97.200 ;
        RECT 1753.160 83.000 1753.420 83.260 ;
        RECT 931.140 67.360 931.400 67.620 ;
        RECT 1753.160 67.360 1753.420 67.620 ;
      LAYER met2 ;
        RECT 1759.130 1626.715 1759.410 1627.085 ;
        RECT 1759.200 1594.250 1759.340 1626.715 ;
        RECT 1754.540 1593.930 1754.800 1594.250 ;
        RECT 1759.140 1593.930 1759.400 1594.250 ;
        RECT 1754.600 1588.210 1754.740 1593.930 ;
        RECT 1754.140 1588.070 1754.740 1588.210 ;
        RECT 1754.140 1545.370 1754.280 1588.070 ;
        RECT 1754.140 1545.290 1754.740 1545.370 ;
        RECT 1754.140 1545.230 1754.800 1545.290 ;
        RECT 1754.540 1544.970 1754.800 1545.230 ;
        RECT 1754.540 1421.780 1754.800 1421.870 ;
        RECT 1754.140 1421.640 1754.800 1421.780 ;
        RECT 1754.140 1307.290 1754.280 1421.640 ;
        RECT 1754.540 1421.550 1754.800 1421.640 ;
        RECT 1754.080 1306.970 1754.340 1307.290 ;
        RECT 1755.460 1306.970 1755.720 1307.290 ;
        RECT 1755.520 1245.750 1755.660 1306.970 ;
        RECT 1754.080 1245.430 1754.340 1245.750 ;
        RECT 1755.460 1245.430 1755.720 1245.750 ;
        RECT 1754.140 909.830 1754.280 1245.430 ;
        RECT 1754.080 909.510 1754.340 909.830 ;
        RECT 1755.460 909.510 1755.720 909.830 ;
        RECT 1755.520 831.290 1755.660 909.510 ;
        RECT 1754.080 830.970 1754.340 831.290 ;
        RECT 1755.460 830.970 1755.720 831.290 ;
        RECT 1754.140 814.290 1754.280 830.970 ;
        RECT 1754.080 813.970 1754.340 814.290 ;
        RECT 1755.460 813.970 1755.720 814.290 ;
        RECT 1755.520 766.205 1755.660 813.970 ;
        RECT 1754.070 765.835 1754.350 766.205 ;
        RECT 1755.450 765.835 1755.730 766.205 ;
        RECT 1754.140 725.405 1754.280 765.835 ;
        RECT 1754.070 725.035 1754.350 725.405 ;
        RECT 1754.070 724.355 1754.350 724.725 ;
        RECT 1754.140 717.730 1754.280 724.355 ;
        RECT 1754.080 717.410 1754.340 717.730 ;
        RECT 1754.080 669.470 1754.340 669.790 ;
        RECT 1754.140 628.845 1754.280 669.470 ;
        RECT 1754.070 628.475 1754.350 628.845 ;
        RECT 1754.070 627.795 1754.350 628.165 ;
        RECT 1754.140 524.270 1754.280 627.795 ;
        RECT 1754.080 523.950 1754.340 524.270 ;
        RECT 1754.080 476.010 1754.340 476.330 ;
        RECT 1754.140 427.710 1754.280 476.010 ;
        RECT 1754.080 427.390 1754.340 427.710 ;
        RECT 1754.080 379.450 1754.340 379.770 ;
        RECT 1754.140 234.590 1754.280 379.450 ;
        RECT 1754.080 234.270 1754.340 234.590 ;
        RECT 1754.080 186.330 1754.340 186.650 ;
        RECT 1754.140 159.450 1754.280 186.330 ;
        RECT 1754.080 159.130 1754.340 159.450 ;
        RECT 1753.160 158.450 1753.420 158.770 ;
        RECT 1753.220 97.230 1753.360 158.450 ;
        RECT 1753.160 96.910 1753.420 97.230 ;
        RECT 1753.160 82.970 1753.420 83.290 ;
        RECT 1753.220 67.650 1753.360 82.970 ;
        RECT 931.140 67.330 931.400 67.650 ;
        RECT 1753.160 67.330 1753.420 67.650 ;
        RECT 931.200 14.010 931.340 67.330 ;
        RECT 930.740 13.870 931.340 14.010 ;
        RECT 930.740 13.330 930.880 13.870 ;
        RECT 930.280 13.190 930.880 13.330 ;
        RECT 930.280 2.400 930.420 13.190 ;
        RECT 930.070 -4.800 930.630 2.400 ;
      LAYER via2 ;
        RECT 1759.130 1626.760 1759.410 1627.040 ;
        RECT 1754.070 765.880 1754.350 766.160 ;
        RECT 1755.450 765.880 1755.730 766.160 ;
        RECT 1754.070 725.080 1754.350 725.360 ;
        RECT 1754.070 724.400 1754.350 724.680 ;
        RECT 1754.070 628.520 1754.350 628.800 ;
        RECT 1754.070 627.840 1754.350 628.120 ;
      LAYER met3 ;
        RECT 1755.835 1629.175 1759.835 1629.775 ;
        RECT 1759.350 1627.065 1759.650 1629.175 ;
        RECT 1759.105 1626.750 1759.650 1627.065 ;
        RECT 1759.105 1626.735 1759.435 1626.750 ;
        RECT 1754.045 766.170 1754.375 766.185 ;
        RECT 1755.425 766.170 1755.755 766.185 ;
        RECT 1754.045 765.870 1755.755 766.170 ;
        RECT 1754.045 765.855 1754.375 765.870 ;
        RECT 1755.425 765.855 1755.755 765.870 ;
        RECT 1754.045 725.370 1754.375 725.385 ;
        RECT 1753.830 725.055 1754.375 725.370 ;
        RECT 1753.830 724.705 1754.130 725.055 ;
        RECT 1753.830 724.390 1754.375 724.705 ;
        RECT 1754.045 724.375 1754.375 724.390 ;
        RECT 1754.045 628.810 1754.375 628.825 ;
        RECT 1753.830 628.495 1754.375 628.810 ;
        RECT 1753.830 628.145 1754.130 628.495 ;
        RECT 1753.830 627.830 1754.375 628.145 ;
        RECT 1754.045 627.815 1754.375 627.830 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 951.810 148.140 952.130 148.200 ;
        RECT 1760.490 148.140 1760.810 148.200 ;
        RECT 951.810 148.000 1760.810 148.140 ;
        RECT 951.810 147.940 952.130 148.000 ;
        RECT 1760.490 147.940 1760.810 148.000 ;
        RECT 948.130 20.640 948.450 20.700 ;
        RECT 951.810 20.640 952.130 20.700 ;
        RECT 948.130 20.500 952.130 20.640 ;
        RECT 948.130 20.440 948.450 20.500 ;
        RECT 951.810 20.440 952.130 20.500 ;
      LAYER via ;
        RECT 951.840 147.940 952.100 148.200 ;
        RECT 1760.520 147.940 1760.780 148.200 ;
        RECT 948.160 20.440 948.420 20.700 ;
        RECT 951.840 20.440 952.100 20.700 ;
      LAYER met2 ;
        RECT 1760.510 2091.835 1760.790 2092.205 ;
        RECT 1760.580 148.230 1760.720 2091.835 ;
        RECT 951.840 147.910 952.100 148.230 ;
        RECT 1760.520 147.910 1760.780 148.230 ;
        RECT 951.900 20.730 952.040 147.910 ;
        RECT 948.160 20.410 948.420 20.730 ;
        RECT 951.840 20.410 952.100 20.730 ;
        RECT 948.220 2.400 948.360 20.410 ;
        RECT 948.010 -4.800 948.570 2.400 ;
      LAYER via2 ;
        RECT 1760.510 2091.880 1760.790 2092.160 ;
      LAYER met3 ;
        RECT 1755.835 2092.170 1759.835 2092.175 ;
        RECT 1760.485 2092.170 1760.815 2092.185 ;
        RECT 1755.835 2091.870 1760.815 2092.170 ;
        RECT 1755.835 2091.575 1759.835 2091.870 ;
        RECT 1760.485 2091.855 1760.815 2091.870 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 967.525 1326.425 967.695 1330.675 ;
        RECT 966.605 48.365 966.775 65.195 ;
      LAYER mcon ;
        RECT 967.525 1330.505 967.695 1330.675 ;
        RECT 966.605 65.025 966.775 65.195 ;
      LAYER met1 ;
        RECT 698.810 2390.100 699.130 2390.160 ;
        RECT 1323.030 2390.100 1323.350 2390.160 ;
        RECT 698.810 2389.960 1323.350 2390.100 ;
        RECT 698.810 2389.900 699.130 2389.960 ;
        RECT 1323.030 2389.900 1323.350 2389.960 ;
        RECT 698.810 1330.660 699.130 1330.720 ;
        RECT 967.465 1330.660 967.755 1330.705 ;
        RECT 698.810 1330.520 967.755 1330.660 ;
        RECT 698.810 1330.460 699.130 1330.520 ;
        RECT 967.465 1330.475 967.755 1330.520 ;
        RECT 967.450 1326.580 967.770 1326.640 ;
        RECT 967.255 1326.440 967.770 1326.580 ;
        RECT 967.450 1326.380 967.770 1326.440 ;
        RECT 966.545 65.180 966.835 65.225 ;
        RECT 967.450 65.180 967.770 65.240 ;
        RECT 966.545 65.040 967.770 65.180 ;
        RECT 966.545 64.995 966.835 65.040 ;
        RECT 967.450 64.980 967.770 65.040 ;
        RECT 966.530 48.520 966.850 48.580 ;
        RECT 966.335 48.380 966.850 48.520 ;
        RECT 966.530 48.320 966.850 48.380 ;
      LAYER via ;
        RECT 698.840 2389.900 699.100 2390.160 ;
        RECT 1323.060 2389.900 1323.320 2390.160 ;
        RECT 698.840 1330.460 699.100 1330.720 ;
        RECT 967.480 1326.380 967.740 1326.640 ;
        RECT 967.480 64.980 967.740 65.240 ;
        RECT 966.560 48.320 966.820 48.580 ;
      LAYER met2 ;
        RECT 698.840 2389.870 699.100 2390.190 ;
        RECT 1323.060 2389.870 1323.320 2390.190 ;
        RECT 698.900 1330.750 699.040 2389.870 ;
        RECT 1323.120 2377.880 1323.260 2389.870 ;
        RECT 1323.100 2373.880 1323.380 2377.880 ;
        RECT 698.840 1330.430 699.100 1330.750 ;
        RECT 967.480 1326.350 967.740 1326.670 ;
        RECT 967.540 65.270 967.680 1326.350 ;
        RECT 967.480 64.950 967.740 65.270 ;
        RECT 966.560 48.290 966.820 48.610 ;
        RECT 966.620 24.890 966.760 48.290 ;
        RECT 966.160 24.750 966.760 24.890 ;
        RECT 966.160 2.400 966.300 24.750 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 717.210 1356.160 717.530 1356.220 ;
        RECT 718.590 1356.160 718.910 1356.220 ;
        RECT 717.210 1356.020 718.910 1356.160 ;
        RECT 717.210 1355.960 717.530 1356.020 ;
        RECT 718.590 1355.960 718.910 1356.020 ;
        RECT 717.670 1309.580 717.990 1309.640 ;
        RECT 979.870 1309.580 980.190 1309.640 ;
        RECT 717.670 1309.440 980.190 1309.580 ;
        RECT 717.670 1309.380 717.990 1309.440 ;
        RECT 979.870 1309.380 980.190 1309.440 ;
        RECT 979.870 37.640 980.190 37.700 ;
        RECT 984.010 37.640 984.330 37.700 ;
        RECT 979.870 37.500 984.330 37.640 ;
        RECT 979.870 37.440 980.190 37.500 ;
        RECT 984.010 37.440 984.330 37.500 ;
      LAYER via ;
        RECT 717.240 1355.960 717.500 1356.220 ;
        RECT 718.620 1355.960 718.880 1356.220 ;
        RECT 717.700 1309.380 717.960 1309.640 ;
        RECT 979.900 1309.380 980.160 1309.640 ;
        RECT 979.900 37.440 980.160 37.700 ;
        RECT 984.040 37.440 984.300 37.700 ;
      LAYER met2 ;
        RECT 718.610 1478.475 718.890 1478.845 ;
        RECT 718.680 1356.250 718.820 1478.475 ;
        RECT 717.240 1355.930 717.500 1356.250 ;
        RECT 718.620 1355.930 718.880 1356.250 ;
        RECT 717.300 1354.290 717.440 1355.930 ;
        RECT 717.300 1354.150 717.900 1354.290 ;
        RECT 717.760 1309.670 717.900 1354.150 ;
        RECT 717.700 1309.350 717.960 1309.670 ;
        RECT 979.900 1309.350 980.160 1309.670 ;
        RECT 979.960 37.730 980.100 1309.350 ;
        RECT 979.900 37.410 980.160 37.730 ;
        RECT 984.040 37.410 984.300 37.730 ;
        RECT 984.100 2.400 984.240 37.410 ;
        RECT 983.890 -4.800 984.450 2.400 ;
      LAYER via2 ;
        RECT 718.610 1478.520 718.890 1478.800 ;
      LAYER met3 ;
        RECT 715.810 1480.935 719.810 1481.535 ;
        RECT 718.830 1478.825 719.130 1480.935 ;
        RECT 718.585 1478.510 719.130 1478.825 ;
        RECT 718.585 1478.495 718.915 1478.510 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 668.450 1939.260 668.770 1939.320 ;
        RECT 706.170 1939.260 706.490 1939.320 ;
        RECT 668.450 1939.120 706.490 1939.260 ;
        RECT 668.450 1939.060 668.770 1939.120 ;
        RECT 706.170 1939.060 706.490 1939.120 ;
        RECT 662.930 17.240 663.250 17.300 ;
        RECT 668.450 17.240 668.770 17.300 ;
        RECT 662.930 17.100 668.770 17.240 ;
        RECT 662.930 17.040 663.250 17.100 ;
        RECT 668.450 17.040 668.770 17.100 ;
      LAYER via ;
        RECT 668.480 1939.060 668.740 1939.320 ;
        RECT 706.200 1939.060 706.460 1939.320 ;
        RECT 662.960 17.040 663.220 17.300 ;
        RECT 668.480 17.040 668.740 17.300 ;
      LAYER met2 ;
        RECT 706.190 1942.235 706.470 1942.605 ;
        RECT 706.260 1939.350 706.400 1942.235 ;
        RECT 668.480 1939.030 668.740 1939.350 ;
        RECT 706.200 1939.030 706.460 1939.350 ;
        RECT 668.540 17.330 668.680 1939.030 ;
        RECT 662.960 17.010 663.220 17.330 ;
        RECT 668.480 17.010 668.740 17.330 ;
        RECT 663.020 2.400 663.160 17.010 ;
        RECT 662.810 -4.800 663.370 2.400 ;
      LAYER via2 ;
        RECT 706.190 1942.280 706.470 1942.560 ;
      LAYER met3 ;
        RECT 706.165 1942.570 706.495 1942.585 ;
        RECT 715.810 1942.570 719.810 1942.575 ;
        RECT 706.165 1942.270 719.810 1942.570 ;
        RECT 706.165 1942.255 706.495 1942.270 ;
        RECT 715.810 1941.975 719.810 1942.270 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1007.010 1317.740 1007.330 1317.800 ;
        RECT 1169.390 1317.740 1169.710 1317.800 ;
        RECT 1007.010 1317.600 1169.710 1317.740 ;
        RECT 1007.010 1317.540 1007.330 1317.600 ;
        RECT 1169.390 1317.540 1169.710 1317.600 ;
        RECT 1001.950 14.860 1002.270 14.920 ;
        RECT 1007.010 14.860 1007.330 14.920 ;
        RECT 1001.950 14.720 1007.330 14.860 ;
        RECT 1001.950 14.660 1002.270 14.720 ;
        RECT 1007.010 14.660 1007.330 14.720 ;
      LAYER via ;
        RECT 1007.040 1317.540 1007.300 1317.800 ;
        RECT 1169.420 1317.540 1169.680 1317.800 ;
        RECT 1001.980 14.660 1002.240 14.920 ;
        RECT 1007.040 14.660 1007.300 14.920 ;
      LAYER met2 ;
        RECT 1169.460 1323.135 1169.740 1327.135 ;
        RECT 1169.480 1317.830 1169.620 1323.135 ;
        RECT 1007.040 1317.510 1007.300 1317.830 ;
        RECT 1169.420 1317.510 1169.680 1317.830 ;
        RECT 1007.100 14.950 1007.240 1317.510 ;
        RECT 1001.980 14.630 1002.240 14.950 ;
        RECT 1007.040 14.630 1007.300 14.950 ;
        RECT 1002.040 2.400 1002.180 14.630 ;
        RECT 1001.830 -4.800 1002.390 2.400 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1757.345 1803.785 1757.515 1838.975 ;
      LAYER mcon ;
        RECT 1757.345 1838.805 1757.515 1838.975 ;
      LAYER met1 ;
        RECT 1757.285 1838.960 1757.575 1839.005 ;
        RECT 1757.730 1838.960 1758.050 1839.020 ;
        RECT 1757.285 1838.820 1758.050 1838.960 ;
        RECT 1757.285 1838.775 1757.575 1838.820 ;
        RECT 1757.730 1838.760 1758.050 1838.820 ;
        RECT 1757.285 1803.940 1757.575 1803.985 ;
        RECT 1757.730 1803.940 1758.050 1804.000 ;
        RECT 1757.285 1803.800 1758.050 1803.940 ;
        RECT 1757.285 1803.755 1757.575 1803.800 ;
        RECT 1757.730 1803.740 1758.050 1803.800 ;
      LAYER via ;
        RECT 1757.760 1838.760 1758.020 1839.020 ;
        RECT 1757.760 1803.740 1758.020 1804.000 ;
      LAYER met2 ;
        RECT 1757.750 1857.915 1758.030 1858.285 ;
        RECT 1757.820 1839.050 1757.960 1857.915 ;
        RECT 1757.760 1838.730 1758.020 1839.050 ;
        RECT 1757.760 1803.885 1758.020 1804.030 ;
        RECT 1757.750 1803.515 1758.030 1803.885 ;
        RECT 1765.110 1548.515 1765.390 1548.885 ;
        RECT 1765.180 1538.685 1765.320 1548.515 ;
        RECT 1765.110 1538.315 1765.390 1538.685 ;
        RECT 1758.210 593.795 1758.490 594.165 ;
        RECT 1758.280 573.085 1758.420 593.795 ;
        RECT 1758.210 572.715 1758.490 573.085 ;
        RECT 1758.210 497.235 1758.490 497.605 ;
        RECT 1758.280 476.525 1758.420 497.235 ;
        RECT 1758.210 476.155 1758.490 476.525 ;
        RECT 1758.210 323.155 1758.490 323.525 ;
        RECT 1758.280 235.125 1758.420 323.155 ;
        RECT 1758.210 234.755 1758.490 235.125 ;
        RECT 1020.370 64.755 1020.650 65.125 ;
        RECT 1020.440 7.210 1020.580 64.755 ;
        RECT 1019.520 7.070 1020.580 7.210 ;
        RECT 1019.520 2.400 1019.660 7.070 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
      LAYER via2 ;
        RECT 1757.750 1857.960 1758.030 1858.240 ;
        RECT 1757.750 1803.560 1758.030 1803.840 ;
        RECT 1765.110 1548.560 1765.390 1548.840 ;
        RECT 1765.110 1538.360 1765.390 1538.640 ;
        RECT 1758.210 593.840 1758.490 594.120 ;
        RECT 1758.210 572.760 1758.490 573.040 ;
        RECT 1758.210 497.280 1758.490 497.560 ;
        RECT 1758.210 476.200 1758.490 476.480 ;
        RECT 1758.210 323.200 1758.490 323.480 ;
        RECT 1758.210 234.800 1758.490 235.080 ;
        RECT 1020.370 64.800 1020.650 65.080 ;
      LAYER met3 ;
        RECT 1755.835 1860.375 1759.835 1860.975 ;
        RECT 1757.510 1858.265 1757.810 1860.375 ;
        RECT 1757.510 1857.950 1758.055 1858.265 ;
        RECT 1757.725 1857.935 1758.055 1857.950 ;
        RECT 1756.550 1803.850 1756.930 1803.860 ;
        RECT 1757.725 1803.850 1758.055 1803.865 ;
        RECT 1756.550 1803.550 1758.055 1803.850 ;
        RECT 1756.550 1803.540 1756.930 1803.550 ;
        RECT 1757.725 1803.535 1758.055 1803.550 ;
        RECT 1756.550 1548.850 1756.930 1548.860 ;
        RECT 1765.085 1548.850 1765.415 1548.865 ;
        RECT 1756.550 1548.550 1765.415 1548.850 ;
        RECT 1756.550 1548.540 1756.930 1548.550 ;
        RECT 1765.085 1548.535 1765.415 1548.550 ;
        RECT 1758.390 1538.650 1758.770 1538.660 ;
        RECT 1765.085 1538.650 1765.415 1538.665 ;
        RECT 1758.390 1538.350 1765.415 1538.650 ;
        RECT 1758.390 1538.340 1758.770 1538.350 ;
        RECT 1765.085 1538.335 1765.415 1538.350 ;
        RECT 1756.550 1409.450 1756.930 1409.460 ;
        RECT 1763.910 1409.450 1764.290 1409.460 ;
        RECT 1756.550 1409.150 1764.290 1409.450 ;
        RECT 1756.550 1409.140 1756.930 1409.150 ;
        RECT 1763.910 1409.140 1764.290 1409.150 ;
        RECT 1757.470 1401.970 1757.850 1401.980 ;
        RECT 1763.910 1401.970 1764.290 1401.980 ;
        RECT 1757.470 1401.670 1764.290 1401.970 ;
        RECT 1757.470 1401.660 1757.850 1401.670 ;
        RECT 1763.910 1401.660 1764.290 1401.670 ;
        RECT 1754.710 1149.010 1755.090 1149.020 ;
        RECT 1758.390 1149.010 1758.770 1149.020 ;
        RECT 1754.710 1148.710 1758.770 1149.010 ;
        RECT 1754.710 1148.700 1755.090 1148.710 ;
        RECT 1758.390 1148.700 1758.770 1148.710 ;
        RECT 1754.710 1078.290 1755.090 1078.300 ;
        RECT 1758.390 1078.290 1758.770 1078.300 ;
        RECT 1754.710 1077.990 1758.770 1078.290 ;
        RECT 1754.710 1077.980 1755.090 1077.990 ;
        RECT 1758.390 1077.980 1758.770 1077.990 ;
        RECT 1754.710 1052.450 1755.090 1052.460 ;
        RECT 1758.390 1052.450 1758.770 1052.460 ;
        RECT 1754.710 1052.150 1758.770 1052.450 ;
        RECT 1754.710 1052.140 1755.090 1052.150 ;
        RECT 1758.390 1052.140 1758.770 1052.150 ;
        RECT 1754.710 981.730 1755.090 981.740 ;
        RECT 1758.390 981.730 1758.770 981.740 ;
        RECT 1754.710 981.430 1758.770 981.730 ;
        RECT 1754.710 981.420 1755.090 981.430 ;
        RECT 1758.390 981.420 1758.770 981.430 ;
        RECT 1754.710 955.890 1755.090 955.900 ;
        RECT 1758.390 955.890 1758.770 955.900 ;
        RECT 1754.710 955.590 1758.770 955.890 ;
        RECT 1754.710 955.580 1755.090 955.590 ;
        RECT 1758.390 955.580 1758.770 955.590 ;
        RECT 1753.790 905.570 1754.170 905.580 ;
        RECT 1758.390 905.570 1758.770 905.580 ;
        RECT 1753.790 905.270 1758.770 905.570 ;
        RECT 1753.790 905.260 1754.170 905.270 ;
        RECT 1758.390 905.260 1758.770 905.270 ;
        RECT 1755.630 796.770 1756.010 796.780 ;
        RECT 1758.390 796.770 1758.770 796.780 ;
        RECT 1755.630 796.470 1758.770 796.770 ;
        RECT 1755.630 796.460 1756.010 796.470 ;
        RECT 1758.390 796.460 1758.770 796.470 ;
        RECT 1754.710 690.690 1755.090 690.700 ;
        RECT 1758.390 690.690 1758.770 690.700 ;
        RECT 1754.710 690.390 1758.770 690.690 ;
        RECT 1754.710 690.380 1755.090 690.390 ;
        RECT 1758.390 690.380 1758.770 690.390 ;
        RECT 1754.710 690.010 1755.090 690.020 ;
        RECT 1758.390 690.010 1758.770 690.020 ;
        RECT 1754.710 689.710 1758.770 690.010 ;
        RECT 1754.710 689.700 1755.090 689.710 ;
        RECT 1758.390 689.700 1758.770 689.710 ;
        RECT 1758.185 594.140 1758.515 594.145 ;
        RECT 1758.185 594.130 1758.770 594.140 ;
        RECT 1757.960 593.830 1758.770 594.130 ;
        RECT 1758.185 593.820 1758.770 593.830 ;
        RECT 1758.185 593.815 1758.515 593.820 ;
        RECT 1758.185 573.060 1758.515 573.065 ;
        RECT 1758.185 573.050 1758.770 573.060 ;
        RECT 1758.185 572.750 1758.970 573.050 ;
        RECT 1758.185 572.740 1758.770 572.750 ;
        RECT 1758.185 572.735 1758.515 572.740 ;
        RECT 1758.185 497.580 1758.515 497.585 ;
        RECT 1758.185 497.570 1758.770 497.580 ;
        RECT 1757.960 497.270 1758.770 497.570 ;
        RECT 1758.185 497.260 1758.770 497.270 ;
        RECT 1758.185 497.255 1758.515 497.260 ;
        RECT 1758.185 476.500 1758.515 476.505 ;
        RECT 1758.185 476.490 1758.770 476.500 ;
        RECT 1758.185 476.190 1758.970 476.490 ;
        RECT 1758.185 476.180 1758.770 476.190 ;
        RECT 1758.185 476.175 1758.515 476.180 ;
        RECT 1755.630 403.730 1756.010 403.740 ;
        RECT 1758.390 403.730 1758.770 403.740 ;
        RECT 1755.630 403.430 1758.770 403.730 ;
        RECT 1755.630 403.420 1756.010 403.430 ;
        RECT 1758.390 403.420 1758.770 403.430 ;
        RECT 1756.550 323.860 1756.930 324.180 ;
        RECT 1756.590 323.490 1756.890 323.860 ;
        RECT 1758.185 323.490 1758.515 323.505 ;
        RECT 1756.590 323.190 1758.515 323.490 ;
        RECT 1758.185 323.175 1758.515 323.190 ;
        RECT 1758.185 235.100 1758.515 235.105 ;
        RECT 1758.185 235.090 1758.770 235.100 ;
        RECT 1758.185 234.790 1758.970 235.090 ;
        RECT 1758.185 234.780 1758.770 234.790 ;
        RECT 1758.185 234.775 1758.515 234.780 ;
        RECT 1756.550 207.210 1756.930 207.220 ;
        RECT 1758.390 207.210 1758.770 207.220 ;
        RECT 1756.550 206.910 1758.770 207.210 ;
        RECT 1756.550 206.900 1756.930 206.910 ;
        RECT 1758.390 206.900 1758.770 206.910 ;
        RECT 1020.345 65.090 1020.675 65.105 ;
        RECT 1753.790 65.090 1754.170 65.100 ;
        RECT 1020.345 64.790 1754.170 65.090 ;
        RECT 1020.345 64.775 1020.675 64.790 ;
        RECT 1753.790 64.780 1754.170 64.790 ;
      LAYER via3 ;
        RECT 1756.580 1803.540 1756.900 1803.860 ;
        RECT 1756.580 1548.540 1756.900 1548.860 ;
        RECT 1758.420 1538.340 1758.740 1538.660 ;
        RECT 1756.580 1409.140 1756.900 1409.460 ;
        RECT 1763.940 1409.140 1764.260 1409.460 ;
        RECT 1757.500 1401.660 1757.820 1401.980 ;
        RECT 1763.940 1401.660 1764.260 1401.980 ;
        RECT 1754.740 1148.700 1755.060 1149.020 ;
        RECT 1758.420 1148.700 1758.740 1149.020 ;
        RECT 1754.740 1077.980 1755.060 1078.300 ;
        RECT 1758.420 1077.980 1758.740 1078.300 ;
        RECT 1754.740 1052.140 1755.060 1052.460 ;
        RECT 1758.420 1052.140 1758.740 1052.460 ;
        RECT 1754.740 981.420 1755.060 981.740 ;
        RECT 1758.420 981.420 1758.740 981.740 ;
        RECT 1754.740 955.580 1755.060 955.900 ;
        RECT 1758.420 955.580 1758.740 955.900 ;
        RECT 1753.820 905.260 1754.140 905.580 ;
        RECT 1758.420 905.260 1758.740 905.580 ;
        RECT 1755.660 796.460 1755.980 796.780 ;
        RECT 1758.420 796.460 1758.740 796.780 ;
        RECT 1754.740 690.380 1755.060 690.700 ;
        RECT 1758.420 690.380 1758.740 690.700 ;
        RECT 1754.740 689.700 1755.060 690.020 ;
        RECT 1758.420 689.700 1758.740 690.020 ;
        RECT 1758.420 593.820 1758.740 594.140 ;
        RECT 1758.420 572.740 1758.740 573.060 ;
        RECT 1758.420 497.260 1758.740 497.580 ;
        RECT 1758.420 476.180 1758.740 476.500 ;
        RECT 1755.660 403.420 1755.980 403.740 ;
        RECT 1758.420 403.420 1758.740 403.740 ;
        RECT 1756.580 323.860 1756.900 324.180 ;
        RECT 1758.420 234.780 1758.740 235.100 ;
        RECT 1756.580 206.900 1756.900 207.220 ;
        RECT 1758.420 206.900 1758.740 207.220 ;
        RECT 1753.820 64.780 1754.140 65.100 ;
      LAYER met4 ;
        RECT 1756.575 1803.850 1756.905 1803.865 ;
        RECT 1755.670 1803.550 1756.905 1803.850 ;
        RECT 1755.670 1752.850 1755.970 1803.550 ;
        RECT 1756.575 1803.535 1756.905 1803.550 ;
        RECT 1754.750 1752.550 1755.970 1752.850 ;
        RECT 1754.750 1573.330 1755.050 1752.550 ;
        RECT 1753.830 1573.030 1755.050 1573.330 ;
        RECT 1753.830 1569.250 1754.130 1573.030 ;
        RECT 1753.830 1568.950 1755.050 1569.250 ;
        RECT 1754.750 1548.850 1755.050 1568.950 ;
        RECT 1756.575 1548.850 1756.905 1548.865 ;
        RECT 1754.750 1548.550 1756.905 1548.850 ;
        RECT 1756.575 1548.535 1756.905 1548.550 ;
        RECT 1758.415 1538.650 1758.745 1538.665 ;
        RECT 1755.670 1538.350 1758.745 1538.650 ;
        RECT 1755.670 1521.650 1755.970 1538.350 ;
        RECT 1758.415 1538.335 1758.745 1538.350 ;
        RECT 1754.750 1521.350 1755.970 1521.650 ;
        RECT 1754.750 1409.450 1755.050 1521.350 ;
        RECT 1756.575 1409.450 1756.905 1409.465 ;
        RECT 1754.750 1409.150 1756.905 1409.450 ;
        RECT 1756.575 1409.135 1756.905 1409.150 ;
        RECT 1763.935 1409.135 1764.265 1409.465 ;
        RECT 1763.950 1401.985 1764.250 1409.135 ;
        RECT 1757.495 1401.655 1757.825 1401.985 ;
        RECT 1763.935 1401.655 1764.265 1401.985 ;
        RECT 1757.510 1367.290 1757.810 1401.655 ;
        RECT 1756.590 1366.990 1757.810 1367.290 ;
        RECT 1756.590 1365.250 1756.890 1366.990 ;
        RECT 1756.360 1364.950 1756.890 1365.250 ;
        RECT 1756.360 1364.570 1756.660 1364.950 ;
        RECT 1754.750 1364.270 1756.660 1364.570 ;
        RECT 1754.750 1290.450 1755.050 1364.270 ;
        RECT 1753.830 1290.150 1755.050 1290.450 ;
        RECT 1753.830 1249.650 1754.130 1290.150 ;
        RECT 1753.830 1249.350 1755.050 1249.650 ;
        RECT 1754.750 1242.850 1755.050 1249.350 ;
        RECT 1754.750 1242.550 1755.970 1242.850 ;
        RECT 1755.670 1178.250 1755.970 1242.550 ;
        RECT 1754.750 1177.950 1755.970 1178.250 ;
        RECT 1754.750 1149.025 1755.050 1177.950 ;
        RECT 1754.735 1148.695 1755.065 1149.025 ;
        RECT 1758.415 1148.695 1758.745 1149.025 ;
        RECT 1758.430 1078.305 1758.730 1148.695 ;
        RECT 1754.735 1077.975 1755.065 1078.305 ;
        RECT 1758.415 1077.975 1758.745 1078.305 ;
        RECT 1754.750 1052.465 1755.050 1077.975 ;
        RECT 1754.735 1052.135 1755.065 1052.465 ;
        RECT 1758.415 1052.135 1758.745 1052.465 ;
        RECT 1758.430 981.745 1758.730 1052.135 ;
        RECT 1754.735 981.415 1755.065 981.745 ;
        RECT 1758.415 981.415 1758.745 981.745 ;
        RECT 1754.750 955.905 1755.050 981.415 ;
        RECT 1754.735 955.575 1755.065 955.905 ;
        RECT 1758.415 955.575 1758.745 955.905 ;
        RECT 1758.430 905.585 1758.730 955.575 ;
        RECT 1753.815 905.255 1754.145 905.585 ;
        RECT 1758.415 905.255 1758.745 905.585 ;
        RECT 1753.830 865.450 1754.130 905.255 ;
        RECT 1753.830 865.150 1755.970 865.450 ;
        RECT 1755.670 796.785 1755.970 865.150 ;
        RECT 1755.655 796.455 1755.985 796.785 ;
        RECT 1758.415 796.455 1758.745 796.785 ;
        RECT 1758.430 690.705 1758.730 796.455 ;
        RECT 1754.735 690.375 1755.065 690.705 ;
        RECT 1758.415 690.375 1758.745 690.705 ;
        RECT 1754.750 690.025 1755.050 690.375 ;
        RECT 1754.735 689.695 1755.065 690.025 ;
        RECT 1758.415 689.695 1758.745 690.025 ;
        RECT 1758.430 594.145 1758.730 689.695 ;
        RECT 1758.415 593.815 1758.745 594.145 ;
        RECT 1758.415 572.735 1758.745 573.065 ;
        RECT 1758.430 497.585 1758.730 572.735 ;
        RECT 1758.415 497.255 1758.745 497.585 ;
        RECT 1758.415 476.175 1758.745 476.505 ;
        RECT 1758.430 403.745 1758.730 476.175 ;
        RECT 1755.655 403.415 1755.985 403.745 ;
        RECT 1758.415 403.415 1758.745 403.745 ;
        RECT 1755.670 324.850 1755.970 403.415 ;
        RECT 1755.670 324.550 1756.890 324.850 ;
        RECT 1756.590 324.185 1756.890 324.550 ;
        RECT 1756.575 323.855 1756.905 324.185 ;
        RECT 1758.415 234.775 1758.745 235.105 ;
        RECT 1758.430 207.225 1758.730 234.775 ;
        RECT 1756.575 206.895 1756.905 207.225 ;
        RECT 1758.415 206.895 1758.745 207.225 ;
        RECT 1756.590 141.250 1756.890 206.895 ;
        RECT 1753.830 140.950 1756.890 141.250 ;
        RECT 1753.830 65.105 1754.130 140.950 ;
        RECT 1753.815 64.775 1754.145 65.105 ;
    END
  END la_oen[21]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1055.310 1293.600 1055.630 1293.660 ;
        RECT 1765.090 1293.600 1765.410 1293.660 ;
        RECT 1055.310 1293.460 1765.410 1293.600 ;
        RECT 1055.310 1293.400 1055.630 1293.460 ;
        RECT 1765.090 1293.400 1765.410 1293.460 ;
      LAYER via ;
        RECT 1055.340 1293.400 1055.600 1293.660 ;
        RECT 1765.120 1293.400 1765.380 1293.660 ;
      LAYER met2 ;
        RECT 1765.110 1475.755 1765.390 1476.125 ;
        RECT 1765.180 1293.690 1765.320 1475.755 ;
        RECT 1055.340 1293.370 1055.600 1293.690 ;
        RECT 1765.120 1293.370 1765.380 1293.690 ;
        RECT 1055.400 2.400 1055.540 1293.370 ;
        RECT 1055.190 -4.800 1055.750 2.400 ;
      LAYER via2 ;
        RECT 1765.110 1475.800 1765.390 1476.080 ;
      LAYER met3 ;
        RECT 1755.835 1476.090 1759.835 1476.095 ;
        RECT 1765.085 1476.090 1765.415 1476.105 ;
        RECT 1755.835 1475.790 1765.415 1476.090 ;
        RECT 1755.835 1475.495 1759.835 1475.790 ;
        RECT 1765.085 1475.775 1765.415 1475.790 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1070.105 1326.425 1070.275 1330.335 ;
      LAYER mcon ;
        RECT 1070.105 1330.165 1070.275 1330.335 ;
      LAYER met1 ;
        RECT 715.830 1330.320 716.150 1330.380 ;
        RECT 1070.045 1330.320 1070.335 1330.365 ;
        RECT 715.830 1330.180 1070.335 1330.320 ;
        RECT 715.830 1330.120 716.150 1330.180 ;
        RECT 1070.045 1330.135 1070.335 1330.180 ;
        RECT 1070.030 1326.580 1070.350 1326.640 ;
        RECT 1069.835 1326.440 1070.350 1326.580 ;
        RECT 1070.030 1326.380 1070.350 1326.440 ;
        RECT 1070.030 2.960 1070.350 3.020 ;
        RECT 1073.250 2.960 1073.570 3.020 ;
        RECT 1070.030 2.820 1073.570 2.960 ;
        RECT 1070.030 2.760 1070.350 2.820 ;
        RECT 1073.250 2.760 1073.570 2.820 ;
      LAYER via ;
        RECT 715.860 1330.120 716.120 1330.380 ;
        RECT 1070.060 1326.380 1070.320 1326.640 ;
        RECT 1070.060 2.760 1070.320 3.020 ;
        RECT 1073.280 2.760 1073.540 3.020 ;
      LAYER met2 ;
        RECT 715.850 2128.555 716.130 2128.925 ;
        RECT 715.920 1330.410 716.060 2128.555 ;
        RECT 715.860 1330.090 716.120 1330.410 ;
        RECT 1070.060 1326.350 1070.320 1326.670 ;
        RECT 1070.120 3.050 1070.260 1326.350 ;
        RECT 1070.060 2.730 1070.320 3.050 ;
        RECT 1073.280 2.730 1073.540 3.050 ;
        RECT 1073.340 2.400 1073.480 2.730 ;
        RECT 1073.130 -4.800 1073.690 2.400 ;
      LAYER via2 ;
        RECT 715.850 2128.600 716.130 2128.880 ;
      LAYER met3 ;
        RECT 715.810 2131.015 719.810 2131.615 ;
        RECT 716.070 2128.905 716.370 2131.015 ;
        RECT 715.825 2128.590 716.370 2128.905 ;
        RECT 715.825 2128.575 716.155 2128.590 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1766.470 1221.180 1766.790 1221.240 ;
        RECT 1768.770 1221.180 1769.090 1221.240 ;
        RECT 1766.470 1221.040 1769.090 1221.180 ;
        RECT 1766.470 1220.980 1766.790 1221.040 ;
        RECT 1768.770 1220.980 1769.090 1221.040 ;
        RECT 1766.470 1173.240 1766.790 1173.300 ;
        RECT 1768.770 1173.240 1769.090 1173.300 ;
        RECT 1766.470 1173.100 1769.090 1173.240 ;
        RECT 1766.470 1173.040 1766.790 1173.100 ;
        RECT 1768.770 1173.040 1769.090 1173.100 ;
        RECT 1766.470 1124.620 1766.790 1124.680 ;
        RECT 1768.770 1124.620 1769.090 1124.680 ;
        RECT 1766.470 1124.480 1769.090 1124.620 ;
        RECT 1766.470 1124.420 1766.790 1124.480 ;
        RECT 1768.770 1124.420 1769.090 1124.480 ;
        RECT 1766.470 1076.680 1766.790 1076.740 ;
        RECT 1768.770 1076.680 1769.090 1076.740 ;
        RECT 1766.470 1076.540 1769.090 1076.680 ;
        RECT 1766.470 1076.480 1766.790 1076.540 ;
        RECT 1768.770 1076.480 1769.090 1076.540 ;
        RECT 1766.470 1027.720 1766.790 1027.780 ;
        RECT 1768.770 1027.720 1769.090 1027.780 ;
        RECT 1766.470 1027.580 1769.090 1027.720 ;
        RECT 1766.470 1027.520 1766.790 1027.580 ;
        RECT 1768.770 1027.520 1769.090 1027.580 ;
        RECT 1766.470 980.120 1766.790 980.180 ;
        RECT 1768.770 980.120 1769.090 980.180 ;
        RECT 1766.470 979.980 1769.090 980.120 ;
        RECT 1766.470 979.920 1766.790 979.980 ;
        RECT 1768.770 979.920 1769.090 979.980 ;
        RECT 1766.470 931.500 1766.790 931.560 ;
        RECT 1768.770 931.500 1769.090 931.560 ;
        RECT 1766.470 931.360 1769.090 931.500 ;
        RECT 1766.470 931.300 1766.790 931.360 ;
        RECT 1768.770 931.300 1769.090 931.360 ;
        RECT 1766.470 883.560 1766.790 883.620 ;
        RECT 1768.770 883.560 1769.090 883.620 ;
        RECT 1766.470 883.420 1769.090 883.560 ;
        RECT 1766.470 883.360 1766.790 883.420 ;
        RECT 1768.770 883.360 1769.090 883.420 ;
        RECT 1766.470 834.940 1766.790 835.000 ;
        RECT 1768.770 834.940 1769.090 835.000 ;
        RECT 1766.470 834.800 1769.090 834.940 ;
        RECT 1766.470 834.740 1766.790 834.800 ;
        RECT 1768.770 834.740 1769.090 834.800 ;
        RECT 1766.470 787.000 1766.790 787.060 ;
        RECT 1768.770 787.000 1769.090 787.060 ;
        RECT 1766.470 786.860 1769.090 787.000 ;
        RECT 1766.470 786.800 1766.790 786.860 ;
        RECT 1768.770 786.800 1769.090 786.860 ;
        RECT 1766.470 738.040 1766.790 738.100 ;
        RECT 1768.770 738.040 1769.090 738.100 ;
        RECT 1766.470 737.900 1769.090 738.040 ;
        RECT 1766.470 737.840 1766.790 737.900 ;
        RECT 1768.770 737.840 1769.090 737.900 ;
        RECT 1766.470 690.100 1766.790 690.160 ;
        RECT 1768.770 690.100 1769.090 690.160 ;
        RECT 1766.470 689.960 1769.090 690.100 ;
        RECT 1766.470 689.900 1766.790 689.960 ;
        RECT 1768.770 689.900 1769.090 689.960 ;
        RECT 1766.470 641.480 1766.790 641.540 ;
        RECT 1768.770 641.480 1769.090 641.540 ;
        RECT 1766.470 641.340 1769.090 641.480 ;
        RECT 1766.470 641.280 1766.790 641.340 ;
        RECT 1768.770 641.280 1769.090 641.340 ;
        RECT 1766.470 593.540 1766.790 593.600 ;
        RECT 1768.770 593.540 1769.090 593.600 ;
        RECT 1766.470 593.400 1769.090 593.540 ;
        RECT 1766.470 593.340 1766.790 593.400 ;
        RECT 1768.770 593.340 1769.090 593.400 ;
        RECT 1766.470 544.920 1766.790 544.980 ;
        RECT 1768.770 544.920 1769.090 544.980 ;
        RECT 1766.470 544.780 1769.090 544.920 ;
        RECT 1766.470 544.720 1766.790 544.780 ;
        RECT 1768.770 544.720 1769.090 544.780 ;
        RECT 1766.470 496.980 1766.790 497.040 ;
        RECT 1768.770 496.980 1769.090 497.040 ;
        RECT 1766.470 496.840 1769.090 496.980 ;
        RECT 1766.470 496.780 1766.790 496.840 ;
        RECT 1768.770 496.780 1769.090 496.840 ;
        RECT 1766.470 351.800 1766.790 351.860 ;
        RECT 1768.770 351.800 1769.090 351.860 ;
        RECT 1766.470 351.660 1769.090 351.800 ;
        RECT 1766.470 351.600 1766.790 351.660 ;
        RECT 1768.770 351.600 1769.090 351.660 ;
        RECT 1766.470 303.860 1766.790 303.920 ;
        RECT 1768.770 303.860 1769.090 303.920 ;
        RECT 1766.470 303.720 1769.090 303.860 ;
        RECT 1766.470 303.660 1766.790 303.720 ;
        RECT 1768.770 303.660 1769.090 303.720 ;
        RECT 1766.470 255.240 1766.790 255.300 ;
        RECT 1768.770 255.240 1769.090 255.300 ;
        RECT 1766.470 255.100 1769.090 255.240 ;
        RECT 1766.470 255.040 1766.790 255.100 ;
        RECT 1768.770 255.040 1769.090 255.100 ;
        RECT 1766.470 207.300 1766.790 207.360 ;
        RECT 1768.770 207.300 1769.090 207.360 ;
        RECT 1766.470 207.160 1769.090 207.300 ;
        RECT 1766.470 207.100 1766.790 207.160 ;
        RECT 1768.770 207.100 1769.090 207.160 ;
        RECT 1096.710 68.240 1097.030 68.300 ;
        RECT 1766.470 68.240 1766.790 68.300 ;
        RECT 1096.710 68.100 1766.790 68.240 ;
        RECT 1096.710 68.040 1097.030 68.100 ;
        RECT 1766.470 68.040 1766.790 68.100 ;
        RECT 1090.730 20.640 1091.050 20.700 ;
        RECT 1096.710 20.640 1097.030 20.700 ;
        RECT 1090.730 20.500 1097.030 20.640 ;
        RECT 1090.730 20.440 1091.050 20.500 ;
        RECT 1096.710 20.440 1097.030 20.500 ;
      LAYER via ;
        RECT 1766.500 1220.980 1766.760 1221.240 ;
        RECT 1768.800 1220.980 1769.060 1221.240 ;
        RECT 1766.500 1173.040 1766.760 1173.300 ;
        RECT 1768.800 1173.040 1769.060 1173.300 ;
        RECT 1766.500 1124.420 1766.760 1124.680 ;
        RECT 1768.800 1124.420 1769.060 1124.680 ;
        RECT 1766.500 1076.480 1766.760 1076.740 ;
        RECT 1768.800 1076.480 1769.060 1076.740 ;
        RECT 1766.500 1027.520 1766.760 1027.780 ;
        RECT 1768.800 1027.520 1769.060 1027.780 ;
        RECT 1766.500 979.920 1766.760 980.180 ;
        RECT 1768.800 979.920 1769.060 980.180 ;
        RECT 1766.500 931.300 1766.760 931.560 ;
        RECT 1768.800 931.300 1769.060 931.560 ;
        RECT 1766.500 883.360 1766.760 883.620 ;
        RECT 1768.800 883.360 1769.060 883.620 ;
        RECT 1766.500 834.740 1766.760 835.000 ;
        RECT 1768.800 834.740 1769.060 835.000 ;
        RECT 1766.500 786.800 1766.760 787.060 ;
        RECT 1768.800 786.800 1769.060 787.060 ;
        RECT 1766.500 737.840 1766.760 738.100 ;
        RECT 1768.800 737.840 1769.060 738.100 ;
        RECT 1766.500 689.900 1766.760 690.160 ;
        RECT 1768.800 689.900 1769.060 690.160 ;
        RECT 1766.500 641.280 1766.760 641.540 ;
        RECT 1768.800 641.280 1769.060 641.540 ;
        RECT 1766.500 593.340 1766.760 593.600 ;
        RECT 1768.800 593.340 1769.060 593.600 ;
        RECT 1766.500 544.720 1766.760 544.980 ;
        RECT 1768.800 544.720 1769.060 544.980 ;
        RECT 1766.500 496.780 1766.760 497.040 ;
        RECT 1768.800 496.780 1769.060 497.040 ;
        RECT 1766.500 351.600 1766.760 351.860 ;
        RECT 1768.800 351.600 1769.060 351.860 ;
        RECT 1766.500 303.660 1766.760 303.920 ;
        RECT 1768.800 303.660 1769.060 303.920 ;
        RECT 1766.500 255.040 1766.760 255.300 ;
        RECT 1768.800 255.040 1769.060 255.300 ;
        RECT 1766.500 207.100 1766.760 207.360 ;
        RECT 1768.800 207.100 1769.060 207.360 ;
        RECT 1096.740 68.040 1097.000 68.300 ;
        RECT 1766.500 68.040 1766.760 68.300 ;
        RECT 1090.760 20.440 1091.020 20.700 ;
        RECT 1096.740 20.440 1097.000 20.700 ;
      LAYER met2 ;
        RECT 1766.490 2049.675 1766.770 2050.045 ;
        RECT 1766.560 1221.270 1766.700 2049.675 ;
        RECT 1766.500 1220.950 1766.760 1221.270 ;
        RECT 1768.800 1220.950 1769.060 1221.270 ;
        RECT 1768.860 1173.330 1769.000 1220.950 ;
        RECT 1766.500 1173.010 1766.760 1173.330 ;
        RECT 1768.800 1173.010 1769.060 1173.330 ;
        RECT 1766.560 1124.710 1766.700 1173.010 ;
        RECT 1766.500 1124.390 1766.760 1124.710 ;
        RECT 1768.800 1124.390 1769.060 1124.710 ;
        RECT 1768.860 1076.770 1769.000 1124.390 ;
        RECT 1766.500 1076.450 1766.760 1076.770 ;
        RECT 1768.800 1076.450 1769.060 1076.770 ;
        RECT 1766.560 1027.810 1766.700 1076.450 ;
        RECT 1766.500 1027.490 1766.760 1027.810 ;
        RECT 1768.800 1027.490 1769.060 1027.810 ;
        RECT 1768.860 980.210 1769.000 1027.490 ;
        RECT 1766.500 979.890 1766.760 980.210 ;
        RECT 1768.800 979.890 1769.060 980.210 ;
        RECT 1766.560 931.590 1766.700 979.890 ;
        RECT 1766.500 931.270 1766.760 931.590 ;
        RECT 1768.800 931.270 1769.060 931.590 ;
        RECT 1768.860 883.650 1769.000 931.270 ;
        RECT 1766.500 883.330 1766.760 883.650 ;
        RECT 1768.800 883.330 1769.060 883.650 ;
        RECT 1766.560 835.030 1766.700 883.330 ;
        RECT 1766.500 834.710 1766.760 835.030 ;
        RECT 1768.800 834.710 1769.060 835.030 ;
        RECT 1768.860 787.090 1769.000 834.710 ;
        RECT 1766.500 786.770 1766.760 787.090 ;
        RECT 1768.800 786.770 1769.060 787.090 ;
        RECT 1766.560 738.130 1766.700 786.770 ;
        RECT 1766.500 737.810 1766.760 738.130 ;
        RECT 1768.800 737.810 1769.060 738.130 ;
        RECT 1768.860 690.190 1769.000 737.810 ;
        RECT 1766.500 689.870 1766.760 690.190 ;
        RECT 1768.800 689.870 1769.060 690.190 ;
        RECT 1766.560 641.570 1766.700 689.870 ;
        RECT 1766.500 641.250 1766.760 641.570 ;
        RECT 1768.800 641.250 1769.060 641.570 ;
        RECT 1768.860 593.630 1769.000 641.250 ;
        RECT 1766.500 593.310 1766.760 593.630 ;
        RECT 1768.800 593.310 1769.060 593.630 ;
        RECT 1766.560 545.010 1766.700 593.310 ;
        RECT 1766.500 544.690 1766.760 545.010 ;
        RECT 1768.800 544.690 1769.060 545.010 ;
        RECT 1768.860 497.070 1769.000 544.690 ;
        RECT 1766.500 496.750 1766.760 497.070 ;
        RECT 1768.800 496.750 1769.060 497.070 ;
        RECT 1766.560 351.890 1766.700 496.750 ;
        RECT 1766.500 351.570 1766.760 351.890 ;
        RECT 1768.800 351.570 1769.060 351.890 ;
        RECT 1768.860 303.950 1769.000 351.570 ;
        RECT 1766.500 303.630 1766.760 303.950 ;
        RECT 1768.800 303.630 1769.060 303.950 ;
        RECT 1766.560 255.330 1766.700 303.630 ;
        RECT 1766.500 255.010 1766.760 255.330 ;
        RECT 1768.800 255.010 1769.060 255.330 ;
        RECT 1768.860 207.390 1769.000 255.010 ;
        RECT 1766.500 207.070 1766.760 207.390 ;
        RECT 1768.800 207.070 1769.060 207.390 ;
        RECT 1766.560 68.330 1766.700 207.070 ;
        RECT 1096.740 68.010 1097.000 68.330 ;
        RECT 1766.500 68.010 1766.760 68.330 ;
        RECT 1096.800 20.730 1096.940 68.010 ;
        RECT 1090.760 20.410 1091.020 20.730 ;
        RECT 1096.740 20.410 1097.000 20.730 ;
        RECT 1090.820 2.400 1090.960 20.410 ;
        RECT 1090.610 -4.800 1091.170 2.400 ;
      LAYER via2 ;
        RECT 1766.490 2049.720 1766.770 2050.000 ;
      LAYER met3 ;
        RECT 1755.835 2050.010 1759.835 2050.015 ;
        RECT 1766.465 2050.010 1766.795 2050.025 ;
        RECT 1755.835 2049.710 1766.795 2050.010 ;
        RECT 1755.835 2049.415 1759.835 2049.710 ;
        RECT 1766.465 2049.695 1766.795 2049.710 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1109.205 1145.545 1109.375 1193.655 ;
        RECT 1110.125 1013.965 1110.295 1055.615 ;
        RECT 1110.585 524.365 1110.755 554.455 ;
        RECT 1110.585 331.245 1110.755 386.155 ;
        RECT 1110.585 48.365 1110.755 113.815 ;
      LAYER mcon ;
        RECT 1109.205 1193.485 1109.375 1193.655 ;
        RECT 1110.125 1055.445 1110.295 1055.615 ;
        RECT 1110.585 554.285 1110.755 554.455 ;
        RECT 1110.585 385.985 1110.755 386.155 ;
        RECT 1110.585 113.645 1110.755 113.815 ;
      LAYER met1 ;
        RECT 1110.510 1313.320 1110.830 1313.380 ;
        RECT 1157.430 1313.320 1157.750 1313.380 ;
        RECT 1110.510 1313.180 1157.750 1313.320 ;
        RECT 1110.510 1313.120 1110.830 1313.180 ;
        RECT 1157.430 1313.120 1157.750 1313.180 ;
        RECT 1109.145 1193.640 1109.435 1193.685 ;
        RECT 1110.050 1193.640 1110.370 1193.700 ;
        RECT 1109.145 1193.500 1110.370 1193.640 ;
        RECT 1109.145 1193.455 1109.435 1193.500 ;
        RECT 1110.050 1193.440 1110.370 1193.500 ;
        RECT 1109.130 1145.700 1109.450 1145.760 ;
        RECT 1108.935 1145.560 1109.450 1145.700 ;
        RECT 1109.130 1145.500 1109.450 1145.560 ;
        RECT 1109.130 1104.220 1109.450 1104.280 ;
        RECT 1110.510 1104.220 1110.830 1104.280 ;
        RECT 1109.130 1104.080 1110.830 1104.220 ;
        RECT 1109.130 1104.020 1109.450 1104.080 ;
        RECT 1110.510 1104.020 1110.830 1104.080 ;
        RECT 1110.050 1055.600 1110.370 1055.660 ;
        RECT 1109.855 1055.460 1110.370 1055.600 ;
        RECT 1110.050 1055.400 1110.370 1055.460 ;
        RECT 1110.050 1014.120 1110.370 1014.180 ;
        RECT 1109.855 1013.980 1110.370 1014.120 ;
        RECT 1110.050 1013.920 1110.370 1013.980 ;
        RECT 1110.510 554.440 1110.830 554.500 ;
        RECT 1110.315 554.300 1110.830 554.440 ;
        RECT 1110.510 554.240 1110.830 554.300 ;
        RECT 1110.510 524.520 1110.830 524.580 ;
        RECT 1110.315 524.380 1110.830 524.520 ;
        RECT 1110.510 524.320 1110.830 524.380 ;
        RECT 1110.510 386.140 1110.830 386.200 ;
        RECT 1110.315 386.000 1110.830 386.140 ;
        RECT 1110.510 385.940 1110.830 386.000 ;
        RECT 1110.510 331.400 1110.830 331.460 ;
        RECT 1110.315 331.260 1110.830 331.400 ;
        RECT 1110.510 331.200 1110.830 331.260 ;
        RECT 1110.510 113.800 1110.830 113.860 ;
        RECT 1110.315 113.660 1110.830 113.800 ;
        RECT 1110.510 113.600 1110.830 113.660 ;
        RECT 1108.670 48.520 1108.990 48.580 ;
        RECT 1110.525 48.520 1110.815 48.565 ;
        RECT 1108.670 48.380 1110.815 48.520 ;
        RECT 1108.670 48.320 1108.990 48.380 ;
        RECT 1110.525 48.335 1110.815 48.380 ;
      LAYER via ;
        RECT 1110.540 1313.120 1110.800 1313.380 ;
        RECT 1157.460 1313.120 1157.720 1313.380 ;
        RECT 1110.080 1193.440 1110.340 1193.700 ;
        RECT 1109.160 1145.500 1109.420 1145.760 ;
        RECT 1109.160 1104.020 1109.420 1104.280 ;
        RECT 1110.540 1104.020 1110.800 1104.280 ;
        RECT 1110.080 1055.400 1110.340 1055.660 ;
        RECT 1110.080 1013.920 1110.340 1014.180 ;
        RECT 1110.540 554.240 1110.800 554.500 ;
        RECT 1110.540 524.320 1110.800 524.580 ;
        RECT 1110.540 385.940 1110.800 386.200 ;
        RECT 1110.540 331.200 1110.800 331.460 ;
        RECT 1110.540 113.600 1110.800 113.860 ;
        RECT 1108.700 48.320 1108.960 48.580 ;
      LAYER met2 ;
        RECT 1157.500 1323.135 1157.780 1327.135 ;
        RECT 1157.520 1313.410 1157.660 1323.135 ;
        RECT 1110.540 1313.090 1110.800 1313.410 ;
        RECT 1157.460 1313.090 1157.720 1313.410 ;
        RECT 1110.600 1200.610 1110.740 1313.090 ;
        RECT 1110.140 1200.470 1110.740 1200.610 ;
        RECT 1110.140 1193.730 1110.280 1200.470 ;
        RECT 1110.080 1193.410 1110.340 1193.730 ;
        RECT 1109.160 1145.470 1109.420 1145.790 ;
        RECT 1109.220 1104.310 1109.360 1145.470 ;
        RECT 1109.160 1103.990 1109.420 1104.310 ;
        RECT 1110.540 1103.990 1110.800 1104.310 ;
        RECT 1110.600 1080.250 1110.740 1103.990 ;
        RECT 1110.140 1080.110 1110.740 1080.250 ;
        RECT 1110.140 1055.690 1110.280 1080.110 ;
        RECT 1110.080 1055.370 1110.340 1055.690 ;
        RECT 1110.080 1013.890 1110.340 1014.210 ;
        RECT 1110.140 1007.490 1110.280 1013.890 ;
        RECT 1110.140 1007.350 1110.740 1007.490 ;
        RECT 1110.600 554.530 1110.740 1007.350 ;
        RECT 1110.540 554.210 1110.800 554.530 ;
        RECT 1110.540 524.290 1110.800 524.610 ;
        RECT 1110.600 386.230 1110.740 524.290 ;
        RECT 1110.540 385.910 1110.800 386.230 ;
        RECT 1110.540 331.170 1110.800 331.490 ;
        RECT 1110.600 241.640 1110.740 331.170 ;
        RECT 1110.140 241.500 1110.740 241.640 ;
        RECT 1110.140 241.130 1110.280 241.500 ;
        RECT 1110.140 240.990 1110.740 241.130 ;
        RECT 1110.600 113.890 1110.740 240.990 ;
        RECT 1110.540 113.570 1110.800 113.890 ;
        RECT 1108.700 48.290 1108.960 48.610 ;
        RECT 1108.760 2.400 1108.900 48.290 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1007.470 1315.020 1007.790 1315.080 ;
        RECT 1124.770 1315.020 1125.090 1315.080 ;
        RECT 1007.470 1314.880 1125.090 1315.020 ;
        RECT 1007.470 1314.820 1007.790 1314.880 ;
        RECT 1124.770 1314.820 1125.090 1314.880 ;
      LAYER via ;
        RECT 1007.500 1314.820 1007.760 1315.080 ;
        RECT 1124.800 1314.820 1125.060 1315.080 ;
      LAYER met2 ;
        RECT 1007.540 1323.135 1007.820 1327.135 ;
        RECT 1007.560 1315.110 1007.700 1323.135 ;
        RECT 1007.500 1314.790 1007.760 1315.110 ;
        RECT 1124.800 1314.790 1125.060 1315.110 ;
        RECT 1124.860 38.490 1125.000 1314.790 ;
        RECT 1124.860 38.350 1126.840 38.490 ;
        RECT 1126.700 2.400 1126.840 38.350 ;
        RECT 1126.490 -4.800 1127.050 2.400 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1144.625 2.805 1144.795 48.195 ;
      LAYER mcon ;
        RECT 1144.625 48.025 1144.795 48.195 ;
      LAYER met1 ;
        RECT 1749.910 1311.280 1750.230 1311.340 ;
        RECT 1753.590 1311.280 1753.910 1311.340 ;
        RECT 1749.910 1311.140 1753.910 1311.280 ;
        RECT 1749.910 1311.080 1750.230 1311.140 ;
        RECT 1753.590 1311.080 1753.910 1311.140 ;
        RECT 1144.090 87.280 1144.410 87.340 ;
        RECT 1749.910 87.280 1750.230 87.340 ;
        RECT 1144.090 87.140 1750.230 87.280 ;
        RECT 1144.090 87.080 1144.410 87.140 ;
        RECT 1749.910 87.080 1750.230 87.140 ;
        RECT 1144.090 48.180 1144.410 48.240 ;
        RECT 1144.565 48.180 1144.855 48.225 ;
        RECT 1144.090 48.040 1144.855 48.180 ;
        RECT 1144.090 47.980 1144.410 48.040 ;
        RECT 1144.565 47.995 1144.855 48.040 ;
        RECT 1144.550 2.960 1144.870 3.020 ;
        RECT 1144.355 2.820 1144.870 2.960 ;
        RECT 1144.550 2.760 1144.870 2.820 ;
      LAYER via ;
        RECT 1749.940 1311.080 1750.200 1311.340 ;
        RECT 1753.620 1311.080 1753.880 1311.340 ;
        RECT 1144.120 87.080 1144.380 87.340 ;
        RECT 1749.940 87.080 1750.200 87.340 ;
        RECT 1144.120 47.980 1144.380 48.240 ;
        RECT 1144.580 2.760 1144.840 3.020 ;
      LAYER met2 ;
        RECT 1753.660 1323.135 1753.940 1327.135 ;
        RECT 1753.680 1311.370 1753.820 1323.135 ;
        RECT 1749.940 1311.050 1750.200 1311.370 ;
        RECT 1753.620 1311.050 1753.880 1311.370 ;
        RECT 1750.000 87.370 1750.140 1311.050 ;
        RECT 1144.120 87.050 1144.380 87.370 ;
        RECT 1749.940 87.050 1750.200 87.370 ;
        RECT 1144.180 48.270 1144.320 87.050 ;
        RECT 1144.120 47.950 1144.380 48.270 ;
        RECT 1144.580 2.730 1144.840 3.050 ;
        RECT 1144.640 2.400 1144.780 2.730 ;
        RECT 1144.430 -4.800 1144.990 2.400 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1165.710 1312.640 1166.030 1312.700 ;
        RECT 1165.710 1312.500 1197.680 1312.640 ;
        RECT 1165.710 1312.440 1166.030 1312.500 ;
        RECT 1197.540 1312.300 1197.680 1312.500 ;
        RECT 1250.350 1312.300 1250.670 1312.360 ;
        RECT 1197.540 1312.160 1250.670 1312.300 ;
        RECT 1250.350 1312.100 1250.670 1312.160 ;
        RECT 1162.490 20.640 1162.810 20.700 ;
        RECT 1165.710 20.640 1166.030 20.700 ;
        RECT 1162.490 20.500 1166.030 20.640 ;
        RECT 1162.490 20.440 1162.810 20.500 ;
        RECT 1165.710 20.440 1166.030 20.500 ;
      LAYER via ;
        RECT 1165.740 1312.440 1166.000 1312.700 ;
        RECT 1250.380 1312.100 1250.640 1312.360 ;
        RECT 1162.520 20.440 1162.780 20.700 ;
        RECT 1165.740 20.440 1166.000 20.700 ;
      LAYER met2 ;
        RECT 1250.420 1323.135 1250.700 1327.135 ;
        RECT 1165.740 1312.410 1166.000 1312.730 ;
        RECT 1165.800 20.730 1165.940 1312.410 ;
        RECT 1250.440 1312.390 1250.580 1323.135 ;
        RECT 1250.380 1312.070 1250.640 1312.390 ;
        RECT 1162.520 20.410 1162.780 20.730 ;
        RECT 1165.740 20.410 1166.000 20.730 ;
        RECT 1162.580 2.400 1162.720 20.410 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 681.330 1300.740 681.650 1300.800 ;
        RECT 1765.550 1300.740 1765.870 1300.800 ;
        RECT 681.330 1300.600 1765.870 1300.740 ;
        RECT 681.330 1300.540 681.650 1300.600 ;
        RECT 1765.550 1300.540 1765.870 1300.600 ;
        RECT 680.410 2.960 680.730 3.020 ;
        RECT 681.330 2.960 681.650 3.020 ;
        RECT 680.410 2.820 681.650 2.960 ;
        RECT 680.410 2.760 680.730 2.820 ;
        RECT 681.330 2.760 681.650 2.820 ;
      LAYER via ;
        RECT 681.360 1300.540 681.620 1300.800 ;
        RECT 1765.580 1300.540 1765.840 1300.800 ;
        RECT 680.440 2.760 680.700 3.020 ;
        RECT 681.360 2.760 681.620 3.020 ;
      LAYER met2 ;
        RECT 1765.570 1415.915 1765.850 1416.285 ;
        RECT 1765.640 1300.830 1765.780 1415.915 ;
        RECT 681.360 1300.510 681.620 1300.830 ;
        RECT 1765.580 1300.510 1765.840 1300.830 ;
        RECT 681.420 3.050 681.560 1300.510 ;
        RECT 680.440 2.730 680.700 3.050 ;
        RECT 681.360 2.730 681.620 3.050 ;
        RECT 680.500 2.400 680.640 2.730 ;
        RECT 680.290 -4.800 680.850 2.400 ;
      LAYER via2 ;
        RECT 1765.570 1415.960 1765.850 1416.240 ;
      LAYER met3 ;
        RECT 1755.835 1416.250 1759.835 1416.255 ;
        RECT 1765.545 1416.250 1765.875 1416.265 ;
        RECT 1755.835 1415.950 1765.875 1416.250 ;
        RECT 1755.835 1415.655 1759.835 1415.950 ;
        RECT 1765.545 1415.935 1765.875 1415.950 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1186.410 1313.320 1186.730 1313.380 ;
        RECT 1255.870 1313.320 1256.190 1313.380 ;
        RECT 1186.410 1313.180 1256.190 1313.320 ;
        RECT 1186.410 1313.120 1186.730 1313.180 ;
        RECT 1255.870 1313.120 1256.190 1313.180 ;
        RECT 1179.970 16.220 1180.290 16.280 ;
        RECT 1186.410 16.220 1186.730 16.280 ;
        RECT 1179.970 16.080 1186.730 16.220 ;
        RECT 1179.970 16.020 1180.290 16.080 ;
        RECT 1186.410 16.020 1186.730 16.080 ;
      LAYER via ;
        RECT 1186.440 1313.120 1186.700 1313.380 ;
        RECT 1255.900 1313.120 1256.160 1313.380 ;
        RECT 1180.000 16.020 1180.260 16.280 ;
        RECT 1186.440 16.020 1186.700 16.280 ;
      LAYER met2 ;
        RECT 1255.940 1323.135 1256.220 1327.135 ;
        RECT 1255.960 1313.410 1256.100 1323.135 ;
        RECT 1186.440 1313.090 1186.700 1313.410 ;
        RECT 1255.900 1313.090 1256.160 1313.410 ;
        RECT 1186.500 16.310 1186.640 1313.090 ;
        RECT 1180.000 15.990 1180.260 16.310 ;
        RECT 1186.440 15.990 1186.700 16.310 ;
        RECT 1180.060 2.400 1180.200 15.990 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1200.210 1316.720 1200.530 1316.780 ;
        RECT 1429.750 1316.720 1430.070 1316.780 ;
        RECT 1200.210 1316.580 1430.070 1316.720 ;
        RECT 1200.210 1316.520 1200.530 1316.580 ;
        RECT 1429.750 1316.520 1430.070 1316.580 ;
        RECT 1197.910 16.560 1198.230 16.620 ;
        RECT 1200.210 16.560 1200.530 16.620 ;
        RECT 1197.910 16.420 1200.530 16.560 ;
        RECT 1197.910 16.360 1198.230 16.420 ;
        RECT 1200.210 16.360 1200.530 16.420 ;
      LAYER via ;
        RECT 1200.240 1316.520 1200.500 1316.780 ;
        RECT 1429.780 1316.520 1430.040 1316.780 ;
        RECT 1197.940 16.360 1198.200 16.620 ;
        RECT 1200.240 16.360 1200.500 16.620 ;
      LAYER met2 ;
        RECT 1429.820 1323.135 1430.100 1327.135 ;
        RECT 1429.840 1316.810 1429.980 1323.135 ;
        RECT 1200.240 1316.490 1200.500 1316.810 ;
        RECT 1429.780 1316.490 1430.040 1316.810 ;
        RECT 1200.300 16.650 1200.440 1316.490 ;
        RECT 1197.940 16.330 1198.200 16.650 ;
        RECT 1200.240 16.330 1200.500 16.650 ;
        RECT 1198.000 2.400 1198.140 16.330 ;
        RECT 1197.790 -4.800 1198.350 2.400 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 724.110 1303.460 724.430 1303.520 ;
        RECT 728.710 1303.460 729.030 1303.520 ;
        RECT 724.110 1303.320 729.030 1303.460 ;
        RECT 724.110 1303.260 724.430 1303.320 ;
        RECT 728.710 1303.260 729.030 1303.320 ;
        RECT 728.710 73.340 729.030 73.400 ;
        RECT 1214.930 73.340 1215.250 73.400 ;
        RECT 728.710 73.200 1215.250 73.340 ;
        RECT 728.710 73.140 729.030 73.200 ;
        RECT 1214.930 73.140 1215.250 73.200 ;
      LAYER via ;
        RECT 724.140 1303.260 724.400 1303.520 ;
        RECT 728.740 1303.260 729.000 1303.520 ;
        RECT 728.740 73.140 729.000 73.400 ;
        RECT 1214.960 73.140 1215.220 73.400 ;
      LAYER met2 ;
        RECT 724.180 1323.135 724.460 1327.135 ;
        RECT 724.200 1303.550 724.340 1323.135 ;
        RECT 724.140 1303.230 724.400 1303.550 ;
        RECT 728.740 1303.230 729.000 1303.550 ;
        RECT 728.800 73.430 728.940 1303.230 ;
        RECT 728.740 73.110 729.000 73.430 ;
        RECT 1214.960 73.110 1215.220 73.430 ;
        RECT 1215.020 16.730 1215.160 73.110 ;
        RECT 1215.020 16.590 1216.080 16.730 ;
        RECT 1215.940 2.400 1216.080 16.590 ;
        RECT 1215.730 -4.800 1216.290 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1233.790 24.040 1234.110 24.100 ;
        RECT 1607.770 24.040 1608.090 24.100 ;
        RECT 1233.790 23.900 1608.090 24.040 ;
        RECT 1233.790 23.840 1234.110 23.900 ;
        RECT 1607.770 23.840 1608.090 23.900 ;
      LAYER via ;
        RECT 1233.820 23.840 1234.080 24.100 ;
        RECT 1607.800 23.840 1608.060 24.100 ;
      LAYER met2 ;
        RECT 1609.220 1323.690 1609.500 1327.135 ;
        RECT 1607.860 1323.550 1609.500 1323.690 ;
        RECT 1607.860 24.130 1608.000 1323.550 ;
        RECT 1609.220 1323.135 1609.500 1323.550 ;
        RECT 1233.820 23.810 1234.080 24.130 ;
        RECT 1607.800 23.810 1608.060 24.130 ;
        RECT 1233.880 2.400 1234.020 23.810 ;
        RECT 1233.670 -4.800 1234.230 2.400 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1251.730 30.500 1252.050 30.560 ;
        RECT 1725.070 30.500 1725.390 30.560 ;
        RECT 1251.730 30.360 1725.390 30.500 ;
        RECT 1251.730 30.300 1252.050 30.360 ;
        RECT 1725.070 30.300 1725.390 30.360 ;
      LAYER via ;
        RECT 1251.760 30.300 1252.020 30.560 ;
        RECT 1725.100 30.300 1725.360 30.560 ;
      LAYER met2 ;
        RECT 1725.140 1323.135 1725.420 1327.135 ;
        RECT 1725.160 30.590 1725.300 1323.135 ;
        RECT 1251.760 30.270 1252.020 30.590 ;
        RECT 1725.100 30.270 1725.360 30.590 ;
        RECT 1251.820 2.400 1251.960 30.270 ;
        RECT 1251.610 -4.800 1252.170 2.400 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 695.590 2374.800 695.910 2374.860 ;
        RECT 956.870 2374.800 957.190 2374.860 ;
        RECT 695.590 2374.660 957.190 2374.800 ;
        RECT 695.590 2374.600 695.910 2374.660 ;
        RECT 956.870 2374.600 957.190 2374.660 ;
        RECT 695.590 16.900 695.910 16.960 ;
        RECT 1269.210 16.900 1269.530 16.960 ;
        RECT 695.590 16.760 1269.530 16.900 ;
        RECT 695.590 16.700 695.910 16.760 ;
        RECT 1269.210 16.700 1269.530 16.760 ;
      LAYER via ;
        RECT 695.620 2374.600 695.880 2374.860 ;
        RECT 956.900 2374.600 957.160 2374.860 ;
        RECT 695.620 16.700 695.880 16.960 ;
        RECT 1269.240 16.700 1269.500 16.960 ;
      LAYER met2 ;
        RECT 958.780 2374.970 959.060 2377.880 ;
        RECT 956.960 2374.890 959.060 2374.970 ;
        RECT 695.620 2374.570 695.880 2374.890 ;
        RECT 956.900 2374.830 959.060 2374.890 ;
        RECT 956.900 2374.570 957.160 2374.830 ;
        RECT 695.680 1393.845 695.820 2374.570 ;
        RECT 958.780 2373.880 959.060 2374.830 ;
        RECT 695.610 1393.475 695.890 1393.845 ;
        RECT 695.610 1390.755 695.890 1391.125 ;
        RECT 695.680 16.990 695.820 1390.755 ;
        RECT 695.620 16.670 695.880 16.990 ;
        RECT 1269.240 16.670 1269.500 16.990 ;
        RECT 1269.300 2.400 1269.440 16.670 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
      LAYER via2 ;
        RECT 695.610 1393.520 695.890 1393.800 ;
        RECT 695.610 1390.800 695.890 1391.080 ;
      LAYER met3 ;
        RECT 695.585 1393.810 695.915 1393.825 ;
        RECT 695.585 1393.495 696.130 1393.810 ;
        RECT 695.830 1391.105 696.130 1393.495 ;
        RECT 695.585 1390.790 696.130 1391.105 ;
        RECT 695.585 1390.775 695.915 1390.790 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 762.365 18.105 762.535 20.315 ;
        RECT 786.285 18.105 786.455 21.335 ;
        RECT 927.505 15.045 927.675 20.315 ;
        RECT 1052.165 15.045 1052.335 20.655 ;
        RECT 1131.745 15.385 1131.915 20.315 ;
        RECT 1192.925 15.385 1193.095 20.315 ;
      LAYER mcon ;
        RECT 786.285 21.165 786.455 21.335 ;
        RECT 762.365 20.145 762.535 20.315 ;
        RECT 1052.165 20.485 1052.335 20.655 ;
        RECT 927.505 20.145 927.675 20.315 ;
        RECT 1131.745 20.145 1131.915 20.315 ;
        RECT 1192.925 20.145 1193.095 20.315 ;
      LAYER met1 ;
        RECT 702.490 2375.820 702.810 2375.880 ;
        RECT 876.370 2375.820 876.690 2375.880 ;
        RECT 702.490 2375.680 876.690 2375.820 ;
        RECT 702.490 2375.620 702.810 2375.680 ;
        RECT 876.370 2375.620 876.690 2375.680 ;
        RECT 786.225 21.320 786.515 21.365 ;
        RECT 786.225 21.180 787.360 21.320 ;
        RECT 786.225 21.135 786.515 21.180 ;
        RECT 702.490 20.300 702.810 20.360 ;
        RECT 762.305 20.300 762.595 20.345 ;
        RECT 702.490 20.160 762.595 20.300 ;
        RECT 787.220 20.300 787.360 21.180 ;
        RECT 1052.105 20.640 1052.395 20.685 ;
        RECT 1052.105 20.500 1084.980 20.640 ;
        RECT 1052.105 20.455 1052.395 20.500 ;
        RECT 927.445 20.300 927.735 20.345 ;
        RECT 787.220 20.160 927.735 20.300 ;
        RECT 1084.840 20.300 1084.980 20.500 ;
        RECT 1131.685 20.300 1131.975 20.345 ;
        RECT 1084.840 20.160 1131.975 20.300 ;
        RECT 702.490 20.100 702.810 20.160 ;
        RECT 762.305 20.115 762.595 20.160 ;
        RECT 927.445 20.115 927.735 20.160 ;
        RECT 1131.685 20.115 1131.975 20.160 ;
        RECT 1192.865 20.300 1193.155 20.345 ;
        RECT 1287.150 20.300 1287.470 20.360 ;
        RECT 1192.865 20.160 1287.470 20.300 ;
        RECT 1192.865 20.115 1193.155 20.160 ;
        RECT 1287.150 20.100 1287.470 20.160 ;
        RECT 762.305 18.260 762.595 18.305 ;
        RECT 786.225 18.260 786.515 18.305 ;
        RECT 762.305 18.120 786.515 18.260 ;
        RECT 762.305 18.075 762.595 18.120 ;
        RECT 786.225 18.075 786.515 18.120 ;
        RECT 1131.685 15.540 1131.975 15.585 ;
        RECT 1192.865 15.540 1193.155 15.585 ;
        RECT 1131.685 15.400 1193.155 15.540 ;
        RECT 1131.685 15.355 1131.975 15.400 ;
        RECT 1192.865 15.355 1193.155 15.400 ;
        RECT 927.445 15.200 927.735 15.245 ;
        RECT 1052.105 15.200 1052.395 15.245 ;
        RECT 927.445 15.060 1052.395 15.200 ;
        RECT 927.445 15.015 927.735 15.060 ;
        RECT 1052.105 15.015 1052.395 15.060 ;
      LAYER via ;
        RECT 702.520 2375.620 702.780 2375.880 ;
        RECT 876.400 2375.620 876.660 2375.880 ;
        RECT 702.520 20.100 702.780 20.360 ;
        RECT 1287.180 20.100 1287.440 20.360 ;
      LAYER met2 ;
        RECT 702.520 2375.590 702.780 2375.910 ;
        RECT 876.400 2375.650 876.660 2375.910 ;
        RECT 877.820 2375.650 878.100 2377.880 ;
        RECT 876.400 2375.590 878.100 2375.650 ;
        RECT 702.580 20.390 702.720 2375.590 ;
        RECT 876.460 2375.510 878.100 2375.590 ;
        RECT 877.820 2373.880 878.100 2375.510 ;
        RECT 702.520 20.070 702.780 20.390 ;
        RECT 1287.180 20.070 1287.440 20.390 ;
        RECT 1287.240 2.400 1287.380 20.070 ;
        RECT 1287.030 -4.800 1287.590 2.400 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 682.710 2379.560 683.030 2379.620 ;
        RECT 773.790 2379.560 774.110 2379.620 ;
        RECT 682.710 2379.420 774.110 2379.560 ;
        RECT 682.710 2379.360 683.030 2379.420 ;
        RECT 773.790 2379.360 774.110 2379.420 ;
        RECT 682.710 34.240 683.030 34.300 ;
        RECT 1305.090 34.240 1305.410 34.300 ;
        RECT 682.710 34.100 1305.410 34.240 ;
        RECT 682.710 34.040 683.030 34.100 ;
        RECT 1305.090 34.040 1305.410 34.100 ;
      LAYER via ;
        RECT 682.740 2379.360 683.000 2379.620 ;
        RECT 773.820 2379.360 774.080 2379.620 ;
        RECT 682.740 34.040 683.000 34.300 ;
        RECT 1305.120 34.040 1305.380 34.300 ;
      LAYER met2 ;
        RECT 682.740 2379.330 683.000 2379.650 ;
        RECT 773.820 2379.330 774.080 2379.650 ;
        RECT 682.800 34.330 682.940 2379.330 ;
        RECT 773.880 2377.880 774.020 2379.330 ;
        RECT 773.860 2373.880 774.140 2377.880 ;
        RECT 682.740 34.010 683.000 34.330 ;
        RECT 1305.120 34.010 1305.380 34.330 ;
        RECT 1305.180 2.400 1305.320 34.010 ;
        RECT 1304.970 -4.800 1305.530 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 708.010 1553.020 708.330 1553.080 ;
        RECT 720.430 1553.020 720.750 1553.080 ;
        RECT 708.010 1552.880 720.750 1553.020 ;
        RECT 708.010 1552.820 708.330 1552.880 ;
        RECT 720.430 1552.820 720.750 1552.880 ;
        RECT 720.430 19.960 720.750 20.020 ;
        RECT 1323.030 19.960 1323.350 20.020 ;
        RECT 720.430 19.820 1323.350 19.960 ;
        RECT 720.430 19.760 720.750 19.820 ;
        RECT 1323.030 19.760 1323.350 19.820 ;
      LAYER via ;
        RECT 708.040 1552.820 708.300 1553.080 ;
        RECT 720.460 1552.820 720.720 1553.080 ;
        RECT 720.460 19.760 720.720 20.020 ;
        RECT 1323.060 19.760 1323.320 20.020 ;
      LAYER met2 ;
        RECT 708.030 2087.755 708.310 2088.125 ;
        RECT 708.100 1553.110 708.240 2087.755 ;
        RECT 708.040 1552.790 708.300 1553.110 ;
        RECT 720.460 1552.790 720.720 1553.110 ;
        RECT 720.520 1525.650 720.660 1552.790 ;
        RECT 720.060 1525.510 720.660 1525.650 ;
        RECT 720.060 1521.570 720.200 1525.510 ;
        RECT 720.060 1521.430 720.660 1521.570 ;
        RECT 720.520 20.050 720.660 1521.430 ;
        RECT 720.460 19.730 720.720 20.050 ;
        RECT 1323.060 19.730 1323.320 20.050 ;
        RECT 1323.120 2.400 1323.260 19.730 ;
        RECT 1322.910 -4.800 1323.470 2.400 ;
      LAYER via2 ;
        RECT 708.030 2087.800 708.310 2088.080 ;
      LAYER met3 ;
        RECT 708.005 2088.090 708.335 2088.105 ;
        RECT 715.810 2088.090 719.810 2088.095 ;
        RECT 708.005 2087.790 719.810 2088.090 ;
        RECT 708.005 2087.775 708.335 2087.790 ;
        RECT 715.810 2087.495 719.810 2087.790 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1338.745 1304.325 1338.915 1309.935 ;
        RECT 1338.745 1207.425 1338.915 1255.875 ;
        RECT 1338.745 531.505 1338.915 579.615 ;
        RECT 1338.745 434.945 1338.915 483.055 ;
        RECT 1338.745 338.045 1338.915 386.155 ;
        RECT 1338.745 241.485 1338.915 289.595 ;
        RECT 1338.745 144.925 1338.915 193.035 ;
        RECT 1340.585 2.805 1340.755 48.195 ;
      LAYER mcon ;
        RECT 1338.745 1309.765 1338.915 1309.935 ;
        RECT 1338.745 1255.705 1338.915 1255.875 ;
        RECT 1338.745 579.445 1338.915 579.615 ;
        RECT 1338.745 482.885 1338.915 483.055 ;
        RECT 1338.745 385.985 1338.915 386.155 ;
        RECT 1338.745 289.425 1338.915 289.595 ;
        RECT 1338.745 192.865 1338.915 193.035 ;
        RECT 1340.585 48.025 1340.755 48.195 ;
      LAYER met1 ;
        RECT 718.130 1309.920 718.450 1309.980 ;
        RECT 1338.685 1309.920 1338.975 1309.965 ;
        RECT 718.130 1309.780 1338.975 1309.920 ;
        RECT 718.130 1309.720 718.450 1309.780 ;
        RECT 1338.685 1309.735 1338.975 1309.780 ;
        RECT 1338.670 1304.480 1338.990 1304.540 ;
        RECT 1338.475 1304.340 1338.990 1304.480 ;
        RECT 1338.670 1304.280 1338.990 1304.340 ;
        RECT 1338.670 1255.860 1338.990 1255.920 ;
        RECT 1338.475 1255.720 1338.990 1255.860 ;
        RECT 1338.670 1255.660 1338.990 1255.720 ;
        RECT 1338.670 1207.580 1338.990 1207.640 ;
        RECT 1338.475 1207.440 1338.990 1207.580 ;
        RECT 1338.670 1207.380 1338.990 1207.440 ;
        RECT 1338.670 1111.020 1338.990 1111.080 ;
        RECT 1339.590 1111.020 1339.910 1111.080 ;
        RECT 1338.670 1110.880 1339.910 1111.020 ;
        RECT 1338.670 1110.820 1338.990 1110.880 ;
        RECT 1339.590 1110.820 1339.910 1110.880 ;
        RECT 1338.670 1014.460 1338.990 1014.520 ;
        RECT 1339.590 1014.460 1339.910 1014.520 ;
        RECT 1338.670 1014.320 1339.910 1014.460 ;
        RECT 1338.670 1014.260 1338.990 1014.320 ;
        RECT 1339.590 1014.260 1339.910 1014.320 ;
        RECT 1338.670 917.900 1338.990 917.960 ;
        RECT 1339.590 917.900 1339.910 917.960 ;
        RECT 1338.670 917.760 1339.910 917.900 ;
        RECT 1338.670 917.700 1338.990 917.760 ;
        RECT 1339.590 917.700 1339.910 917.760 ;
        RECT 1338.670 772.720 1338.990 772.780 ;
        RECT 1339.590 772.720 1339.910 772.780 ;
        RECT 1338.670 772.580 1339.910 772.720 ;
        RECT 1338.670 772.520 1338.990 772.580 ;
        RECT 1339.590 772.520 1339.910 772.580 ;
        RECT 1338.670 676.160 1338.990 676.220 ;
        RECT 1339.590 676.160 1339.910 676.220 ;
        RECT 1338.670 676.020 1339.910 676.160 ;
        RECT 1338.670 675.960 1338.990 676.020 ;
        RECT 1339.590 675.960 1339.910 676.020 ;
        RECT 1338.670 579.600 1338.990 579.660 ;
        RECT 1338.475 579.460 1338.990 579.600 ;
        RECT 1338.670 579.400 1338.990 579.460 ;
        RECT 1338.670 531.660 1338.990 531.720 ;
        RECT 1338.475 531.520 1338.990 531.660 ;
        RECT 1338.670 531.460 1338.990 531.520 ;
        RECT 1338.670 483.040 1338.990 483.100 ;
        RECT 1338.475 482.900 1338.990 483.040 ;
        RECT 1338.670 482.840 1338.990 482.900 ;
        RECT 1338.670 435.100 1338.990 435.160 ;
        RECT 1338.475 434.960 1338.990 435.100 ;
        RECT 1338.670 434.900 1338.990 434.960 ;
        RECT 1338.670 386.140 1338.990 386.200 ;
        RECT 1338.475 386.000 1338.990 386.140 ;
        RECT 1338.670 385.940 1338.990 386.000 ;
        RECT 1338.670 338.200 1338.990 338.260 ;
        RECT 1338.475 338.060 1338.990 338.200 ;
        RECT 1338.670 338.000 1338.990 338.060 ;
        RECT 1338.670 289.580 1338.990 289.640 ;
        RECT 1338.475 289.440 1338.990 289.580 ;
        RECT 1338.670 289.380 1338.990 289.440 ;
        RECT 1338.670 241.640 1338.990 241.700 ;
        RECT 1338.475 241.500 1338.990 241.640 ;
        RECT 1338.670 241.440 1338.990 241.500 ;
        RECT 1338.670 193.020 1338.990 193.080 ;
        RECT 1338.475 192.880 1338.990 193.020 ;
        RECT 1338.670 192.820 1338.990 192.880 ;
        RECT 1338.670 145.080 1338.990 145.140 ;
        RECT 1338.475 144.940 1338.990 145.080 ;
        RECT 1338.670 144.880 1338.990 144.940 ;
        RECT 1337.750 96.460 1338.070 96.520 ;
        RECT 1338.670 96.460 1338.990 96.520 ;
        RECT 1337.750 96.320 1338.990 96.460 ;
        RECT 1337.750 96.260 1338.070 96.320 ;
        RECT 1338.670 96.260 1338.990 96.320 ;
        RECT 1338.670 48.180 1338.990 48.240 ;
        RECT 1340.525 48.180 1340.815 48.225 ;
        RECT 1338.670 48.040 1340.815 48.180 ;
        RECT 1338.670 47.980 1338.990 48.040 ;
        RECT 1340.525 47.995 1340.815 48.040 ;
        RECT 1340.510 2.960 1340.830 3.020 ;
        RECT 1340.315 2.820 1340.830 2.960 ;
        RECT 1340.510 2.760 1340.830 2.820 ;
      LAYER via ;
        RECT 718.160 1309.720 718.420 1309.980 ;
        RECT 1338.700 1304.280 1338.960 1304.540 ;
        RECT 1338.700 1255.660 1338.960 1255.920 ;
        RECT 1338.700 1207.380 1338.960 1207.640 ;
        RECT 1338.700 1110.820 1338.960 1111.080 ;
        RECT 1339.620 1110.820 1339.880 1111.080 ;
        RECT 1338.700 1014.260 1338.960 1014.520 ;
        RECT 1339.620 1014.260 1339.880 1014.520 ;
        RECT 1338.700 917.700 1338.960 917.960 ;
        RECT 1339.620 917.700 1339.880 917.960 ;
        RECT 1338.700 772.520 1338.960 772.780 ;
        RECT 1339.620 772.520 1339.880 772.780 ;
        RECT 1338.700 675.960 1338.960 676.220 ;
        RECT 1339.620 675.960 1339.880 676.220 ;
        RECT 1338.700 579.400 1338.960 579.660 ;
        RECT 1338.700 531.460 1338.960 531.720 ;
        RECT 1338.700 482.840 1338.960 483.100 ;
        RECT 1338.700 434.900 1338.960 435.160 ;
        RECT 1338.700 385.940 1338.960 386.200 ;
        RECT 1338.700 338.000 1338.960 338.260 ;
        RECT 1338.700 289.380 1338.960 289.640 ;
        RECT 1338.700 241.440 1338.960 241.700 ;
        RECT 1338.700 192.820 1338.960 193.080 ;
        RECT 1338.700 144.880 1338.960 145.140 ;
        RECT 1337.780 96.260 1338.040 96.520 ;
        RECT 1338.700 96.260 1338.960 96.520 ;
        RECT 1338.700 47.980 1338.960 48.240 ;
        RECT 1340.540 2.760 1340.800 3.020 ;
      LAYER met2 ;
        RECT 717.690 1855.195 717.970 1855.565 ;
        RECT 717.760 1354.970 717.900 1855.195 ;
        RECT 717.760 1354.830 718.360 1354.970 ;
        RECT 718.220 1310.010 718.360 1354.830 ;
        RECT 718.160 1309.690 718.420 1310.010 ;
        RECT 1338.700 1304.250 1338.960 1304.570 ;
        RECT 1338.760 1255.950 1338.900 1304.250 ;
        RECT 1338.700 1255.630 1338.960 1255.950 ;
        RECT 1338.700 1207.350 1338.960 1207.670 ;
        RECT 1338.760 1159.245 1338.900 1207.350 ;
        RECT 1338.690 1158.875 1338.970 1159.245 ;
        RECT 1339.610 1158.875 1339.890 1159.245 ;
        RECT 1339.680 1111.110 1339.820 1158.875 ;
        RECT 1338.700 1110.790 1338.960 1111.110 ;
        RECT 1339.620 1110.790 1339.880 1111.110 ;
        RECT 1338.760 1062.685 1338.900 1110.790 ;
        RECT 1338.690 1062.315 1338.970 1062.685 ;
        RECT 1339.610 1062.315 1339.890 1062.685 ;
        RECT 1339.680 1014.550 1339.820 1062.315 ;
        RECT 1338.700 1014.230 1338.960 1014.550 ;
        RECT 1339.620 1014.230 1339.880 1014.550 ;
        RECT 1338.760 966.125 1338.900 1014.230 ;
        RECT 1338.690 965.755 1338.970 966.125 ;
        RECT 1339.610 965.755 1339.890 966.125 ;
        RECT 1339.680 917.990 1339.820 965.755 ;
        RECT 1338.700 917.670 1338.960 917.990 ;
        RECT 1339.620 917.670 1339.880 917.990 ;
        RECT 1338.760 869.565 1338.900 917.670 ;
        RECT 1338.690 869.195 1338.970 869.565 ;
        RECT 1339.610 869.195 1339.890 869.565 ;
        RECT 1339.680 821.285 1339.820 869.195 ;
        RECT 1338.690 820.915 1338.970 821.285 ;
        RECT 1339.610 820.915 1339.890 821.285 ;
        RECT 1338.760 772.810 1338.900 820.915 ;
        RECT 1338.700 772.490 1338.960 772.810 ;
        RECT 1339.620 772.490 1339.880 772.810 ;
        RECT 1339.680 724.725 1339.820 772.490 ;
        RECT 1338.690 724.355 1338.970 724.725 ;
        RECT 1339.610 724.355 1339.890 724.725 ;
        RECT 1338.760 676.250 1338.900 724.355 ;
        RECT 1338.700 675.930 1338.960 676.250 ;
        RECT 1339.620 675.930 1339.880 676.250 ;
        RECT 1339.680 628.165 1339.820 675.930 ;
        RECT 1338.690 627.795 1338.970 628.165 ;
        RECT 1339.610 627.795 1339.890 628.165 ;
        RECT 1338.760 579.690 1338.900 627.795 ;
        RECT 1338.700 579.370 1338.960 579.690 ;
        RECT 1338.700 531.430 1338.960 531.750 ;
        RECT 1338.760 483.130 1338.900 531.430 ;
        RECT 1338.700 482.810 1338.960 483.130 ;
        RECT 1338.700 434.870 1338.960 435.190 ;
        RECT 1338.760 386.230 1338.900 434.870 ;
        RECT 1338.700 385.910 1338.960 386.230 ;
        RECT 1338.700 337.970 1338.960 338.290 ;
        RECT 1338.760 289.670 1338.900 337.970 ;
        RECT 1338.700 289.350 1338.960 289.670 ;
        RECT 1338.700 241.410 1338.960 241.730 ;
        RECT 1338.760 193.110 1338.900 241.410 ;
        RECT 1338.700 192.790 1338.960 193.110 ;
        RECT 1338.700 144.850 1338.960 145.170 ;
        RECT 1338.760 96.550 1338.900 144.850 ;
        RECT 1337.780 96.230 1338.040 96.550 ;
        RECT 1338.700 96.230 1338.960 96.550 ;
        RECT 1337.840 48.805 1337.980 96.230 ;
        RECT 1337.770 48.435 1338.050 48.805 ;
        RECT 1338.690 48.435 1338.970 48.805 ;
        RECT 1338.760 48.270 1338.900 48.435 ;
        RECT 1338.700 47.950 1338.960 48.270 ;
        RECT 1340.540 2.730 1340.800 3.050 ;
        RECT 1340.600 2.400 1340.740 2.730 ;
        RECT 1340.390 -4.800 1340.950 2.400 ;
      LAYER via2 ;
        RECT 717.690 1855.240 717.970 1855.520 ;
        RECT 1338.690 1158.920 1338.970 1159.200 ;
        RECT 1339.610 1158.920 1339.890 1159.200 ;
        RECT 1338.690 1062.360 1338.970 1062.640 ;
        RECT 1339.610 1062.360 1339.890 1062.640 ;
        RECT 1338.690 965.800 1338.970 966.080 ;
        RECT 1339.610 965.800 1339.890 966.080 ;
        RECT 1338.690 869.240 1338.970 869.520 ;
        RECT 1339.610 869.240 1339.890 869.520 ;
        RECT 1338.690 820.960 1338.970 821.240 ;
        RECT 1339.610 820.960 1339.890 821.240 ;
        RECT 1338.690 724.400 1338.970 724.680 ;
        RECT 1339.610 724.400 1339.890 724.680 ;
        RECT 1338.690 627.840 1338.970 628.120 ;
        RECT 1339.610 627.840 1339.890 628.120 ;
        RECT 1337.770 48.480 1338.050 48.760 ;
        RECT 1338.690 48.480 1338.970 48.760 ;
      LAYER met3 ;
        RECT 715.810 1856.295 719.810 1856.895 ;
        RECT 717.910 1855.545 718.210 1856.295 ;
        RECT 717.665 1855.230 718.210 1855.545 ;
        RECT 717.665 1855.215 717.995 1855.230 ;
        RECT 1338.665 1159.210 1338.995 1159.225 ;
        RECT 1339.585 1159.210 1339.915 1159.225 ;
        RECT 1338.665 1158.910 1339.915 1159.210 ;
        RECT 1338.665 1158.895 1338.995 1158.910 ;
        RECT 1339.585 1158.895 1339.915 1158.910 ;
        RECT 1338.665 1062.650 1338.995 1062.665 ;
        RECT 1339.585 1062.650 1339.915 1062.665 ;
        RECT 1338.665 1062.350 1339.915 1062.650 ;
        RECT 1338.665 1062.335 1338.995 1062.350 ;
        RECT 1339.585 1062.335 1339.915 1062.350 ;
        RECT 1338.665 966.090 1338.995 966.105 ;
        RECT 1339.585 966.090 1339.915 966.105 ;
        RECT 1338.665 965.790 1339.915 966.090 ;
        RECT 1338.665 965.775 1338.995 965.790 ;
        RECT 1339.585 965.775 1339.915 965.790 ;
        RECT 1338.665 869.530 1338.995 869.545 ;
        RECT 1339.585 869.530 1339.915 869.545 ;
        RECT 1338.665 869.230 1339.915 869.530 ;
        RECT 1338.665 869.215 1338.995 869.230 ;
        RECT 1339.585 869.215 1339.915 869.230 ;
        RECT 1338.665 821.250 1338.995 821.265 ;
        RECT 1339.585 821.250 1339.915 821.265 ;
        RECT 1338.665 820.950 1339.915 821.250 ;
        RECT 1338.665 820.935 1338.995 820.950 ;
        RECT 1339.585 820.935 1339.915 820.950 ;
        RECT 1338.665 724.690 1338.995 724.705 ;
        RECT 1339.585 724.690 1339.915 724.705 ;
        RECT 1338.665 724.390 1339.915 724.690 ;
        RECT 1338.665 724.375 1338.995 724.390 ;
        RECT 1339.585 724.375 1339.915 724.390 ;
        RECT 1338.665 628.130 1338.995 628.145 ;
        RECT 1339.585 628.130 1339.915 628.145 ;
        RECT 1338.665 627.830 1339.915 628.130 ;
        RECT 1338.665 627.815 1338.995 627.830 ;
        RECT 1339.585 627.815 1339.915 627.830 ;
        RECT 1337.745 48.770 1338.075 48.785 ;
        RECT 1338.665 48.770 1338.995 48.785 ;
        RECT 1337.745 48.470 1338.995 48.770 ;
        RECT 1337.745 48.455 1338.075 48.470 ;
        RECT 1338.665 48.455 1338.995 48.470 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 698.350 61.440 698.670 61.500 ;
        RECT 1760.030 61.440 1760.350 61.500 ;
        RECT 698.350 61.300 1760.350 61.440 ;
        RECT 698.350 61.240 698.670 61.300 ;
        RECT 1760.030 61.240 1760.350 61.300 ;
      LAYER via ;
        RECT 698.380 61.240 698.640 61.500 ;
        RECT 1760.060 61.240 1760.320 61.500 ;
      LAYER met2 ;
        RECT 1760.050 2063.275 1760.330 2063.645 ;
        RECT 1760.120 61.530 1760.260 2063.275 ;
        RECT 698.380 61.210 698.640 61.530 ;
        RECT 1760.060 61.210 1760.320 61.530 ;
        RECT 698.440 2.400 698.580 61.210 ;
        RECT 698.230 -4.800 698.790 2.400 ;
      LAYER via2 ;
        RECT 1760.050 2063.320 1760.330 2063.600 ;
      LAYER met3 ;
        RECT 1755.835 2065.735 1759.835 2066.335 ;
        RECT 1759.350 2063.610 1759.650 2065.735 ;
        RECT 1760.025 2063.610 1760.355 2063.625 ;
        RECT 1759.350 2063.310 1760.355 2063.610 ;
        RECT 1760.025 2063.295 1760.355 2063.310 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1358.450 196.760 1358.770 196.820 ;
        RECT 1759.570 196.760 1759.890 196.820 ;
        RECT 1358.450 196.620 1759.890 196.760 ;
        RECT 1358.450 196.560 1358.770 196.620 ;
        RECT 1759.570 196.560 1759.890 196.620 ;
      LAYER via ;
        RECT 1358.480 196.560 1358.740 196.820 ;
        RECT 1759.600 196.560 1759.860 196.820 ;
      LAYER met2 ;
        RECT 1759.590 2227.835 1759.870 2228.205 ;
        RECT 1759.660 196.850 1759.800 2227.835 ;
        RECT 1358.480 196.530 1358.740 196.850 ;
        RECT 1759.600 196.530 1759.860 196.850 ;
        RECT 1358.540 2.400 1358.680 196.530 ;
        RECT 1358.330 -4.800 1358.890 2.400 ;
      LAYER via2 ;
        RECT 1759.590 2227.880 1759.870 2228.160 ;
      LAYER met3 ;
        RECT 1755.835 2228.935 1759.835 2229.535 ;
        RECT 1759.350 2228.185 1759.650 2228.935 ;
        RECT 1759.350 2227.870 1759.895 2228.185 ;
        RECT 1759.565 2227.855 1759.895 2227.870 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1633.145 2387.905 1633.315 2389.435 ;
      LAYER mcon ;
        RECT 1633.145 2389.265 1633.315 2389.435 ;
      LAYER met1 ;
        RECT 1611.910 2389.420 1612.230 2389.480 ;
        RECT 1633.085 2389.420 1633.375 2389.465 ;
        RECT 1611.910 2389.280 1633.375 2389.420 ;
        RECT 1611.910 2389.220 1612.230 2389.280 ;
        RECT 1633.085 2389.235 1633.375 2389.280 ;
        RECT 1633.085 2388.060 1633.375 2388.105 ;
        RECT 1781.650 2388.060 1781.970 2388.120 ;
        RECT 1633.085 2387.920 1781.970 2388.060 ;
        RECT 1633.085 2387.875 1633.375 2387.920 ;
        RECT 1781.650 2387.860 1781.970 2387.920 ;
        RECT 1379.610 1323.520 1379.930 1323.580 ;
        RECT 1781.650 1323.520 1781.970 1323.580 ;
        RECT 1379.610 1323.380 1781.970 1323.520 ;
        RECT 1379.610 1323.320 1379.930 1323.380 ;
        RECT 1781.650 1323.320 1781.970 1323.380 ;
        RECT 1376.390 20.640 1376.710 20.700 ;
        RECT 1379.610 20.640 1379.930 20.700 ;
        RECT 1376.390 20.500 1379.930 20.640 ;
        RECT 1376.390 20.440 1376.710 20.500 ;
        RECT 1379.610 20.440 1379.930 20.500 ;
      LAYER via ;
        RECT 1611.940 2389.220 1612.200 2389.480 ;
        RECT 1781.680 2387.860 1781.940 2388.120 ;
        RECT 1379.640 1323.320 1379.900 1323.580 ;
        RECT 1781.680 1323.320 1781.940 1323.580 ;
        RECT 1376.420 20.440 1376.680 20.700 ;
        RECT 1379.640 20.440 1379.900 20.700 ;
      LAYER met2 ;
        RECT 1611.940 2389.190 1612.200 2389.510 ;
        RECT 1612.000 2377.880 1612.140 2389.190 ;
        RECT 1781.680 2387.830 1781.940 2388.150 ;
        RECT 1611.980 2373.880 1612.260 2377.880 ;
        RECT 1781.740 1323.610 1781.880 2387.830 ;
        RECT 1379.640 1323.290 1379.900 1323.610 ;
        RECT 1781.680 1323.290 1781.940 1323.610 ;
        RECT 1379.700 20.730 1379.840 1323.290 ;
        RECT 1376.420 20.410 1376.680 20.730 ;
        RECT 1379.640 20.410 1379.900 20.730 ;
        RECT 1376.480 2.400 1376.620 20.410 ;
        RECT 1376.270 -4.800 1376.830 2.400 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1763.785 1341.045 1763.955 1342.575 ;
      LAYER mcon ;
        RECT 1763.785 1342.405 1763.955 1342.575 ;
      LAYER met1 ;
        RECT 1763.710 1342.560 1764.030 1342.620 ;
        RECT 1763.515 1342.420 1764.030 1342.560 ;
        RECT 1763.710 1342.360 1764.030 1342.420 ;
        RECT 1763.710 1341.200 1764.030 1341.260 ;
        RECT 1763.515 1341.060 1764.030 1341.200 ;
        RECT 1763.710 1341.000 1764.030 1341.060 ;
        RECT 1399.850 1280.340 1400.170 1280.400 ;
        RECT 1763.710 1280.340 1764.030 1280.400 ;
        RECT 1399.850 1280.200 1764.030 1280.340 ;
        RECT 1399.850 1280.140 1400.170 1280.200 ;
        RECT 1763.710 1280.140 1764.030 1280.200 ;
        RECT 1394.330 16.220 1394.650 16.280 ;
        RECT 1399.850 16.220 1400.170 16.280 ;
        RECT 1394.330 16.080 1400.170 16.220 ;
        RECT 1394.330 16.020 1394.650 16.080 ;
        RECT 1399.850 16.020 1400.170 16.080 ;
      LAYER via ;
        RECT 1763.740 1342.360 1764.000 1342.620 ;
        RECT 1763.740 1341.000 1764.000 1341.260 ;
        RECT 1399.880 1280.140 1400.140 1280.400 ;
        RECT 1763.740 1280.140 1764.000 1280.400 ;
        RECT 1394.360 16.020 1394.620 16.280 ;
        RECT 1399.880 16.020 1400.140 16.280 ;
      LAYER met2 ;
        RECT 1763.730 2083.675 1764.010 2084.045 ;
        RECT 1763.800 1342.650 1763.940 2083.675 ;
        RECT 1763.740 1342.330 1764.000 1342.650 ;
        RECT 1763.740 1340.970 1764.000 1341.290 ;
        RECT 1763.800 1280.430 1763.940 1340.970 ;
        RECT 1399.880 1280.110 1400.140 1280.430 ;
        RECT 1763.740 1280.110 1764.000 1280.430 ;
        RECT 1399.940 16.310 1400.080 1280.110 ;
        RECT 1394.360 15.990 1394.620 16.310 ;
        RECT 1399.880 15.990 1400.140 16.310 ;
        RECT 1394.420 2.400 1394.560 15.990 ;
        RECT 1394.210 -4.800 1394.770 2.400 ;
      LAYER via2 ;
        RECT 1763.730 2083.720 1764.010 2084.000 ;
      LAYER met3 ;
        RECT 1755.835 2084.010 1759.835 2084.015 ;
        RECT 1763.705 2084.010 1764.035 2084.025 ;
        RECT 1755.835 2083.710 1764.035 2084.010 ;
        RECT 1755.835 2083.415 1759.835 2083.710 ;
        RECT 1763.705 2083.695 1764.035 2083.710 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 689.610 2366.980 689.930 2367.040 ;
        RECT 709.390 2366.980 709.710 2367.040 ;
        RECT 689.610 2366.840 709.710 2366.980 ;
        RECT 689.610 2366.780 689.930 2366.840 ;
        RECT 709.390 2366.780 709.710 2366.840 ;
        RECT 689.610 33.900 689.930 33.960 ;
        RECT 1412.270 33.900 1412.590 33.960 ;
        RECT 689.610 33.760 1412.590 33.900 ;
        RECT 689.610 33.700 689.930 33.760 ;
        RECT 1412.270 33.700 1412.590 33.760 ;
      LAYER via ;
        RECT 689.640 2366.780 689.900 2367.040 ;
        RECT 709.420 2366.780 709.680 2367.040 ;
        RECT 689.640 33.700 689.900 33.960 ;
        RECT 1412.300 33.700 1412.560 33.960 ;
      LAYER met2 ;
        RECT 709.410 2370.635 709.690 2371.005 ;
        RECT 709.480 2367.070 709.620 2370.635 ;
        RECT 689.640 2366.750 689.900 2367.070 ;
        RECT 709.420 2366.750 709.680 2367.070 ;
        RECT 689.700 33.990 689.840 2366.750 ;
        RECT 689.640 33.670 689.900 33.990 ;
        RECT 1412.300 33.670 1412.560 33.990 ;
        RECT 1412.360 2.400 1412.500 33.670 ;
        RECT 1412.150 -4.800 1412.710 2.400 ;
      LAYER via2 ;
        RECT 709.410 2370.680 709.690 2370.960 ;
      LAYER met3 ;
        RECT 709.385 2370.970 709.715 2370.985 ;
        RECT 715.810 2370.970 719.810 2370.975 ;
        RECT 709.385 2370.670 719.810 2370.970 ;
        RECT 709.385 2370.655 709.715 2370.670 ;
        RECT 715.810 2370.375 719.810 2370.670 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1755.965 1313.165 1756.135 1329.995 ;
      LAYER mcon ;
        RECT 1755.965 1329.825 1756.135 1329.995 ;
      LAYER met1 ;
        RECT 1755.905 1329.980 1756.195 1330.025 ;
        RECT 1756.350 1329.980 1756.670 1330.040 ;
        RECT 1755.905 1329.840 1756.670 1329.980 ;
        RECT 1755.905 1329.795 1756.195 1329.840 ;
        RECT 1756.350 1329.780 1756.670 1329.840 ;
        RECT 1434.810 1313.320 1435.130 1313.380 ;
        RECT 1755.905 1313.320 1756.195 1313.365 ;
        RECT 1434.810 1313.180 1756.195 1313.320 ;
        RECT 1434.810 1313.120 1435.130 1313.180 ;
        RECT 1755.905 1313.135 1756.195 1313.180 ;
        RECT 1429.750 16.900 1430.070 16.960 ;
        RECT 1434.810 16.900 1435.130 16.960 ;
        RECT 1429.750 16.760 1435.130 16.900 ;
        RECT 1429.750 16.700 1430.070 16.760 ;
        RECT 1434.810 16.700 1435.130 16.760 ;
      LAYER via ;
        RECT 1756.380 1329.780 1756.640 1330.040 ;
        RECT 1434.840 1313.120 1435.100 1313.380 ;
        RECT 1429.780 16.700 1430.040 16.960 ;
        RECT 1434.840 16.700 1435.100 16.960 ;
      LAYER met2 ;
        RECT 1756.370 1370.355 1756.650 1370.725 ;
        RECT 1756.440 1330.070 1756.580 1370.355 ;
        RECT 1756.380 1329.750 1756.640 1330.070 ;
        RECT 1434.840 1313.090 1435.100 1313.410 ;
        RECT 1434.900 16.990 1435.040 1313.090 ;
        RECT 1429.780 16.670 1430.040 16.990 ;
        RECT 1434.840 16.670 1435.100 16.990 ;
        RECT 1429.840 2.400 1429.980 16.670 ;
        RECT 1429.630 -4.800 1430.190 2.400 ;
      LAYER via2 ;
        RECT 1756.370 1370.400 1756.650 1370.680 ;
      LAYER met3 ;
        RECT 1755.835 1373.495 1759.835 1374.095 ;
        RECT 1756.590 1372.730 1756.890 1373.495 ;
        RECT 1756.590 1372.430 1757.120 1372.730 ;
        RECT 1756.820 1372.050 1757.120 1372.430 ;
        RECT 1756.820 1371.750 1757.810 1372.050 ;
        RECT 1756.345 1370.690 1756.675 1370.705 ;
        RECT 1757.510 1370.690 1757.810 1371.750 ;
        RECT 1756.345 1370.390 1757.810 1370.690 ;
        RECT 1756.345 1370.375 1756.675 1370.390 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1447.690 2.960 1448.010 3.020 ;
        RECT 1448.610 2.960 1448.930 3.020 ;
        RECT 1447.690 2.820 1448.930 2.960 ;
        RECT 1447.690 2.760 1448.010 2.820 ;
        RECT 1448.610 2.760 1448.930 2.820 ;
      LAYER via ;
        RECT 1447.720 2.760 1447.980 3.020 ;
        RECT 1448.640 2.760 1448.900 3.020 ;
      LAYER met2 ;
        RECT 1583.410 2392.395 1583.690 2392.765 ;
        RECT 1583.480 2377.880 1583.620 2392.395 ;
        RECT 1583.460 2373.880 1583.740 2377.880 ;
        RECT 1448.630 1326.155 1448.910 1326.525 ;
        RECT 1448.700 3.050 1448.840 1326.155 ;
        RECT 1447.720 2.730 1447.980 3.050 ;
        RECT 1448.640 2.730 1448.900 3.050 ;
        RECT 1447.780 2.400 1447.920 2.730 ;
        RECT 1447.570 -4.800 1448.130 2.400 ;
      LAYER via2 ;
        RECT 1583.410 2392.440 1583.690 2392.720 ;
        RECT 1448.630 1326.200 1448.910 1326.480 ;
      LAYER met3 ;
        RECT 1583.385 2392.730 1583.715 2392.745 ;
        RECT 1747.350 2392.730 1747.730 2392.740 ;
        RECT 1583.385 2392.430 1747.730 2392.730 ;
        RECT 1583.385 2392.415 1583.715 2392.430 ;
        RECT 1747.350 2392.420 1747.730 2392.430 ;
        RECT 1448.605 1326.490 1448.935 1326.505 ;
        RECT 1747.350 1326.490 1747.730 1326.500 ;
        RECT 1448.605 1326.190 1747.730 1326.490 ;
        RECT 1448.605 1326.175 1448.935 1326.190 ;
        RECT 1747.350 1326.180 1747.730 1326.190 ;
      LAYER via3 ;
        RECT 1747.380 2392.420 1747.700 2392.740 ;
        RECT 1747.380 1326.180 1747.700 1326.500 ;
      LAYER met4 ;
        RECT 1747.375 2392.415 1747.705 2392.745 ;
        RECT 1747.390 1326.505 1747.690 2392.415 ;
        RECT 1747.375 1326.175 1747.705 1326.505 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1469.385 1326.425 1469.555 1331.355 ;
      LAYER mcon ;
        RECT 1469.385 1331.185 1469.555 1331.355 ;
      LAYER met1 ;
        RECT 1469.325 1331.340 1469.615 1331.385 ;
        RECT 1761.410 1331.340 1761.730 1331.400 ;
        RECT 1469.325 1331.200 1761.730 1331.340 ;
        RECT 1469.325 1331.155 1469.615 1331.200 ;
        RECT 1761.410 1331.140 1761.730 1331.200 ;
        RECT 1469.310 1326.580 1469.630 1326.640 ;
        RECT 1469.115 1326.440 1469.630 1326.580 ;
        RECT 1469.310 1326.380 1469.630 1326.440 ;
        RECT 1465.630 15.200 1465.950 15.260 ;
        RECT 1469.310 15.200 1469.630 15.260 ;
        RECT 1465.630 15.060 1469.630 15.200 ;
        RECT 1465.630 15.000 1465.950 15.060 ;
        RECT 1469.310 15.000 1469.630 15.060 ;
      LAYER via ;
        RECT 1761.440 1331.140 1761.700 1331.400 ;
        RECT 1469.340 1326.380 1469.600 1326.640 ;
        RECT 1465.660 15.000 1465.920 15.260 ;
        RECT 1469.340 15.000 1469.600 15.260 ;
      LAYER met2 ;
        RECT 1761.430 2014.315 1761.710 2014.685 ;
        RECT 1761.500 1331.430 1761.640 2014.315 ;
        RECT 1761.440 1331.110 1761.700 1331.430 ;
        RECT 1469.340 1326.350 1469.600 1326.670 ;
        RECT 1469.400 15.290 1469.540 1326.350 ;
        RECT 1465.660 14.970 1465.920 15.290 ;
        RECT 1469.340 14.970 1469.600 15.290 ;
        RECT 1465.720 2.400 1465.860 14.970 ;
        RECT 1465.510 -4.800 1466.070 2.400 ;
      LAYER via2 ;
        RECT 1761.430 2014.360 1761.710 2014.640 ;
      LAYER met3 ;
        RECT 1755.835 2014.650 1759.835 2014.655 ;
        RECT 1761.405 2014.650 1761.735 2014.665 ;
        RECT 1755.835 2014.350 1761.735 2014.650 ;
        RECT 1755.835 2014.055 1759.835 2014.350 ;
        RECT 1761.405 2014.335 1761.735 2014.350 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1629.005 1325.745 1629.175 1327.955 ;
        RECT 1679.605 1325.745 1679.775 1327.955 ;
        RECT 1728.365 1327.785 1728.535 1328.975 ;
      LAYER mcon ;
        RECT 1728.365 1328.805 1728.535 1328.975 ;
        RECT 1629.005 1327.785 1629.175 1327.955 ;
        RECT 1679.605 1327.785 1679.775 1327.955 ;
      LAYER met1 ;
        RECT 1728.305 1328.960 1728.595 1329.005 ;
        RECT 1764.630 1328.960 1764.950 1329.020 ;
        RECT 1728.305 1328.820 1764.950 1328.960 ;
        RECT 1728.305 1328.775 1728.595 1328.820 ;
        RECT 1764.630 1328.760 1764.950 1328.820 ;
        RECT 1628.945 1327.940 1629.235 1327.985 ;
        RECT 1579.800 1327.800 1629.235 1327.940 ;
        RECT 1579.800 1327.600 1579.940 1327.800 ;
        RECT 1628.945 1327.755 1629.235 1327.800 ;
        RECT 1679.545 1327.940 1679.835 1327.985 ;
        RECT 1728.305 1327.940 1728.595 1327.985 ;
        RECT 1679.545 1327.800 1728.595 1327.940 ;
        RECT 1679.545 1327.755 1679.835 1327.800 ;
        RECT 1728.305 1327.755 1728.595 1327.800 ;
        RECT 1489.640 1327.460 1579.940 1327.600 ;
        RECT 1489.640 1326.640 1489.780 1327.460 ;
        RECT 1489.550 1326.380 1489.870 1326.640 ;
        RECT 1628.945 1325.900 1629.235 1325.945 ;
        RECT 1679.545 1325.900 1679.835 1325.945 ;
        RECT 1628.945 1325.760 1679.835 1325.900 ;
        RECT 1628.945 1325.715 1629.235 1325.760 ;
        RECT 1679.545 1325.715 1679.835 1325.760 ;
        RECT 1483.570 20.640 1483.890 20.700 ;
        RECT 1489.550 20.640 1489.870 20.700 ;
        RECT 1483.570 20.500 1489.870 20.640 ;
        RECT 1483.570 20.440 1483.890 20.500 ;
        RECT 1489.550 20.440 1489.870 20.500 ;
      LAYER via ;
        RECT 1764.660 1328.760 1764.920 1329.020 ;
        RECT 1489.580 1326.380 1489.840 1326.640 ;
        RECT 1483.600 20.440 1483.860 20.700 ;
        RECT 1489.580 20.440 1489.840 20.700 ;
      LAYER met2 ;
        RECT 1764.650 1647.115 1764.930 1647.485 ;
        RECT 1764.720 1329.050 1764.860 1647.115 ;
        RECT 1764.660 1328.730 1764.920 1329.050 ;
        RECT 1489.580 1326.350 1489.840 1326.670 ;
        RECT 1489.640 20.730 1489.780 1326.350 ;
        RECT 1483.600 20.410 1483.860 20.730 ;
        RECT 1489.580 20.410 1489.840 20.730 ;
        RECT 1483.660 2.400 1483.800 20.410 ;
        RECT 1483.450 -4.800 1484.010 2.400 ;
      LAYER via2 ;
        RECT 1764.650 1647.160 1764.930 1647.440 ;
      LAYER met3 ;
        RECT 1755.835 1647.450 1759.835 1647.455 ;
        RECT 1764.625 1647.450 1764.955 1647.465 ;
        RECT 1755.835 1647.150 1764.955 1647.450 ;
        RECT 1755.835 1646.855 1759.835 1647.150 ;
        RECT 1764.625 1647.135 1764.955 1647.150 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1265.090 2378.795 1265.370 2379.165 ;
        RECT 1265.160 2377.880 1265.300 2378.795 ;
        RECT 1265.140 2373.880 1265.420 2377.880 ;
        RECT 1501.530 15.795 1501.810 16.165 ;
        RECT 1501.600 2.400 1501.740 15.795 ;
        RECT 1501.390 -4.800 1501.950 2.400 ;
      LAYER via2 ;
        RECT 1265.090 2378.840 1265.370 2379.120 ;
        RECT 1501.530 15.840 1501.810 16.120 ;
      LAYER met3 ;
        RECT 1265.065 2379.130 1265.395 2379.145 ;
        RECT 1743.670 2379.130 1744.050 2379.140 ;
        RECT 1265.065 2378.830 1744.050 2379.130 ;
        RECT 1265.065 2378.815 1265.395 2378.830 ;
        RECT 1743.670 2378.820 1744.050 2378.830 ;
        RECT 1501.505 16.130 1501.835 16.145 ;
        RECT 1743.670 16.130 1744.050 16.140 ;
        RECT 1501.505 15.830 1744.050 16.130 ;
        RECT 1501.505 15.815 1501.835 15.830 ;
        RECT 1743.670 15.820 1744.050 15.830 ;
      LAYER via3 ;
        RECT 1743.700 2378.820 1744.020 2379.140 ;
        RECT 1743.700 15.820 1744.020 16.140 ;
      LAYER met4 ;
        RECT 1743.695 2378.815 1744.025 2379.145 ;
        RECT 1743.710 16.145 1744.010 2378.815 ;
        RECT 1743.695 15.815 1744.025 16.145 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1334.090 2393.755 1334.370 2394.125 ;
        RECT 1334.160 2377.880 1334.300 2393.755 ;
        RECT 1334.140 2373.880 1334.420 2377.880 ;
        RECT 1519.010 15.115 1519.290 15.485 ;
        RECT 1519.080 2.400 1519.220 15.115 ;
        RECT 1518.870 -4.800 1519.430 2.400 ;
      LAYER via2 ;
        RECT 1334.090 2393.800 1334.370 2394.080 ;
        RECT 1519.010 15.160 1519.290 15.440 ;
      LAYER met3 ;
        RECT 1334.065 2394.090 1334.395 2394.105 ;
        RECT 1763.910 2394.090 1764.290 2394.100 ;
        RECT 1334.065 2393.790 1764.290 2394.090 ;
        RECT 1334.065 2393.775 1334.395 2393.790 ;
        RECT 1763.910 2393.780 1764.290 2393.790 ;
        RECT 1763.910 1498.900 1764.290 1499.220 ;
        RECT 1763.950 1498.530 1764.250 1498.900 ;
        RECT 1764.830 1498.530 1765.210 1498.540 ;
        RECT 1763.950 1498.230 1765.210 1498.530 ;
        RECT 1764.830 1498.220 1765.210 1498.230 ;
        RECT 1518.985 15.450 1519.315 15.465 ;
        RECT 1751.030 15.450 1751.410 15.460 ;
        RECT 1518.985 15.150 1751.410 15.450 ;
        RECT 1518.985 15.135 1519.315 15.150 ;
        RECT 1751.030 15.140 1751.410 15.150 ;
      LAYER via3 ;
        RECT 1763.940 2393.780 1764.260 2394.100 ;
        RECT 1763.940 1498.900 1764.260 1499.220 ;
        RECT 1764.860 1498.220 1765.180 1498.540 ;
        RECT 1751.060 15.140 1751.380 15.460 ;
      LAYER met4 ;
        RECT 1763.935 2393.775 1764.265 2394.105 ;
        RECT 1763.950 1499.225 1764.250 2393.775 ;
        RECT 1763.935 1498.895 1764.265 1499.225 ;
        RECT 1764.855 1498.215 1765.185 1498.545 ;
        RECT 1764.870 1494.890 1765.170 1498.215 ;
        RECT 1750.630 1493.710 1751.810 1494.890 ;
        RECT 1764.430 1493.710 1765.610 1494.890 ;
        RECT 1751.070 15.465 1751.370 1493.710 ;
        RECT 1751.055 15.135 1751.385 15.465 ;
      LAYER met5 ;
        RECT 1750.420 1493.500 1765.820 1495.100 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 687.770 2376.160 688.090 2376.220 ;
        RECT 1101.310 2376.160 1101.630 2376.220 ;
        RECT 687.770 2376.020 1101.630 2376.160 ;
        RECT 687.770 2375.960 688.090 2376.020 ;
        RECT 1101.310 2375.960 1101.630 2376.020 ;
        RECT 687.770 1324.200 688.090 1324.260 ;
        RECT 712.610 1324.200 712.930 1324.260 ;
        RECT 687.770 1324.060 712.930 1324.200 ;
        RECT 687.770 1324.000 688.090 1324.060 ;
        RECT 712.610 1324.000 712.930 1324.060 ;
        RECT 712.610 20.640 712.930 20.700 ;
        RECT 716.290 20.640 716.610 20.700 ;
        RECT 712.610 20.500 716.610 20.640 ;
        RECT 712.610 20.440 712.930 20.500 ;
        RECT 716.290 20.440 716.610 20.500 ;
      LAYER via ;
        RECT 687.800 2375.960 688.060 2376.220 ;
        RECT 1101.340 2375.960 1101.600 2376.220 ;
        RECT 687.800 1324.000 688.060 1324.260 ;
        RECT 712.640 1324.000 712.900 1324.260 ;
        RECT 712.640 20.440 712.900 20.700 ;
        RECT 716.320 20.440 716.580 20.700 ;
      LAYER met2 ;
        RECT 1103.220 2376.330 1103.500 2377.880 ;
        RECT 1101.400 2376.250 1103.500 2376.330 ;
        RECT 687.800 2375.930 688.060 2376.250 ;
        RECT 1101.340 2376.190 1103.500 2376.250 ;
        RECT 1101.340 2375.930 1101.600 2376.190 ;
        RECT 687.860 1324.290 688.000 2375.930 ;
        RECT 1103.220 2373.880 1103.500 2376.190 ;
        RECT 687.800 1323.970 688.060 1324.290 ;
        RECT 712.640 1323.970 712.900 1324.290 ;
        RECT 712.700 20.730 712.840 1323.970 ;
        RECT 712.640 20.410 712.900 20.730 ;
        RECT 716.320 20.410 716.580 20.730 ;
        RECT 716.380 2.400 716.520 20.410 ;
        RECT 716.170 -4.800 716.730 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1629.465 1327.445 1629.635 1328.975 ;
        RECT 1680.065 1327.445 1680.235 1328.975 ;
        RECT 1704.445 1325.405 1704.615 1327.615 ;
        RECT 1752.285 1325.745 1752.455 1327.955 ;
      LAYER mcon ;
        RECT 1629.465 1328.805 1629.635 1328.975 ;
        RECT 1680.065 1328.805 1680.235 1328.975 ;
        RECT 1752.285 1327.785 1752.455 1327.955 ;
        RECT 1704.445 1327.445 1704.615 1327.615 ;
      LAYER met1 ;
        RECT 1560.390 2394.180 1560.710 2394.240 ;
        RECT 1784.870 2394.180 1785.190 2394.240 ;
        RECT 1560.390 2394.040 1785.190 2394.180 ;
        RECT 1560.390 2393.980 1560.710 2394.040 ;
        RECT 1784.870 2393.980 1785.190 2394.040 ;
        RECT 1629.405 1328.960 1629.695 1329.005 ;
        RECT 1680.005 1328.960 1680.295 1329.005 ;
        RECT 1629.405 1328.820 1680.295 1328.960 ;
        RECT 1629.405 1328.775 1629.695 1328.820 ;
        RECT 1680.005 1328.775 1680.295 1328.820 ;
        RECT 1752.225 1327.940 1752.515 1327.985 ;
        RECT 1784.870 1327.940 1785.190 1328.000 ;
        RECT 1752.225 1327.800 1785.190 1327.940 ;
        RECT 1752.225 1327.755 1752.515 1327.800 ;
        RECT 1784.870 1327.740 1785.190 1327.800 ;
        RECT 1629.405 1327.600 1629.695 1327.645 ;
        RECT 1604.180 1327.460 1629.695 1327.600 ;
        RECT 1604.180 1327.260 1604.320 1327.460 ;
        RECT 1629.405 1327.415 1629.695 1327.460 ;
        RECT 1680.005 1327.600 1680.295 1327.645 ;
        RECT 1704.385 1327.600 1704.675 1327.645 ;
        RECT 1680.005 1327.460 1704.675 1327.600 ;
        RECT 1680.005 1327.415 1680.295 1327.460 ;
        RECT 1704.385 1327.415 1704.675 1327.460 ;
        RECT 1579.800 1327.120 1604.320 1327.260 ;
        RECT 1538.310 1326.240 1538.630 1326.300 ;
        RECT 1579.800 1326.240 1579.940 1327.120 ;
        RECT 1538.310 1326.100 1579.940 1326.240 ;
        RECT 1538.310 1326.040 1538.630 1326.100 ;
        RECT 1752.225 1325.900 1752.515 1325.945 ;
        RECT 1750.000 1325.760 1752.515 1325.900 ;
        RECT 1704.385 1325.560 1704.675 1325.605 ;
        RECT 1750.000 1325.560 1750.140 1325.760 ;
        RECT 1752.225 1325.715 1752.515 1325.760 ;
        RECT 1704.385 1325.420 1750.140 1325.560 ;
        RECT 1704.385 1325.375 1704.675 1325.420 ;
      LAYER via ;
        RECT 1560.420 2393.980 1560.680 2394.240 ;
        RECT 1784.900 2393.980 1785.160 2394.240 ;
        RECT 1784.900 1327.740 1785.160 1328.000 ;
        RECT 1538.340 1326.040 1538.600 1326.300 ;
      LAYER met2 ;
        RECT 1560.420 2393.950 1560.680 2394.270 ;
        RECT 1784.900 2393.950 1785.160 2394.270 ;
        RECT 1560.480 2377.880 1560.620 2393.950 ;
        RECT 1560.460 2373.880 1560.740 2377.880 ;
        RECT 1784.960 1328.030 1785.100 2393.950 ;
        RECT 1784.900 1327.710 1785.160 1328.030 ;
        RECT 1538.340 1326.010 1538.600 1326.330 ;
        RECT 1538.400 7.210 1538.540 1326.010 ;
        RECT 1537.020 7.070 1538.540 7.210 ;
        RECT 1537.020 2.400 1537.160 7.070 ;
        RECT 1536.810 -4.800 1537.370 2.400 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1197.910 1312.640 1198.230 1312.700 ;
        RECT 1552.570 1312.640 1552.890 1312.700 ;
        RECT 1197.910 1312.500 1552.890 1312.640 ;
        RECT 1197.910 1312.440 1198.230 1312.500 ;
        RECT 1552.570 1312.440 1552.890 1312.500 ;
      LAYER via ;
        RECT 1197.940 1312.440 1198.200 1312.700 ;
        RECT 1552.600 1312.440 1552.860 1312.700 ;
      LAYER met2 ;
        RECT 1197.980 1323.135 1198.260 1327.135 ;
        RECT 1198.000 1312.730 1198.140 1323.135 ;
        RECT 1197.940 1312.410 1198.200 1312.730 ;
        RECT 1552.600 1312.410 1552.860 1312.730 ;
        RECT 1552.660 7.210 1552.800 1312.410 ;
        RECT 1552.660 7.070 1555.100 7.210 ;
        RECT 1554.960 2.400 1555.100 7.070 ;
        RECT 1554.750 -4.800 1555.310 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1607.385 1311.805 1608.015 1311.975 ;
        RECT 1690.645 1311.465 1690.815 1312.315 ;
        RECT 1703.985 1311.975 1704.155 1312.315 ;
        RECT 1703.985 1311.805 1704.615 1311.975 ;
        RECT 1571.965 48.365 1572.135 62.475 ;
      LAYER mcon ;
        RECT 1690.645 1312.145 1690.815 1312.315 ;
        RECT 1607.845 1311.805 1608.015 1311.975 ;
        RECT 1703.985 1312.145 1704.155 1312.315 ;
        RECT 1704.445 1311.805 1704.615 1311.975 ;
        RECT 1571.965 62.305 1572.135 62.475 ;
      LAYER met1 ;
        RECT 1763.250 1345.620 1763.570 1345.680 ;
        RECT 1764.170 1345.620 1764.490 1345.680 ;
        RECT 1763.250 1345.480 1764.490 1345.620 ;
        RECT 1763.250 1345.420 1763.570 1345.480 ;
        RECT 1764.170 1345.420 1764.490 1345.480 ;
        RECT 1690.585 1312.300 1690.875 1312.345 ;
        RECT 1703.925 1312.300 1704.215 1312.345 ;
        RECT 1763.250 1312.300 1763.570 1312.360 ;
        RECT 1690.585 1312.160 1704.215 1312.300 ;
        RECT 1690.585 1312.115 1690.875 1312.160 ;
        RECT 1703.925 1312.115 1704.215 1312.160 ;
        RECT 1738.500 1312.160 1763.570 1312.300 ;
        RECT 1572.350 1311.960 1572.670 1312.020 ;
        RECT 1607.325 1311.960 1607.615 1312.005 ;
        RECT 1572.350 1311.820 1607.615 1311.960 ;
        RECT 1572.350 1311.760 1572.670 1311.820 ;
        RECT 1607.325 1311.775 1607.615 1311.820 ;
        RECT 1607.785 1311.960 1608.075 1312.005 ;
        RECT 1704.385 1311.960 1704.675 1312.005 ;
        RECT 1738.500 1311.960 1738.640 1312.160 ;
        RECT 1763.250 1312.100 1763.570 1312.160 ;
        RECT 1607.785 1311.820 1642.960 1311.960 ;
        RECT 1607.785 1311.775 1608.075 1311.820 ;
        RECT 1642.820 1311.620 1642.960 1311.820 ;
        RECT 1704.385 1311.820 1738.640 1311.960 ;
        RECT 1704.385 1311.775 1704.675 1311.820 ;
        RECT 1690.585 1311.620 1690.875 1311.665 ;
        RECT 1642.820 1311.480 1690.875 1311.620 ;
        RECT 1690.585 1311.435 1690.875 1311.480 ;
        RECT 1571.905 62.460 1572.195 62.505 ;
        RECT 1572.350 62.460 1572.670 62.520 ;
        RECT 1571.905 62.320 1572.670 62.460 ;
        RECT 1571.905 62.275 1572.195 62.320 ;
        RECT 1572.350 62.260 1572.670 62.320 ;
        RECT 1571.890 48.520 1572.210 48.580 ;
        RECT 1571.695 48.380 1572.210 48.520 ;
        RECT 1571.890 48.320 1572.210 48.380 ;
      LAYER via ;
        RECT 1763.280 1345.420 1763.540 1345.680 ;
        RECT 1764.200 1345.420 1764.460 1345.680 ;
        RECT 1572.380 1311.760 1572.640 1312.020 ;
        RECT 1763.280 1312.100 1763.540 1312.360 ;
        RECT 1572.380 62.260 1572.640 62.520 ;
        RECT 1571.920 48.320 1572.180 48.580 ;
      LAYER met2 ;
        RECT 1764.190 1954.475 1764.470 1954.845 ;
        RECT 1764.260 1345.710 1764.400 1954.475 ;
        RECT 1763.280 1345.390 1763.540 1345.710 ;
        RECT 1764.200 1345.390 1764.460 1345.710 ;
        RECT 1763.340 1312.390 1763.480 1345.390 ;
        RECT 1763.280 1312.070 1763.540 1312.390 ;
        RECT 1572.380 1311.730 1572.640 1312.050 ;
        RECT 1572.440 62.550 1572.580 1311.730 ;
        RECT 1572.380 62.230 1572.640 62.550 ;
        RECT 1571.920 48.290 1572.180 48.610 ;
        RECT 1571.980 17.410 1572.120 48.290 ;
        RECT 1571.980 17.270 1573.040 17.410 ;
        RECT 1572.900 2.400 1573.040 17.270 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
      LAYER via2 ;
        RECT 1764.190 1954.520 1764.470 1954.800 ;
      LAYER met3 ;
        RECT 1755.835 1954.810 1759.835 1954.815 ;
        RECT 1764.165 1954.810 1764.495 1954.825 ;
        RECT 1755.835 1954.510 1764.495 1954.810 ;
        RECT 1755.835 1954.215 1759.835 1954.510 ;
        RECT 1764.165 1954.495 1764.495 1954.510 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1754.585 1326.085 1754.755 1368.415 ;
      LAYER mcon ;
        RECT 1754.585 1368.245 1754.755 1368.415 ;
      LAYER met1 ;
        RECT 1754.525 1368.400 1754.815 1368.445 ;
        RECT 1756.810 1368.400 1757.130 1368.460 ;
        RECT 1754.525 1368.260 1757.130 1368.400 ;
        RECT 1754.525 1368.215 1754.815 1368.260 ;
        RECT 1756.810 1368.200 1757.130 1368.260 ;
        RECT 1751.750 1326.240 1752.070 1326.300 ;
        RECT 1754.525 1326.240 1754.815 1326.285 ;
        RECT 1751.750 1326.100 1754.815 1326.240 ;
        RECT 1751.750 1326.040 1752.070 1326.100 ;
        RECT 1754.525 1326.055 1754.815 1326.100 ;
      LAYER via ;
        RECT 1756.840 1368.200 1757.100 1368.460 ;
        RECT 1751.780 1326.040 1752.040 1326.300 ;
      LAYER met2 ;
        RECT 923.770 2393.755 924.050 2394.125 ;
        RECT 976.210 2393.755 976.490 2394.125 ;
        RECT 923.840 2377.880 923.980 2393.755 ;
        RECT 976.280 2392.085 976.420 2393.755 ;
        RECT 976.210 2391.715 976.490 2392.085 ;
        RECT 923.820 2373.880 924.100 2377.880 ;
        RECT 1759.130 2342.075 1759.410 2342.445 ;
        RECT 1759.200 2319.325 1759.340 2342.075 ;
        RECT 1759.130 2318.955 1759.410 2319.325 ;
        RECT 1757.750 2148.955 1758.030 2149.325 ;
        RECT 1757.820 2077.245 1757.960 2148.955 ;
        RECT 1757.750 2076.875 1758.030 2077.245 ;
        RECT 1757.750 2076.195 1758.030 2076.565 ;
        RECT 1757.820 2011.285 1757.960 2076.195 ;
        RECT 1757.750 2010.915 1758.030 2011.285 ;
        RECT 1759.130 1848.395 1759.410 1848.765 ;
        RECT 1759.200 1789.605 1759.340 1848.395 ;
        RECT 1759.130 1789.235 1759.410 1789.605 ;
        RECT 1759.130 1728.715 1759.410 1729.085 ;
        RECT 1759.200 1723.645 1759.340 1728.715 ;
        RECT 1759.130 1723.275 1759.410 1723.645 ;
        RECT 1756.830 1368.995 1757.110 1369.365 ;
        RECT 1756.900 1368.490 1757.040 1368.995 ;
        RECT 1756.840 1368.170 1757.100 1368.490 ;
        RECT 1751.780 1326.010 1752.040 1326.330 ;
        RECT 1751.840 1325.845 1751.980 1326.010 ;
        RECT 1751.770 1325.475 1752.050 1325.845 ;
        RECT 1590.310 14.435 1590.590 14.805 ;
        RECT 1590.380 2.400 1590.520 14.435 ;
        RECT 1590.170 -4.800 1590.730 2.400 ;
      LAYER via2 ;
        RECT 923.770 2393.800 924.050 2394.080 ;
        RECT 976.210 2393.800 976.490 2394.080 ;
        RECT 976.210 2391.760 976.490 2392.040 ;
        RECT 1759.130 2342.120 1759.410 2342.400 ;
        RECT 1759.130 2319.000 1759.410 2319.280 ;
        RECT 1757.750 2149.000 1758.030 2149.280 ;
        RECT 1757.750 2076.920 1758.030 2077.200 ;
        RECT 1757.750 2076.240 1758.030 2076.520 ;
        RECT 1757.750 2010.960 1758.030 2011.240 ;
        RECT 1759.130 1848.440 1759.410 1848.720 ;
        RECT 1759.130 1789.280 1759.410 1789.560 ;
        RECT 1759.130 1728.760 1759.410 1729.040 ;
        RECT 1759.130 1723.320 1759.410 1723.600 ;
        RECT 1756.830 1369.040 1757.110 1369.320 ;
        RECT 1751.770 1325.520 1752.050 1325.800 ;
        RECT 1590.310 14.480 1590.590 14.760 ;
      LAYER met3 ;
        RECT 923.745 2394.090 924.075 2394.105 ;
        RECT 976.185 2394.090 976.515 2394.105 ;
        RECT 923.745 2393.790 976.515 2394.090 ;
        RECT 923.745 2393.775 924.075 2393.790 ;
        RECT 976.185 2393.775 976.515 2393.790 ;
        RECT 976.185 2392.050 976.515 2392.065 ;
        RECT 1756.550 2392.050 1756.930 2392.060 ;
        RECT 976.185 2391.750 1756.930 2392.050 ;
        RECT 976.185 2391.735 976.515 2391.750 ;
        RECT 1756.550 2391.740 1756.930 2391.750 ;
        RECT 1756.550 2342.410 1756.930 2342.420 ;
        RECT 1759.105 2342.410 1759.435 2342.425 ;
        RECT 1756.550 2342.110 1759.435 2342.410 ;
        RECT 1756.550 2342.100 1756.930 2342.110 ;
        RECT 1759.105 2342.095 1759.435 2342.110 ;
        RECT 1757.470 2319.290 1757.850 2319.300 ;
        RECT 1759.105 2319.290 1759.435 2319.305 ;
        RECT 1757.470 2318.990 1759.435 2319.290 ;
        RECT 1757.470 2318.980 1757.850 2318.990 ;
        RECT 1759.105 2318.975 1759.435 2318.990 ;
        RECT 1758.390 2260.130 1758.770 2260.140 ;
        RECT 1757.510 2259.830 1758.770 2260.130 ;
        RECT 1757.510 2258.780 1757.810 2259.830 ;
        RECT 1758.390 2259.820 1758.770 2259.830 ;
        RECT 1757.470 2258.460 1757.850 2258.780 ;
        RECT 1757.725 2149.300 1758.055 2149.305 ;
        RECT 1757.470 2149.290 1758.055 2149.300 ;
        RECT 1757.270 2148.990 1758.055 2149.290 ;
        RECT 1757.470 2148.980 1758.055 2148.990 ;
        RECT 1757.725 2148.975 1758.055 2148.980 ;
        RECT 1757.725 2077.220 1758.055 2077.225 ;
        RECT 1757.470 2077.210 1758.055 2077.220 ;
        RECT 1757.270 2076.910 1758.055 2077.210 ;
        RECT 1757.470 2076.900 1758.055 2076.910 ;
        RECT 1757.725 2076.895 1758.055 2076.900 ;
        RECT 1757.725 2076.540 1758.055 2076.545 ;
        RECT 1757.470 2076.530 1758.055 2076.540 ;
        RECT 1757.470 2076.230 1758.280 2076.530 ;
        RECT 1757.470 2076.220 1758.055 2076.230 ;
        RECT 1757.725 2076.215 1758.055 2076.220 ;
        RECT 1756.550 2011.250 1756.930 2011.260 ;
        RECT 1757.725 2011.250 1758.055 2011.265 ;
        RECT 1756.550 2010.950 1758.055 2011.250 ;
        RECT 1756.550 2010.940 1756.930 2010.950 ;
        RECT 1757.725 2010.935 1758.055 2010.950 ;
        RECT 1758.390 1848.730 1758.770 1848.740 ;
        RECT 1759.105 1848.730 1759.435 1848.745 ;
        RECT 1758.390 1848.430 1759.435 1848.730 ;
        RECT 1758.390 1848.420 1758.770 1848.430 ;
        RECT 1759.105 1848.415 1759.435 1848.430 ;
        RECT 1756.550 1789.570 1756.930 1789.580 ;
        RECT 1759.105 1789.570 1759.435 1789.585 ;
        RECT 1756.550 1789.270 1759.435 1789.570 ;
        RECT 1756.550 1789.260 1756.930 1789.270 ;
        RECT 1759.105 1789.255 1759.435 1789.270 ;
        RECT 1756.550 1770.530 1756.930 1770.540 ;
        RECT 1758.390 1770.530 1758.770 1770.540 ;
        RECT 1756.550 1770.230 1758.770 1770.530 ;
        RECT 1756.550 1770.220 1756.930 1770.230 ;
        RECT 1758.390 1770.220 1758.770 1770.230 ;
        RECT 1758.390 1729.050 1758.770 1729.060 ;
        RECT 1759.105 1729.050 1759.435 1729.065 ;
        RECT 1758.390 1728.750 1759.435 1729.050 ;
        RECT 1758.390 1728.740 1758.770 1728.750 ;
        RECT 1759.105 1728.735 1759.435 1728.750 ;
        RECT 1756.550 1723.610 1756.930 1723.620 ;
        RECT 1759.105 1723.610 1759.435 1723.625 ;
        RECT 1756.550 1723.310 1759.435 1723.610 ;
        RECT 1756.550 1723.300 1756.930 1723.310 ;
        RECT 1759.105 1723.295 1759.435 1723.310 ;
        RECT 1757.470 1607.700 1757.850 1608.020 ;
        RECT 1757.510 1605.980 1757.810 1607.700 ;
        RECT 1757.470 1605.660 1757.850 1605.980 ;
        RECT 1757.470 1556.020 1757.850 1556.340 ;
        RECT 1757.510 1554.980 1757.810 1556.020 ;
        RECT 1757.470 1554.660 1757.850 1554.980 ;
        RECT 1757.470 1539.020 1757.850 1539.340 ;
        RECT 1757.510 1537.980 1757.810 1539.020 ;
        RECT 1757.470 1537.660 1757.850 1537.980 ;
        RECT 1756.805 1369.340 1757.135 1369.345 ;
        RECT 1756.550 1369.330 1757.135 1369.340 ;
        RECT 1756.550 1369.030 1757.360 1369.330 ;
        RECT 1756.550 1369.020 1757.135 1369.030 ;
        RECT 1756.805 1369.015 1757.135 1369.020 ;
        RECT 1751.745 1325.810 1752.075 1325.825 ;
        RECT 1751.745 1325.495 1752.290 1325.810 ;
        RECT 1751.990 1325.140 1752.290 1325.495 ;
        RECT 1751.950 1324.820 1752.330 1325.140 ;
        RECT 1590.285 14.770 1590.615 14.785 ;
        RECT 1751.950 14.770 1752.330 14.780 ;
        RECT 1590.285 14.470 1752.330 14.770 ;
        RECT 1590.285 14.455 1590.615 14.470 ;
        RECT 1751.950 14.460 1752.330 14.470 ;
      LAYER via3 ;
        RECT 1756.580 2391.740 1756.900 2392.060 ;
        RECT 1756.580 2342.100 1756.900 2342.420 ;
        RECT 1757.500 2318.980 1757.820 2319.300 ;
        RECT 1758.420 2259.820 1758.740 2260.140 ;
        RECT 1757.500 2258.460 1757.820 2258.780 ;
        RECT 1757.500 2148.980 1757.820 2149.300 ;
        RECT 1757.500 2076.900 1757.820 2077.220 ;
        RECT 1757.500 2076.220 1757.820 2076.540 ;
        RECT 1756.580 2010.940 1756.900 2011.260 ;
        RECT 1758.420 1848.420 1758.740 1848.740 ;
        RECT 1756.580 1789.260 1756.900 1789.580 ;
        RECT 1756.580 1770.220 1756.900 1770.540 ;
        RECT 1758.420 1770.220 1758.740 1770.540 ;
        RECT 1758.420 1728.740 1758.740 1729.060 ;
        RECT 1756.580 1723.300 1756.900 1723.620 ;
        RECT 1757.500 1607.700 1757.820 1608.020 ;
        RECT 1757.500 1605.660 1757.820 1605.980 ;
        RECT 1757.500 1556.020 1757.820 1556.340 ;
        RECT 1757.500 1554.660 1757.820 1554.980 ;
        RECT 1757.500 1539.020 1757.820 1539.340 ;
        RECT 1757.500 1537.660 1757.820 1537.980 ;
        RECT 1756.580 1369.020 1756.900 1369.340 ;
        RECT 1751.980 1324.820 1752.300 1325.140 ;
        RECT 1751.980 14.460 1752.300 14.780 ;
      LAYER met4 ;
        RECT 1756.575 2391.735 1756.905 2392.065 ;
        RECT 1756.590 2342.425 1756.890 2391.735 ;
        RECT 1756.575 2342.095 1756.905 2342.425 ;
        RECT 1757.495 2318.975 1757.825 2319.305 ;
        RECT 1757.510 2307.050 1757.810 2318.975 ;
        RECT 1757.510 2306.750 1759.650 2307.050 ;
        RECT 1759.350 2293.450 1759.650 2306.750 ;
        RECT 1758.430 2293.150 1759.650 2293.450 ;
        RECT 1758.430 2260.145 1758.730 2293.150 ;
        RECT 1758.415 2259.815 1758.745 2260.145 ;
        RECT 1757.495 2258.455 1757.825 2258.785 ;
        RECT 1757.510 2149.305 1757.810 2258.455 ;
        RECT 1757.495 2148.975 1757.825 2149.305 ;
        RECT 1757.495 2076.895 1757.825 2077.225 ;
        RECT 1757.510 2076.545 1757.810 2076.895 ;
        RECT 1757.495 2076.215 1757.825 2076.545 ;
        RECT 1756.575 2011.250 1756.905 2011.265 ;
        RECT 1754.750 2010.950 1756.905 2011.250 ;
        RECT 1754.750 2007.850 1755.050 2010.950 ;
        RECT 1756.575 2010.935 1756.905 2010.950 ;
        RECT 1752.910 2007.550 1755.050 2007.850 ;
        RECT 1752.910 1956.850 1753.210 2007.550 ;
        RECT 1752.910 1956.550 1756.890 1956.850 ;
        RECT 1756.590 1950.050 1756.890 1956.550 ;
        RECT 1756.590 1949.750 1758.730 1950.050 ;
        RECT 1758.430 1848.745 1758.730 1949.750 ;
        RECT 1758.415 1848.415 1758.745 1848.745 ;
        RECT 1756.575 1789.255 1756.905 1789.585 ;
        RECT 1756.590 1770.545 1756.890 1789.255 ;
        RECT 1756.575 1770.215 1756.905 1770.545 ;
        RECT 1758.415 1770.215 1758.745 1770.545 ;
        RECT 1758.430 1729.065 1758.730 1770.215 ;
        RECT 1758.415 1728.735 1758.745 1729.065 ;
        RECT 1756.575 1723.295 1756.905 1723.625 ;
        RECT 1756.590 1722.250 1756.890 1723.295 ;
        RECT 1755.670 1721.950 1756.890 1722.250 ;
        RECT 1755.670 1664.450 1755.970 1721.950 ;
        RECT 1755.670 1664.150 1757.810 1664.450 ;
        RECT 1757.510 1608.025 1757.810 1664.150 ;
        RECT 1757.495 1607.695 1757.825 1608.025 ;
        RECT 1757.495 1605.655 1757.825 1605.985 ;
        RECT 1757.510 1556.345 1757.810 1605.655 ;
        RECT 1757.495 1556.015 1757.825 1556.345 ;
        RECT 1757.495 1554.655 1757.825 1554.985 ;
        RECT 1757.510 1539.345 1757.810 1554.655 ;
        RECT 1757.495 1539.015 1757.825 1539.345 ;
        RECT 1757.495 1537.655 1757.825 1537.985 ;
        RECT 1757.510 1404.010 1757.810 1537.655 ;
        RECT 1756.590 1403.710 1757.810 1404.010 ;
        RECT 1756.590 1369.345 1756.890 1403.710 ;
        RECT 1756.575 1369.015 1756.905 1369.345 ;
        RECT 1751.975 1324.815 1752.305 1325.145 ;
        RECT 1751.990 14.785 1752.290 1324.815 ;
        RECT 1751.975 14.455 1752.305 14.785 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1710.350 2390.780 1710.670 2390.840 ;
        RECT 1782.570 2390.780 1782.890 2390.840 ;
        RECT 1710.350 2390.640 1782.890 2390.780 ;
        RECT 1710.350 2390.580 1710.670 2390.640 ;
        RECT 1782.570 2390.580 1782.890 2390.640 ;
        RECT 1782.570 1326.920 1782.890 1326.980 ;
        RECT 1614.300 1326.780 1782.890 1326.920 ;
        RECT 1614.300 1326.640 1614.440 1326.780 ;
        RECT 1782.570 1326.720 1782.890 1326.780 ;
        RECT 1614.210 1326.380 1614.530 1326.640 ;
        RECT 1608.230 20.640 1608.550 20.700 ;
        RECT 1614.210 20.640 1614.530 20.700 ;
        RECT 1608.230 20.500 1614.530 20.640 ;
        RECT 1608.230 20.440 1608.550 20.500 ;
        RECT 1614.210 20.440 1614.530 20.500 ;
      LAYER via ;
        RECT 1710.380 2390.580 1710.640 2390.840 ;
        RECT 1782.600 2390.580 1782.860 2390.840 ;
        RECT 1782.600 1326.720 1782.860 1326.980 ;
        RECT 1614.240 1326.380 1614.500 1326.640 ;
        RECT 1608.260 20.440 1608.520 20.700 ;
        RECT 1614.240 20.440 1614.500 20.700 ;
      LAYER met2 ;
        RECT 1710.380 2390.550 1710.640 2390.870 ;
        RECT 1782.600 2390.550 1782.860 2390.870 ;
        RECT 1710.440 2377.880 1710.580 2390.550 ;
        RECT 1710.420 2373.880 1710.700 2377.880 ;
        RECT 1782.660 1327.010 1782.800 2390.550 ;
        RECT 1782.600 1326.690 1782.860 1327.010 ;
        RECT 1614.240 1326.350 1614.500 1326.670 ;
        RECT 1614.300 20.730 1614.440 1326.350 ;
        RECT 1608.260 20.410 1608.520 20.730 ;
        RECT 1614.240 20.410 1614.500 20.730 ;
        RECT 1608.320 2.400 1608.460 20.410 ;
        RECT 1608.110 -4.800 1608.670 2.400 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 951.885 2388.925 952.055 2394.535 ;
      LAYER mcon ;
        RECT 951.885 2394.365 952.055 2394.535 ;
      LAYER met1 ;
        RECT 951.825 2394.520 952.115 2394.565 ;
        RECT 951.825 2394.380 952.500 2394.520 ;
        RECT 951.825 2394.335 952.115 2394.380 ;
        RECT 952.360 2394.180 952.500 2394.380 ;
        RECT 952.360 2394.040 952.960 2394.180 ;
        RECT 952.820 2393.840 952.960 2394.040 ;
        RECT 1773.830 2393.840 1774.150 2393.900 ;
        RECT 952.820 2393.700 1774.150 2393.840 ;
        RECT 1773.830 2393.640 1774.150 2393.700 ;
        RECT 906.270 2389.080 906.590 2389.140 ;
        RECT 951.825 2389.080 952.115 2389.125 ;
        RECT 906.270 2388.940 952.115 2389.080 ;
        RECT 906.270 2388.880 906.590 2388.940 ;
        RECT 951.825 2388.895 952.115 2388.940 ;
        RECT 1626.170 16.220 1626.490 16.280 ;
        RECT 1773.830 16.220 1774.150 16.280 ;
        RECT 1626.170 16.080 1774.150 16.220 ;
        RECT 1626.170 16.020 1626.490 16.080 ;
        RECT 1773.830 16.020 1774.150 16.080 ;
      LAYER via ;
        RECT 1773.860 2393.640 1774.120 2393.900 ;
        RECT 906.300 2388.880 906.560 2389.140 ;
        RECT 1626.200 16.020 1626.460 16.280 ;
        RECT 1773.860 16.020 1774.120 16.280 ;
      LAYER met2 ;
        RECT 1773.860 2393.610 1774.120 2393.930 ;
        RECT 906.300 2388.850 906.560 2389.170 ;
        RECT 906.360 2377.880 906.500 2388.850 ;
        RECT 906.340 2373.880 906.620 2377.880 ;
        RECT 1773.920 16.310 1774.060 2393.610 ;
        RECT 1626.200 15.990 1626.460 16.310 ;
        RECT 1773.860 15.990 1774.120 16.310 ;
        RECT 1626.260 2.400 1626.400 15.990 ;
        RECT 1626.050 -4.800 1626.610 2.400 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1467.470 2392.820 1467.790 2392.880 ;
        RECT 1787.170 2392.820 1787.490 2392.880 ;
        RECT 1467.470 2392.680 1787.490 2392.820 ;
        RECT 1467.470 2392.620 1467.790 2392.680 ;
        RECT 1787.170 2392.620 1787.490 2392.680 ;
        RECT 1787.170 15.540 1787.490 15.600 ;
        RECT 1664.900 15.400 1787.490 15.540 ;
        RECT 1644.110 15.200 1644.430 15.260 ;
        RECT 1664.900 15.200 1665.040 15.400 ;
        RECT 1787.170 15.340 1787.490 15.400 ;
        RECT 1644.110 15.060 1665.040 15.200 ;
        RECT 1644.110 15.000 1644.430 15.060 ;
      LAYER via ;
        RECT 1467.500 2392.620 1467.760 2392.880 ;
        RECT 1787.200 2392.620 1787.460 2392.880 ;
        RECT 1644.140 15.000 1644.400 15.260 ;
        RECT 1787.200 15.340 1787.460 15.600 ;
      LAYER met2 ;
        RECT 1467.500 2392.590 1467.760 2392.910 ;
        RECT 1787.200 2392.590 1787.460 2392.910 ;
        RECT 1467.560 2377.880 1467.700 2392.590 ;
        RECT 1467.540 2373.880 1467.820 2377.880 ;
        RECT 1787.260 15.630 1787.400 2392.590 ;
        RECT 1787.200 15.310 1787.460 15.630 ;
        RECT 1644.140 14.970 1644.400 15.290 ;
        RECT 1644.200 2.400 1644.340 14.970 ;
        RECT 1643.990 -4.800 1644.550 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 711.230 73.000 711.550 73.060 ;
        RECT 1656.990 73.000 1657.310 73.060 ;
        RECT 711.230 72.860 1657.310 73.000 ;
        RECT 711.230 72.800 711.550 72.860 ;
        RECT 1656.990 72.800 1657.310 72.860 ;
      LAYER via ;
        RECT 711.260 72.800 711.520 73.060 ;
        RECT 1657.020 72.800 1657.280 73.060 ;
      LAYER met2 ;
        RECT 711.250 2225.115 711.530 2225.485 ;
        RECT 711.320 73.090 711.460 2225.115 ;
        RECT 711.260 72.770 711.520 73.090 ;
        RECT 1657.020 72.770 1657.280 73.090 ;
        RECT 1657.080 7.210 1657.220 72.770 ;
        RECT 1657.080 7.070 1662.280 7.210 ;
        RECT 1662.140 2.400 1662.280 7.070 ;
        RECT 1661.930 -4.800 1662.490 2.400 ;
      LAYER via2 ;
        RECT 711.250 2225.160 711.530 2225.440 ;
      LAYER met3 ;
        RECT 711.225 2225.450 711.555 2225.465 ;
        RECT 715.810 2225.450 719.810 2225.455 ;
        RECT 711.225 2225.150 719.810 2225.450 ;
        RECT 711.225 2225.135 711.555 2225.150 ;
        RECT 715.810 2224.855 719.810 2225.150 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 705.710 1308.560 706.030 1308.620 ;
        RECT 1676.770 1308.560 1677.090 1308.620 ;
        RECT 705.710 1308.420 1677.090 1308.560 ;
        RECT 705.710 1308.360 706.030 1308.420 ;
        RECT 1676.770 1308.360 1677.090 1308.420 ;
      LAYER via ;
        RECT 705.740 1308.360 706.000 1308.620 ;
        RECT 1676.800 1308.360 1677.060 1308.620 ;
      LAYER met2 ;
        RECT 705.730 1780.395 706.010 1780.765 ;
        RECT 705.800 1308.650 705.940 1780.395 ;
        RECT 705.740 1308.330 706.000 1308.650 ;
        RECT 1676.800 1308.330 1677.060 1308.650 ;
        RECT 1676.860 37.810 1677.000 1308.330 ;
        RECT 1676.860 37.670 1679.760 37.810 ;
        RECT 1679.620 2.400 1679.760 37.670 ;
        RECT 1679.410 -4.800 1679.970 2.400 ;
      LAYER via2 ;
        RECT 705.730 1780.440 706.010 1780.720 ;
      LAYER met3 ;
        RECT 705.705 1780.730 706.035 1780.745 ;
        RECT 715.810 1780.730 719.810 1780.735 ;
        RECT 705.705 1780.430 719.810 1780.730 ;
        RECT 705.705 1780.415 706.035 1780.430 ;
        RECT 715.810 1780.135 719.810 1780.430 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1762.865 1340.705 1763.035 1348.695 ;
      LAYER mcon ;
        RECT 1762.865 1348.525 1763.035 1348.695 ;
      LAYER met1 ;
        RECT 1762.790 1348.680 1763.110 1348.740 ;
        RECT 1762.595 1348.540 1763.110 1348.680 ;
        RECT 1762.790 1348.480 1763.110 1348.540 ;
        RECT 1761.870 1340.860 1762.190 1340.920 ;
        RECT 1762.805 1340.860 1763.095 1340.905 ;
        RECT 1761.870 1340.720 1763.095 1340.860 ;
        RECT 1761.870 1340.660 1762.190 1340.720 ;
        RECT 1762.805 1340.675 1763.095 1340.720 ;
        RECT 1703.910 1321.480 1704.230 1321.540 ;
        RECT 1761.870 1321.480 1762.190 1321.540 ;
        RECT 1703.910 1321.340 1762.190 1321.480 ;
        RECT 1703.910 1321.280 1704.230 1321.340 ;
        RECT 1761.870 1321.280 1762.190 1321.340 ;
        RECT 1697.470 18.940 1697.790 19.000 ;
        RECT 1703.910 18.940 1704.230 19.000 ;
        RECT 1697.470 18.800 1704.230 18.940 ;
        RECT 1697.470 18.740 1697.790 18.800 ;
        RECT 1703.910 18.740 1704.230 18.800 ;
      LAYER via ;
        RECT 1762.820 1348.480 1763.080 1348.740 ;
        RECT 1761.900 1340.660 1762.160 1340.920 ;
        RECT 1703.940 1321.280 1704.200 1321.540 ;
        RECT 1761.900 1321.280 1762.160 1321.540 ;
        RECT 1697.500 18.740 1697.760 19.000 ;
        RECT 1703.940 18.740 1704.200 19.000 ;
      LAYER met2 ;
        RECT 1762.810 2185.675 1763.090 2186.045 ;
        RECT 1762.880 1348.770 1763.020 2185.675 ;
        RECT 1762.820 1348.450 1763.080 1348.770 ;
        RECT 1761.900 1340.630 1762.160 1340.950 ;
        RECT 1761.960 1321.570 1762.100 1340.630 ;
        RECT 1703.940 1321.250 1704.200 1321.570 ;
        RECT 1761.900 1321.250 1762.160 1321.570 ;
        RECT 1704.000 19.030 1704.140 1321.250 ;
        RECT 1697.500 18.710 1697.760 19.030 ;
        RECT 1703.940 18.710 1704.200 19.030 ;
        RECT 1697.560 2.400 1697.700 18.710 ;
        RECT 1697.350 -4.800 1697.910 2.400 ;
      LAYER via2 ;
        RECT 1762.810 2185.720 1763.090 2186.000 ;
      LAYER met3 ;
        RECT 1755.835 2186.010 1759.835 2186.015 ;
        RECT 1762.785 2186.010 1763.115 2186.025 ;
        RECT 1755.835 2185.710 1763.115 2186.010 ;
        RECT 1755.835 2185.415 1759.835 2185.710 ;
        RECT 1762.785 2185.695 1763.115 2185.710 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 786.745 2394.025 787.835 2394.195 ;
      LAYER mcon ;
        RECT 787.665 2394.025 787.835 2394.195 ;
      LAYER met1 ;
        RECT 681.330 2394.180 681.650 2394.240 ;
        RECT 786.685 2394.180 786.975 2394.225 ;
        RECT 681.330 2394.040 786.975 2394.180 ;
        RECT 681.330 2393.980 681.650 2394.040 ;
        RECT 786.685 2393.995 786.975 2394.040 ;
        RECT 787.605 2394.180 787.895 2394.225 ;
        RECT 941.230 2394.180 941.550 2394.240 ;
        RECT 787.605 2394.040 941.550 2394.180 ;
        RECT 787.605 2393.995 787.895 2394.040 ;
        RECT 941.230 2393.980 941.550 2394.040 ;
        RECT 710.310 1310.600 710.630 1310.660 ;
        RECT 731.930 1310.600 732.250 1310.660 ;
        RECT 710.310 1310.460 732.250 1310.600 ;
        RECT 710.310 1310.400 710.630 1310.460 ;
        RECT 731.930 1310.400 732.250 1310.460 ;
        RECT 731.930 20.640 732.250 20.700 ;
        RECT 734.230 20.640 734.550 20.700 ;
        RECT 731.930 20.500 734.550 20.640 ;
        RECT 731.930 20.440 732.250 20.500 ;
        RECT 734.230 20.440 734.550 20.500 ;
      LAYER via ;
        RECT 681.360 2393.980 681.620 2394.240 ;
        RECT 941.260 2393.980 941.520 2394.240 ;
        RECT 710.340 1310.400 710.600 1310.660 ;
        RECT 731.960 1310.400 732.220 1310.660 ;
        RECT 731.960 20.440 732.220 20.700 ;
        RECT 734.260 20.440 734.520 20.700 ;
      LAYER met2 ;
        RECT 681.360 2393.950 681.620 2394.270 ;
        RECT 941.260 2393.950 941.520 2394.270 ;
        RECT 681.420 1327.885 681.560 2393.950 ;
        RECT 941.320 2377.880 941.460 2393.950 ;
        RECT 941.300 2373.880 941.580 2377.880 ;
        RECT 681.350 1327.515 681.630 1327.885 ;
        RECT 710.330 1327.515 710.610 1327.885 ;
        RECT 710.400 1310.690 710.540 1327.515 ;
        RECT 710.340 1310.370 710.600 1310.690 ;
        RECT 731.960 1310.370 732.220 1310.690 ;
        RECT 732.020 20.730 732.160 1310.370 ;
        RECT 731.960 20.410 732.220 20.730 ;
        RECT 734.260 20.410 734.520 20.730 ;
        RECT 734.320 2.400 734.460 20.410 ;
        RECT 734.110 -4.800 734.670 2.400 ;
      LAYER via2 ;
        RECT 681.350 1327.560 681.630 1327.840 ;
        RECT 710.330 1327.560 710.610 1327.840 ;
      LAYER met3 ;
        RECT 681.325 1327.850 681.655 1327.865 ;
        RECT 710.305 1327.850 710.635 1327.865 ;
        RECT 681.325 1327.550 710.635 1327.850 ;
        RECT 681.325 1327.535 681.655 1327.550 ;
        RECT 710.305 1327.535 710.635 1327.550 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1715.485 2.805 1715.655 48.195 ;
      LAYER mcon ;
        RECT 1715.485 48.025 1715.655 48.195 ;
      LAYER met1 ;
        RECT 710.770 72.660 711.090 72.720 ;
        RECT 1711.270 72.660 1711.590 72.720 ;
        RECT 710.770 72.520 1711.590 72.660 ;
        RECT 710.770 72.460 711.090 72.520 ;
        RECT 1711.270 72.460 1711.590 72.520 ;
        RECT 1711.270 48.180 1711.590 48.240 ;
        RECT 1715.425 48.180 1715.715 48.225 ;
        RECT 1711.270 48.040 1715.715 48.180 ;
        RECT 1711.270 47.980 1711.590 48.040 ;
        RECT 1715.425 47.995 1715.715 48.040 ;
        RECT 1715.410 2.960 1715.730 3.020 ;
        RECT 1715.215 2.820 1715.730 2.960 ;
        RECT 1715.410 2.760 1715.730 2.820 ;
      LAYER via ;
        RECT 710.800 72.460 711.060 72.720 ;
        RECT 1711.300 72.460 1711.560 72.720 ;
        RECT 1711.300 47.980 1711.560 48.240 ;
        RECT 1715.440 2.760 1715.700 3.020 ;
      LAYER met2 ;
        RECT 710.790 2233.275 711.070 2233.645 ;
        RECT 710.860 72.750 711.000 2233.275 ;
        RECT 710.800 72.430 711.060 72.750 ;
        RECT 1711.300 72.430 1711.560 72.750 ;
        RECT 1711.360 48.270 1711.500 72.430 ;
        RECT 1711.300 47.950 1711.560 48.270 ;
        RECT 1715.440 2.730 1715.700 3.050 ;
        RECT 1715.500 2.400 1715.640 2.730 ;
        RECT 1715.290 -4.800 1715.850 2.400 ;
      LAYER via2 ;
        RECT 710.790 2233.320 711.070 2233.600 ;
      LAYER met3 ;
        RECT 710.765 2233.610 711.095 2233.625 ;
        RECT 715.810 2233.610 719.810 2233.615 ;
        RECT 710.765 2233.310 719.810 2233.610 ;
        RECT 710.765 2233.295 711.095 2233.310 ;
        RECT 715.810 2233.015 719.810 2233.310 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1219.070 2382.960 1219.390 2383.020 ;
        RECT 1787.630 2382.960 1787.950 2383.020 ;
        RECT 1219.070 2382.820 1787.950 2382.960 ;
        RECT 1219.070 2382.760 1219.390 2382.820 ;
        RECT 1787.630 2382.760 1787.950 2382.820 ;
        RECT 1733.350 14.860 1733.670 14.920 ;
        RECT 1787.630 14.860 1787.950 14.920 ;
        RECT 1733.350 14.720 1787.950 14.860 ;
        RECT 1733.350 14.660 1733.670 14.720 ;
        RECT 1787.630 14.660 1787.950 14.720 ;
      LAYER via ;
        RECT 1219.100 2382.760 1219.360 2383.020 ;
        RECT 1787.660 2382.760 1787.920 2383.020 ;
        RECT 1733.380 14.660 1733.640 14.920 ;
        RECT 1787.660 14.660 1787.920 14.920 ;
      LAYER met2 ;
        RECT 1219.100 2382.730 1219.360 2383.050 ;
        RECT 1787.660 2382.730 1787.920 2383.050 ;
        RECT 1219.160 2377.880 1219.300 2382.730 ;
        RECT 1219.140 2373.880 1219.420 2377.880 ;
        RECT 1787.720 14.950 1787.860 2382.730 ;
        RECT 1733.380 14.630 1733.640 14.950 ;
        RECT 1787.660 14.630 1787.920 14.950 ;
        RECT 1733.440 2.400 1733.580 14.630 ;
        RECT 1733.230 -4.800 1733.790 2.400 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1276.110 33.560 1276.430 33.620 ;
        RECT 1751.290 33.560 1751.610 33.620 ;
        RECT 1276.110 33.420 1751.610 33.560 ;
        RECT 1276.110 33.360 1276.430 33.420 ;
        RECT 1751.290 33.360 1751.610 33.420 ;
      LAYER via ;
        RECT 1276.140 33.360 1276.400 33.620 ;
        RECT 1751.320 33.360 1751.580 33.620 ;
      LAYER met2 ;
        RECT 1273.420 1323.690 1273.700 1327.135 ;
        RECT 1273.420 1323.550 1276.340 1323.690 ;
        RECT 1273.420 1323.135 1273.700 1323.550 ;
        RECT 1276.200 33.650 1276.340 1323.550 ;
        RECT 1276.140 33.330 1276.400 33.650 ;
        RECT 1751.320 33.330 1751.580 33.650 ;
        RECT 1751.380 2.400 1751.520 33.330 ;
        RECT 1751.170 -4.800 1751.730 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1767.410 1689.275 1767.690 1689.645 ;
        RECT 1767.480 3.130 1767.620 1689.275 ;
        RECT 1767.480 2.990 1769.000 3.130 ;
        RECT 1768.860 2.400 1769.000 2.990 ;
        RECT 1768.650 -4.800 1769.210 2.400 ;
      LAYER via2 ;
        RECT 1767.410 1689.320 1767.690 1689.600 ;
      LAYER met3 ;
        RECT 1755.835 1689.610 1759.835 1689.615 ;
        RECT 1767.385 1689.610 1767.715 1689.625 ;
        RECT 1755.835 1689.310 1767.715 1689.610 ;
        RECT 1755.835 1689.015 1759.835 1689.310 ;
        RECT 1767.385 1689.295 1767.715 1689.310 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1498.750 1311.280 1499.070 1311.340 ;
        RECT 1503.810 1311.280 1504.130 1311.340 ;
        RECT 1498.750 1311.140 1504.130 1311.280 ;
        RECT 1498.750 1311.080 1499.070 1311.140 ;
        RECT 1503.810 1311.080 1504.130 1311.140 ;
        RECT 1503.810 32.200 1504.130 32.260 ;
        RECT 1786.710 32.200 1787.030 32.260 ;
        RECT 1503.810 32.060 1787.030 32.200 ;
        RECT 1503.810 32.000 1504.130 32.060 ;
        RECT 1786.710 32.000 1787.030 32.060 ;
      LAYER via ;
        RECT 1498.780 1311.080 1499.040 1311.340 ;
        RECT 1503.840 1311.080 1504.100 1311.340 ;
        RECT 1503.840 32.000 1504.100 32.260 ;
        RECT 1786.740 32.000 1787.000 32.260 ;
      LAYER met2 ;
        RECT 1498.820 1323.135 1499.100 1327.135 ;
        RECT 1498.840 1311.370 1498.980 1323.135 ;
        RECT 1498.780 1311.050 1499.040 1311.370 ;
        RECT 1503.840 1311.050 1504.100 1311.370 ;
        RECT 1503.900 32.290 1504.040 1311.050 ;
        RECT 1503.840 31.970 1504.100 32.290 ;
        RECT 1786.740 31.970 1787.000 32.290 ;
        RECT 1786.800 2.400 1786.940 31.970 ;
        RECT 1786.590 -4.800 1787.150 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 955.030 1311.280 955.350 1311.340 ;
        RECT 958.710 1311.280 959.030 1311.340 ;
        RECT 955.030 1311.140 959.030 1311.280 ;
        RECT 955.030 1311.080 955.350 1311.140 ;
        RECT 958.710 1311.080 959.030 1311.140 ;
        RECT 958.710 41.040 959.030 41.100 ;
        RECT 1804.650 41.040 1804.970 41.100 ;
        RECT 958.710 40.900 1804.970 41.040 ;
        RECT 958.710 40.840 959.030 40.900 ;
        RECT 1804.650 40.840 1804.970 40.900 ;
      LAYER via ;
        RECT 955.060 1311.080 955.320 1311.340 ;
        RECT 958.740 1311.080 959.000 1311.340 ;
        RECT 958.740 40.840 959.000 41.100 ;
        RECT 1804.680 40.840 1804.940 41.100 ;
      LAYER met2 ;
        RECT 955.100 1323.135 955.380 1327.135 ;
        RECT 955.120 1311.370 955.260 1323.135 ;
        RECT 955.060 1311.050 955.320 1311.370 ;
        RECT 958.740 1311.050 959.000 1311.370 ;
        RECT 958.800 41.130 958.940 1311.050 ;
        RECT 958.740 40.810 959.000 41.130 ;
        RECT 1804.680 40.810 1804.940 41.130 ;
        RECT 1804.740 2.400 1804.880 40.810 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1652.925 2387.565 1653.095 2389.435 ;
      LAYER mcon ;
        RECT 1652.925 2389.265 1653.095 2389.435 ;
      LAYER met1 ;
        RECT 1633.530 2389.420 1633.850 2389.480 ;
        RECT 1652.865 2389.420 1653.155 2389.465 ;
        RECT 1633.530 2389.280 1653.155 2389.420 ;
        RECT 1633.530 2389.220 1633.850 2389.280 ;
        RECT 1652.865 2389.235 1653.155 2389.280 ;
        RECT 1652.865 2387.720 1653.155 2387.765 ;
        RECT 1757.270 2387.720 1757.590 2387.780 ;
        RECT 1652.865 2387.580 1757.590 2387.720 ;
        RECT 1652.865 2387.535 1653.155 2387.580 ;
        RECT 1757.270 2387.520 1757.590 2387.580 ;
        RECT 1757.730 2308.160 1758.050 2308.220 ;
        RECT 1821.670 2308.160 1821.990 2308.220 ;
        RECT 1757.730 2308.020 1821.990 2308.160 ;
        RECT 1757.730 2307.960 1758.050 2308.020 ;
        RECT 1821.670 2307.960 1821.990 2308.020 ;
      LAYER via ;
        RECT 1633.560 2389.220 1633.820 2389.480 ;
        RECT 1757.300 2387.520 1757.560 2387.780 ;
        RECT 1757.760 2307.960 1758.020 2308.220 ;
        RECT 1821.700 2307.960 1821.960 2308.220 ;
      LAYER met2 ;
        RECT 1633.560 2389.190 1633.820 2389.510 ;
        RECT 1633.620 2378.370 1633.760 2389.190 ;
        RECT 1757.300 2387.490 1757.560 2387.810 ;
        RECT 1631.320 2378.230 1633.760 2378.370 ;
        RECT 1629.460 2377.690 1629.740 2377.880 ;
        RECT 1631.320 2377.690 1631.460 2378.230 ;
        RECT 1629.460 2377.550 1631.460 2377.690 ;
        RECT 1629.460 2373.880 1629.740 2377.550 ;
        RECT 1757.360 2314.450 1757.500 2387.490 ;
        RECT 1757.360 2314.310 1757.960 2314.450 ;
        RECT 1757.820 2308.250 1757.960 2314.310 ;
        RECT 1757.760 2307.930 1758.020 2308.250 ;
        RECT 1821.700 2307.930 1821.960 2308.250 ;
        RECT 1821.760 16.730 1821.900 2307.930 ;
        RECT 1821.760 16.590 1822.820 16.730 ;
        RECT 1822.680 2.400 1822.820 16.590 ;
        RECT 1822.470 -4.800 1823.030 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 718.665 1884.705 718.835 1928.735 ;
        RECT 718.665 1802.085 718.835 1845.775 ;
        RECT 718.665 1476.705 718.835 1658.775 ;
        RECT 716.825 1429.445 716.995 1453.075 ;
        RECT 717.285 1403.265 717.455 1406.495 ;
        RECT 717.285 1353.625 717.455 1374.535 ;
      LAYER mcon ;
        RECT 718.665 1928.565 718.835 1928.735 ;
        RECT 718.665 1845.605 718.835 1845.775 ;
        RECT 718.665 1658.605 718.835 1658.775 ;
        RECT 716.825 1452.905 716.995 1453.075 ;
        RECT 717.285 1406.325 717.455 1406.495 ;
        RECT 717.285 1374.365 717.455 1374.535 ;
      LAYER met1 ;
        RECT 718.590 1928.720 718.910 1928.780 ;
        RECT 718.395 1928.580 718.910 1928.720 ;
        RECT 718.590 1928.520 718.910 1928.580 ;
        RECT 718.590 1884.860 718.910 1884.920 ;
        RECT 718.395 1884.720 718.910 1884.860 ;
        RECT 718.590 1884.660 718.910 1884.720 ;
        RECT 718.590 1845.760 718.910 1845.820 ;
        RECT 718.395 1845.620 718.910 1845.760 ;
        RECT 718.590 1845.560 718.910 1845.620 ;
        RECT 718.590 1802.240 718.910 1802.300 ;
        RECT 718.395 1802.100 718.910 1802.240 ;
        RECT 718.590 1802.040 718.910 1802.100 ;
        RECT 718.590 1658.760 718.910 1658.820 ;
        RECT 718.395 1658.620 718.910 1658.760 ;
        RECT 718.590 1658.560 718.910 1658.620 ;
        RECT 717.210 1476.860 717.530 1476.920 ;
        RECT 718.605 1476.860 718.895 1476.905 ;
        RECT 717.210 1476.720 718.895 1476.860 ;
        RECT 717.210 1476.660 717.530 1476.720 ;
        RECT 718.605 1476.675 718.895 1476.720 ;
        RECT 716.750 1453.060 717.070 1453.120 ;
        RECT 716.555 1452.920 717.070 1453.060 ;
        RECT 716.750 1452.860 717.070 1452.920 ;
        RECT 716.765 1429.600 717.055 1429.645 ;
        RECT 717.210 1429.600 717.530 1429.660 ;
        RECT 716.765 1429.460 717.530 1429.600 ;
        RECT 716.765 1429.415 717.055 1429.460 ;
        RECT 717.210 1429.400 717.530 1429.460 ;
        RECT 717.210 1406.480 717.530 1406.540 ;
        RECT 717.015 1406.340 717.530 1406.480 ;
        RECT 717.210 1406.280 717.530 1406.340 ;
        RECT 717.210 1403.420 717.530 1403.480 ;
        RECT 717.015 1403.280 717.530 1403.420 ;
        RECT 717.210 1403.220 717.530 1403.280 ;
        RECT 717.210 1374.520 717.530 1374.580 ;
        RECT 717.015 1374.380 717.530 1374.520 ;
        RECT 717.210 1374.320 717.530 1374.380 ;
        RECT 717.210 1353.780 717.530 1353.840 ;
        RECT 717.015 1353.640 717.530 1353.780 ;
        RECT 717.210 1353.580 717.530 1353.640 ;
      LAYER via ;
        RECT 718.620 1928.520 718.880 1928.780 ;
        RECT 718.620 1884.660 718.880 1884.920 ;
        RECT 718.620 1845.560 718.880 1845.820 ;
        RECT 718.620 1802.040 718.880 1802.300 ;
        RECT 718.620 1658.560 718.880 1658.820 ;
        RECT 717.240 1476.660 717.500 1476.920 ;
        RECT 716.780 1452.860 717.040 1453.120 ;
        RECT 717.240 1429.400 717.500 1429.660 ;
        RECT 717.240 1406.280 717.500 1406.540 ;
        RECT 717.240 1403.220 717.500 1403.480 ;
        RECT 717.240 1374.320 717.500 1374.580 ;
        RECT 717.240 1353.580 717.500 1353.840 ;
      LAYER met2 ;
        RECT 718.610 1991.195 718.890 1991.565 ;
        RECT 718.680 1928.810 718.820 1991.195 ;
        RECT 718.620 1928.490 718.880 1928.810 ;
        RECT 718.620 1884.630 718.880 1884.950 ;
        RECT 718.680 1845.850 718.820 1884.630 ;
        RECT 718.620 1845.530 718.880 1845.850 ;
        RECT 718.620 1802.010 718.880 1802.330 ;
        RECT 718.680 1658.850 718.820 1802.010 ;
        RECT 718.620 1658.530 718.880 1658.850 ;
        RECT 717.240 1476.805 717.500 1476.950 ;
        RECT 717.230 1476.435 717.510 1476.805 ;
        RECT 716.770 1468.275 717.050 1468.645 ;
        RECT 716.840 1453.150 716.980 1468.275 ;
        RECT 716.780 1452.830 717.040 1453.150 ;
        RECT 717.240 1429.370 717.500 1429.690 ;
        RECT 717.300 1406.570 717.440 1429.370 ;
        RECT 717.240 1406.250 717.500 1406.570 ;
        RECT 717.240 1403.190 717.500 1403.510 ;
        RECT 717.300 1374.610 717.440 1403.190 ;
        RECT 717.240 1374.290 717.500 1374.610 ;
        RECT 717.240 1353.725 717.500 1353.870 ;
        RECT 717.230 1353.355 717.510 1353.725 ;
        RECT 1835.490 888.915 1835.770 889.285 ;
        RECT 1835.560 16.730 1835.700 888.915 ;
        RECT 1835.560 16.590 1840.300 16.730 ;
        RECT 1840.160 2.400 1840.300 16.590 ;
        RECT 1839.950 -4.800 1840.510 2.400 ;
      LAYER via2 ;
        RECT 718.610 1991.240 718.890 1991.520 ;
        RECT 717.230 1476.480 717.510 1476.760 ;
        RECT 716.770 1468.320 717.050 1468.600 ;
        RECT 717.230 1353.400 717.510 1353.680 ;
        RECT 1835.490 888.960 1835.770 889.240 ;
      LAYER met3 ;
        RECT 715.810 1993.655 719.810 1994.255 ;
        RECT 718.830 1991.545 719.130 1993.655 ;
        RECT 718.585 1991.230 719.130 1991.545 ;
        RECT 718.585 1991.215 718.915 1991.230 ;
        RECT 717.205 1476.770 717.535 1476.785 ;
        RECT 718.790 1476.770 719.170 1476.780 ;
        RECT 717.205 1476.470 719.170 1476.770 ;
        RECT 717.205 1476.455 717.535 1476.470 ;
        RECT 718.790 1476.460 719.170 1476.470 ;
        RECT 718.790 1468.980 719.170 1469.300 ;
        RECT 716.745 1468.610 717.075 1468.625 ;
        RECT 718.830 1468.610 719.130 1468.980 ;
        RECT 716.745 1468.310 719.130 1468.610 ;
        RECT 716.745 1468.295 717.075 1468.310 ;
        RECT 717.205 1353.700 717.535 1353.705 ;
        RECT 716.950 1353.690 717.535 1353.700 ;
        RECT 716.750 1353.390 717.535 1353.690 ;
        RECT 716.950 1353.380 717.535 1353.390 ;
        RECT 717.205 1353.375 717.535 1353.380 ;
        RECT 716.950 1340.770 717.330 1340.780 ;
        RECT 718.790 1340.770 719.170 1340.780 ;
        RECT 716.950 1340.470 719.170 1340.770 ;
        RECT 716.950 1340.460 717.330 1340.470 ;
        RECT 718.790 1340.460 719.170 1340.470 ;
        RECT 718.790 889.250 719.170 889.260 ;
        RECT 1835.465 889.250 1835.795 889.265 ;
        RECT 718.790 888.950 1835.795 889.250 ;
        RECT 718.790 888.940 719.170 888.950 ;
        RECT 1835.465 888.935 1835.795 888.950 ;
      LAYER via3 ;
        RECT 718.820 1476.460 719.140 1476.780 ;
        RECT 718.820 1468.980 719.140 1469.300 ;
        RECT 716.980 1353.380 717.300 1353.700 ;
        RECT 716.980 1340.460 717.300 1340.780 ;
        RECT 718.820 1340.460 719.140 1340.780 ;
        RECT 718.820 888.940 719.140 889.260 ;
      LAYER met4 ;
        RECT 718.815 1476.455 719.145 1476.785 ;
        RECT 718.830 1469.305 719.130 1476.455 ;
        RECT 718.815 1468.975 719.145 1469.305 ;
        RECT 716.975 1353.375 717.305 1353.705 ;
        RECT 716.990 1340.785 717.290 1353.375 ;
        RECT 716.975 1340.455 717.305 1340.785 ;
        RECT 718.815 1340.455 719.145 1340.785 ;
        RECT 718.830 889.265 719.130 1340.455 ;
        RECT 718.815 888.935 719.145 889.265 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 701.645 1352.605 701.815 1393.575 ;
      LAYER mcon ;
        RECT 701.645 1393.405 701.815 1393.575 ;
      LAYER met1 ;
        RECT 701.570 1393.560 701.890 1393.620 ;
        RECT 701.570 1393.420 702.085 1393.560 ;
        RECT 701.570 1393.360 701.890 1393.420 ;
        RECT 701.570 1352.760 701.890 1352.820 ;
        RECT 701.375 1352.620 701.890 1352.760 ;
        RECT 701.570 1352.560 701.890 1352.620 ;
        RECT 701.570 93.060 701.890 93.120 ;
        RECT 1856.170 93.060 1856.490 93.120 ;
        RECT 701.570 92.920 1856.490 93.060 ;
        RECT 701.570 92.860 701.890 92.920 ;
        RECT 1856.170 92.860 1856.490 92.920 ;
      LAYER via ;
        RECT 701.600 1393.360 701.860 1393.620 ;
        RECT 701.600 1352.560 701.860 1352.820 ;
        RECT 701.600 92.860 701.860 93.120 ;
        RECT 1856.200 92.860 1856.460 93.120 ;
      LAYER met2 ;
        RECT 701.590 1925.915 701.870 1926.285 ;
        RECT 701.660 1393.650 701.800 1925.915 ;
        RECT 701.600 1393.330 701.860 1393.650 ;
        RECT 701.600 1352.530 701.860 1352.850 ;
        RECT 701.660 93.150 701.800 1352.530 ;
        RECT 701.600 92.830 701.860 93.150 ;
        RECT 1856.200 92.830 1856.460 93.150 ;
        RECT 1856.260 19.960 1856.400 92.830 ;
        RECT 1856.260 19.820 1857.320 19.960 ;
        RECT 1857.180 12.650 1857.320 19.820 ;
        RECT 1857.180 12.510 1858.240 12.650 ;
        RECT 1858.100 2.400 1858.240 12.510 ;
        RECT 1857.890 -4.800 1858.450 2.400 ;
      LAYER via2 ;
        RECT 701.590 1925.960 701.870 1926.240 ;
      LAYER met3 ;
        RECT 701.565 1926.250 701.895 1926.265 ;
        RECT 715.810 1926.250 719.810 1926.255 ;
        RECT 701.565 1925.950 719.810 1926.250 ;
        RECT 701.565 1925.935 701.895 1925.950 ;
        RECT 715.810 1925.655 719.810 1925.950 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1771.990 2242.880 1772.310 2242.940 ;
        RECT 1824.890 2242.880 1825.210 2242.940 ;
        RECT 1771.990 2242.740 1825.210 2242.880 ;
        RECT 1771.990 2242.680 1772.310 2242.740 ;
        RECT 1824.890 2242.680 1825.210 2242.740 ;
        RECT 1824.890 19.280 1825.210 19.340 ;
        RECT 1875.950 19.280 1876.270 19.340 ;
        RECT 1824.890 19.140 1876.270 19.280 ;
        RECT 1824.890 19.080 1825.210 19.140 ;
        RECT 1875.950 19.080 1876.270 19.140 ;
      LAYER via ;
        RECT 1772.020 2242.680 1772.280 2242.940 ;
        RECT 1824.920 2242.680 1825.180 2242.940 ;
        RECT 1824.920 19.080 1825.180 19.340 ;
        RECT 1875.980 19.080 1876.240 19.340 ;
      LAYER met2 ;
        RECT 1772.010 2245.515 1772.290 2245.885 ;
        RECT 1772.080 2242.970 1772.220 2245.515 ;
        RECT 1772.020 2242.650 1772.280 2242.970 ;
        RECT 1824.920 2242.650 1825.180 2242.970 ;
        RECT 1824.980 19.370 1825.120 2242.650 ;
        RECT 1824.920 19.050 1825.180 19.370 ;
        RECT 1875.980 19.050 1876.240 19.370 ;
        RECT 1876.040 2.400 1876.180 19.050 ;
        RECT 1875.830 -4.800 1876.390 2.400 ;
      LAYER via2 ;
        RECT 1772.010 2245.560 1772.290 2245.840 ;
      LAYER met3 ;
        RECT 1755.835 2245.850 1759.835 2245.855 ;
        RECT 1771.985 2245.850 1772.315 2245.865 ;
        RECT 1755.835 2245.550 1772.315 2245.850 ;
        RECT 1755.835 2245.255 1759.835 2245.550 ;
        RECT 1771.985 2245.535 1772.315 2245.550 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 710.310 1567.640 710.630 1567.700 ;
        RECT 713.990 1567.640 714.310 1567.700 ;
        RECT 710.310 1567.500 714.310 1567.640 ;
        RECT 710.310 1567.440 710.630 1567.500 ;
        RECT 713.990 1567.440 714.310 1567.500 ;
        RECT 713.990 15.200 714.310 15.260 ;
        RECT 752.170 15.200 752.490 15.260 ;
        RECT 713.990 15.060 752.490 15.200 ;
        RECT 713.990 15.000 714.310 15.060 ;
        RECT 752.170 15.000 752.490 15.060 ;
      LAYER via ;
        RECT 710.340 1567.440 710.600 1567.700 ;
        RECT 714.020 1567.440 714.280 1567.700 ;
        RECT 714.020 15.000 714.280 15.260 ;
        RECT 752.200 15.000 752.460 15.260 ;
      LAYER met2 ;
        RECT 710.330 1575.035 710.610 1575.405 ;
        RECT 710.400 1567.730 710.540 1575.035 ;
        RECT 710.340 1567.410 710.600 1567.730 ;
        RECT 714.020 1567.410 714.280 1567.730 ;
        RECT 714.080 15.290 714.220 1567.410 ;
        RECT 714.020 14.970 714.280 15.290 ;
        RECT 752.200 14.970 752.460 15.290 ;
        RECT 752.260 2.400 752.400 14.970 ;
        RECT 752.050 -4.800 752.610 2.400 ;
      LAYER via2 ;
        RECT 710.330 1575.080 710.610 1575.360 ;
      LAYER met3 ;
        RECT 710.305 1575.370 710.635 1575.385 ;
        RECT 715.810 1575.370 719.810 1575.375 ;
        RECT 710.305 1575.070 719.810 1575.370 ;
        RECT 710.305 1575.055 710.635 1575.070 ;
        RECT 715.810 1574.775 719.810 1575.070 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1890.690 93.315 1890.970 93.685 ;
        RECT 1890.760 18.770 1890.900 93.315 ;
        RECT 1890.760 18.630 1894.120 18.770 ;
        RECT 1893.980 2.400 1894.120 18.630 ;
        RECT 1893.770 -4.800 1894.330 2.400 ;
      LAYER via2 ;
        RECT 1890.690 93.360 1890.970 93.640 ;
      LAYER met3 ;
        RECT 702.230 2251.290 702.610 2251.300 ;
        RECT 715.810 2251.290 719.810 2251.295 ;
        RECT 702.230 2250.990 719.810 2251.290 ;
        RECT 702.230 2250.980 702.610 2250.990 ;
        RECT 715.810 2250.695 719.810 2250.990 ;
        RECT 702.230 93.650 702.610 93.660 ;
        RECT 1890.665 93.650 1890.995 93.665 ;
        RECT 702.230 93.350 1890.995 93.650 ;
        RECT 702.230 93.340 702.610 93.350 ;
        RECT 1890.665 93.335 1890.995 93.350 ;
      LAYER via3 ;
        RECT 702.260 2250.980 702.580 2251.300 ;
        RECT 702.260 93.340 702.580 93.660 ;
      LAYER met4 ;
        RECT 702.255 2250.975 702.585 2251.305 ;
        RECT 702.270 93.665 702.570 2250.975 ;
        RECT 702.255 93.335 702.585 93.665 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1432.510 2390.440 1432.830 2390.500 ;
        RECT 1873.190 2390.440 1873.510 2390.500 ;
        RECT 1432.510 2390.300 1873.510 2390.440 ;
        RECT 1432.510 2390.240 1432.830 2390.300 ;
        RECT 1873.190 2390.240 1873.510 2390.300 ;
        RECT 1873.190 19.620 1873.510 19.680 ;
        RECT 1911.830 19.620 1912.150 19.680 ;
        RECT 1873.190 19.480 1912.150 19.620 ;
        RECT 1873.190 19.420 1873.510 19.480 ;
        RECT 1911.830 19.420 1912.150 19.480 ;
      LAYER via ;
        RECT 1432.540 2390.240 1432.800 2390.500 ;
        RECT 1873.220 2390.240 1873.480 2390.500 ;
        RECT 1873.220 19.420 1873.480 19.680 ;
        RECT 1911.860 19.420 1912.120 19.680 ;
      LAYER met2 ;
        RECT 1432.540 2390.210 1432.800 2390.530 ;
        RECT 1873.220 2390.210 1873.480 2390.530 ;
        RECT 1432.600 2377.880 1432.740 2390.210 ;
        RECT 1432.580 2373.880 1432.860 2377.880 ;
        RECT 1873.280 19.710 1873.420 2390.210 ;
        RECT 1873.220 19.390 1873.480 19.710 ;
        RECT 1911.860 19.390 1912.120 19.710 ;
        RECT 1911.920 2.400 1912.060 19.390 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1652.465 2389.605 1652.635 2391.135 ;
      LAYER mcon ;
        RECT 1652.465 2390.965 1652.635 2391.135 ;
      LAYER met1 ;
        RECT 1652.405 2391.120 1652.695 2391.165 ;
        RECT 1914.590 2391.120 1914.910 2391.180 ;
        RECT 1652.405 2390.980 1914.910 2391.120 ;
        RECT 1652.405 2390.935 1652.695 2390.980 ;
        RECT 1914.590 2390.920 1914.910 2390.980 ;
        RECT 1600.870 2389.760 1601.190 2389.820 ;
        RECT 1652.405 2389.760 1652.695 2389.805 ;
        RECT 1600.870 2389.620 1652.695 2389.760 ;
        RECT 1600.870 2389.560 1601.190 2389.620 ;
        RECT 1652.405 2389.575 1652.695 2389.620 ;
        RECT 1914.590 20.640 1914.910 20.700 ;
        RECT 1929.310 20.640 1929.630 20.700 ;
        RECT 1914.590 20.500 1929.630 20.640 ;
        RECT 1914.590 20.440 1914.910 20.500 ;
        RECT 1929.310 20.440 1929.630 20.500 ;
      LAYER via ;
        RECT 1914.620 2390.920 1914.880 2391.180 ;
        RECT 1600.900 2389.560 1601.160 2389.820 ;
        RECT 1914.620 20.440 1914.880 20.700 ;
        RECT 1929.340 20.440 1929.600 20.700 ;
      LAYER met2 ;
        RECT 1914.620 2390.890 1914.880 2391.210 ;
        RECT 1600.900 2389.530 1601.160 2389.850 ;
        RECT 1600.960 2377.880 1601.100 2389.530 ;
        RECT 1600.940 2373.880 1601.220 2377.880 ;
        RECT 1914.680 20.730 1914.820 2390.890 ;
        RECT 1914.620 20.410 1914.880 20.730 ;
        RECT 1929.340 20.410 1929.600 20.730 ;
        RECT 1929.400 2.400 1929.540 20.410 ;
        RECT 1929.190 -4.800 1929.750 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1937.130 48.520 1937.450 48.580 ;
        RECT 1947.250 48.520 1947.570 48.580 ;
        RECT 1937.130 48.380 1947.570 48.520 ;
        RECT 1937.130 48.320 1937.450 48.380 ;
        RECT 1947.250 48.320 1947.570 48.380 ;
      LAYER via ;
        RECT 1937.160 48.320 1937.420 48.580 ;
        RECT 1947.280 48.320 1947.540 48.580 ;
      LAYER met2 ;
        RECT 1937.150 92.635 1937.430 93.005 ;
        RECT 1937.220 48.610 1937.360 92.635 ;
        RECT 1937.160 48.290 1937.420 48.610 ;
        RECT 1947.280 48.290 1947.540 48.610 ;
        RECT 1947.340 2.400 1947.480 48.290 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
      LAYER via2 ;
        RECT 1937.150 92.680 1937.430 92.960 ;
      LAYER met3 ;
        RECT 703.150 2293.450 703.530 2293.460 ;
        RECT 715.810 2293.450 719.810 2293.455 ;
        RECT 703.150 2293.150 719.810 2293.450 ;
        RECT 703.150 2293.140 703.530 2293.150 ;
        RECT 715.810 2292.855 719.810 2293.150 ;
        RECT 703.150 92.970 703.530 92.980 ;
        RECT 1937.125 92.970 1937.455 92.985 ;
        RECT 703.150 92.670 1937.455 92.970 ;
        RECT 703.150 92.660 703.530 92.670 ;
        RECT 1937.125 92.655 1937.455 92.670 ;
      LAYER via3 ;
        RECT 703.180 2293.140 703.500 2293.460 ;
        RECT 703.180 92.660 703.500 92.980 ;
      LAYER met4 ;
        RECT 703.175 2293.135 703.505 2293.465 ;
        RECT 703.190 92.985 703.490 2293.135 ;
        RECT 703.175 92.655 703.505 92.985 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1772.910 1594.160 1773.230 1594.220 ;
        RECT 1949.090 1594.160 1949.410 1594.220 ;
        RECT 1772.910 1594.020 1949.410 1594.160 ;
        RECT 1772.910 1593.960 1773.230 1594.020 ;
        RECT 1949.090 1593.960 1949.410 1594.020 ;
        RECT 1949.090 20.640 1949.410 20.700 ;
        RECT 1965.190 20.640 1965.510 20.700 ;
        RECT 1949.090 20.500 1965.510 20.640 ;
        RECT 1949.090 20.440 1949.410 20.500 ;
        RECT 1965.190 20.440 1965.510 20.500 ;
      LAYER via ;
        RECT 1772.940 1593.960 1773.200 1594.220 ;
        RECT 1949.120 1593.960 1949.380 1594.220 ;
        RECT 1949.120 20.440 1949.380 20.700 ;
        RECT 1965.220 20.440 1965.480 20.700 ;
      LAYER met2 ;
        RECT 1772.930 1595.435 1773.210 1595.805 ;
        RECT 1773.000 1594.250 1773.140 1595.435 ;
        RECT 1772.940 1593.930 1773.200 1594.250 ;
        RECT 1949.120 1593.930 1949.380 1594.250 ;
        RECT 1949.180 20.730 1949.320 1593.930 ;
        RECT 1949.120 20.410 1949.380 20.730 ;
        RECT 1965.220 20.410 1965.480 20.730 ;
        RECT 1965.280 2.400 1965.420 20.410 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
      LAYER via2 ;
        RECT 1772.930 1595.480 1773.210 1595.760 ;
      LAYER met3 ;
        RECT 1755.835 1595.770 1759.835 1595.775 ;
        RECT 1772.905 1595.770 1773.235 1595.785 ;
        RECT 1755.835 1595.470 1773.235 1595.770 ;
        RECT 1755.835 1595.175 1759.835 1595.470 ;
        RECT 1772.905 1595.455 1773.235 1595.470 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1020.810 40.360 1021.130 40.420 ;
        RECT 1983.130 40.360 1983.450 40.420 ;
        RECT 1020.810 40.220 1983.450 40.360 ;
        RECT 1020.810 40.160 1021.130 40.220 ;
        RECT 1983.130 40.160 1983.450 40.220 ;
      LAYER via ;
        RECT 1020.840 40.160 1021.100 40.420 ;
        RECT 1983.160 40.160 1983.420 40.420 ;
      LAYER met2 ;
        RECT 1018.580 1323.690 1018.860 1327.135 ;
        RECT 1018.580 1323.550 1021.040 1323.690 ;
        RECT 1018.580 1323.135 1018.860 1323.550 ;
        RECT 1020.900 40.450 1021.040 1323.550 ;
        RECT 1020.840 40.130 1021.100 40.450 ;
        RECT 1983.160 40.130 1983.420 40.450 ;
        RECT 1983.220 2.400 1983.360 40.130 ;
        RECT 1983.010 -4.800 1983.570 2.400 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1151.910 40.700 1152.230 40.760 ;
        RECT 2001.070 40.700 2001.390 40.760 ;
        RECT 1151.910 40.560 2001.390 40.700 ;
        RECT 1151.910 40.500 1152.230 40.560 ;
        RECT 2001.070 40.500 2001.390 40.560 ;
      LAYER via ;
        RECT 1151.940 40.500 1152.200 40.760 ;
        RECT 2001.100 40.500 2001.360 40.760 ;
      LAYER met2 ;
        RECT 1151.980 1323.135 1152.260 1327.135 ;
        RECT 1152.000 40.790 1152.140 1323.135 ;
        RECT 1151.940 40.470 1152.200 40.790 ;
        RECT 2001.100 40.470 2001.360 40.790 ;
        RECT 2001.160 2.400 2001.300 40.470 ;
        RECT 2000.950 -4.800 2001.510 2.400 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 969.750 2389.080 970.070 2389.140 ;
        RECT 1757.730 2389.080 1758.050 2389.140 ;
        RECT 969.750 2388.940 1758.050 2389.080 ;
        RECT 969.750 2388.880 970.070 2388.940 ;
        RECT 1757.730 2388.880 1758.050 2388.940 ;
        RECT 1757.730 2314.960 1758.050 2315.020 ;
        RECT 2014.870 2314.960 2015.190 2315.020 ;
        RECT 1757.730 2314.820 2015.190 2314.960 ;
        RECT 1757.730 2314.760 1758.050 2314.820 ;
        RECT 2014.870 2314.760 2015.190 2314.820 ;
        RECT 2014.870 2.960 2015.190 3.020 ;
        RECT 2018.550 2.960 2018.870 3.020 ;
        RECT 2014.870 2.820 2018.870 2.960 ;
        RECT 2014.870 2.760 2015.190 2.820 ;
        RECT 2018.550 2.760 2018.870 2.820 ;
      LAYER via ;
        RECT 969.780 2388.880 970.040 2389.140 ;
        RECT 1757.760 2388.880 1758.020 2389.140 ;
        RECT 1757.760 2314.760 1758.020 2315.020 ;
        RECT 2014.900 2314.760 2015.160 2315.020 ;
        RECT 2014.900 2.760 2015.160 3.020 ;
        RECT 2018.580 2.760 2018.840 3.020 ;
      LAYER met2 ;
        RECT 969.780 2388.850 970.040 2389.170 ;
        RECT 1757.760 2388.850 1758.020 2389.170 ;
        RECT 969.840 2377.880 969.980 2388.850 ;
        RECT 969.820 2373.880 970.100 2377.880 ;
        RECT 1757.820 2315.050 1757.960 2388.850 ;
        RECT 1757.760 2314.730 1758.020 2315.050 ;
        RECT 2014.900 2314.730 2015.160 2315.050 ;
        RECT 2014.960 3.050 2015.100 2314.730 ;
        RECT 2014.900 2.730 2015.160 3.050 ;
        RECT 2018.580 2.730 2018.840 3.050 ;
        RECT 2018.640 2.400 2018.780 2.730 ;
        RECT 2018.430 -4.800 2018.990 2.400 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1259.550 2388.740 1259.870 2388.800 ;
        RECT 2035.570 2388.740 2035.890 2388.800 ;
        RECT 1259.550 2388.600 2035.890 2388.740 ;
        RECT 1259.550 2388.540 1259.870 2388.600 ;
        RECT 2035.570 2388.540 2035.890 2388.600 ;
      LAYER via ;
        RECT 1259.580 2388.540 1259.840 2388.800 ;
        RECT 2035.600 2388.540 2035.860 2388.800 ;
      LAYER met2 ;
        RECT 1259.580 2388.510 1259.840 2388.830 ;
        RECT 2035.600 2388.510 2035.860 2388.830 ;
        RECT 1259.640 2377.880 1259.780 2388.510 ;
        RECT 1259.620 2373.880 1259.900 2377.880 ;
        RECT 2035.660 3.130 2035.800 2388.510 ;
        RECT 2035.660 2.990 2036.720 3.130 ;
        RECT 2036.580 2.400 2036.720 2.990 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1772.450 2001.140 1772.770 2001.200 ;
        RECT 1893.890 2001.140 1894.210 2001.200 ;
        RECT 1772.450 2001.000 1894.210 2001.140 ;
        RECT 1772.450 2000.940 1772.770 2001.000 ;
        RECT 1893.890 2000.940 1894.210 2001.000 ;
        RECT 2054.430 19.960 2054.750 20.020 ;
        RECT 1995.640 19.820 2054.750 19.960 ;
        RECT 1893.890 19.280 1894.210 19.340 ;
        RECT 1995.640 19.280 1995.780 19.820 ;
        RECT 2054.430 19.760 2054.750 19.820 ;
        RECT 1893.890 19.140 1995.780 19.280 ;
        RECT 1893.890 19.080 1894.210 19.140 ;
      LAYER via ;
        RECT 1772.480 2000.940 1772.740 2001.200 ;
        RECT 1893.920 2000.940 1894.180 2001.200 ;
        RECT 1893.920 19.080 1894.180 19.340 ;
        RECT 2054.460 19.760 2054.720 20.020 ;
      LAYER met2 ;
        RECT 1772.470 2006.155 1772.750 2006.525 ;
        RECT 1772.540 2001.230 1772.680 2006.155 ;
        RECT 1772.480 2000.910 1772.740 2001.230 ;
        RECT 1893.920 2000.910 1894.180 2001.230 ;
        RECT 1893.980 19.370 1894.120 2000.910 ;
        RECT 2054.460 19.730 2054.720 20.050 ;
        RECT 1893.920 19.050 1894.180 19.370 ;
        RECT 2054.520 2.400 2054.660 19.730 ;
        RECT 2054.310 -4.800 2054.870 2.400 ;
      LAYER via2 ;
        RECT 1772.470 2006.200 1772.750 2006.480 ;
      LAYER met3 ;
        RECT 1755.835 2006.490 1759.835 2006.495 ;
        RECT 1772.445 2006.490 1772.775 2006.505 ;
        RECT 1755.835 2006.190 1772.775 2006.490 ;
        RECT 1755.835 2005.895 1759.835 2006.190 ;
        RECT 1772.445 2006.175 1772.775 2006.190 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 686.925 1369.605 687.095 1393.575 ;
        RECT 717.285 1325.065 717.455 1337.475 ;
      LAYER mcon ;
        RECT 686.925 1393.405 687.095 1393.575 ;
        RECT 717.285 1337.305 717.455 1337.475 ;
      LAYER met1 ;
        RECT 686.850 2377.180 687.170 2377.240 ;
        RECT 898.910 2377.180 899.230 2377.240 ;
        RECT 686.850 2377.040 899.230 2377.180 ;
        RECT 686.850 2376.980 687.170 2377.040 ;
        RECT 898.910 2376.980 899.230 2377.040 ;
        RECT 686.850 1393.560 687.170 1393.620 ;
        RECT 686.655 1393.420 687.170 1393.560 ;
        RECT 686.850 1393.360 687.170 1393.420 ;
        RECT 686.850 1369.760 687.170 1369.820 ;
        RECT 686.655 1369.620 687.170 1369.760 ;
        RECT 686.850 1369.560 687.170 1369.620 ;
        RECT 686.850 1337.460 687.170 1337.520 ;
        RECT 717.225 1337.460 717.515 1337.505 ;
        RECT 686.850 1337.320 717.515 1337.460 ;
        RECT 686.850 1337.260 687.170 1337.320 ;
        RECT 717.225 1337.275 717.515 1337.320 ;
        RECT 717.225 1325.220 717.515 1325.265 ;
        RECT 766.430 1325.220 766.750 1325.280 ;
        RECT 717.225 1325.080 766.750 1325.220 ;
        RECT 717.225 1325.035 717.515 1325.080 ;
        RECT 766.430 1325.020 766.750 1325.080 ;
        RECT 766.430 20.300 766.750 20.360 ;
        RECT 769.650 20.300 769.970 20.360 ;
        RECT 766.430 20.160 769.970 20.300 ;
        RECT 766.430 20.100 766.750 20.160 ;
        RECT 769.650 20.100 769.970 20.160 ;
      LAYER via ;
        RECT 686.880 2376.980 687.140 2377.240 ;
        RECT 898.940 2376.980 899.200 2377.240 ;
        RECT 686.880 1393.360 687.140 1393.620 ;
        RECT 686.880 1369.560 687.140 1369.820 ;
        RECT 686.880 1337.260 687.140 1337.520 ;
        RECT 766.460 1325.020 766.720 1325.280 ;
        RECT 766.460 20.100 766.720 20.360 ;
        RECT 769.680 20.100 769.940 20.360 ;
      LAYER met2 ;
        RECT 686.880 2376.950 687.140 2377.270 ;
        RECT 898.940 2377.010 899.200 2377.270 ;
        RECT 900.820 2377.010 901.100 2377.880 ;
        RECT 898.940 2376.950 901.100 2377.010 ;
        RECT 686.940 1393.650 687.080 2376.950 ;
        RECT 899.000 2376.870 901.100 2376.950 ;
        RECT 900.820 2373.880 901.100 2376.870 ;
        RECT 686.880 1393.330 687.140 1393.650 ;
        RECT 686.880 1369.530 687.140 1369.850 ;
        RECT 686.940 1337.550 687.080 1369.530 ;
        RECT 686.880 1337.230 687.140 1337.550 ;
        RECT 766.460 1324.990 766.720 1325.310 ;
        RECT 766.520 20.390 766.660 1324.990 ;
        RECT 766.460 20.070 766.720 20.390 ;
        RECT 769.680 20.070 769.940 20.390 ;
        RECT 769.740 2.400 769.880 20.070 ;
        RECT 769.530 -4.800 770.090 2.400 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 713.145 1927.885 713.315 1947.095 ;
        RECT 713.605 1766.385 713.775 1798.855 ;
        RECT 713.605 1637.185 713.775 1653.335 ;
        RECT 718.205 1528.385 718.375 1572.415 ;
        RECT 2072.445 2.805 2072.615 48.195 ;
      LAYER mcon ;
        RECT 713.145 1946.925 713.315 1947.095 ;
        RECT 713.605 1798.685 713.775 1798.855 ;
        RECT 713.605 1653.165 713.775 1653.335 ;
        RECT 718.205 1572.245 718.375 1572.415 ;
        RECT 2072.445 48.025 2072.615 48.195 ;
      LAYER met1 ;
        RECT 717.210 2218.400 717.530 2218.460 ;
        RECT 719.050 2218.400 719.370 2218.460 ;
        RECT 717.210 2218.260 719.370 2218.400 ;
        RECT 717.210 2218.200 717.530 2218.260 ;
        RECT 719.050 2218.200 719.370 2218.260 ;
        RECT 713.070 1947.080 713.390 1947.140 ;
        RECT 712.875 1946.940 713.390 1947.080 ;
        RECT 713.070 1946.880 713.390 1946.940 ;
        RECT 713.085 1928.040 713.375 1928.085 ;
        RECT 718.590 1928.040 718.910 1928.100 ;
        RECT 713.085 1927.900 718.910 1928.040 ;
        RECT 713.085 1927.855 713.375 1927.900 ;
        RECT 718.590 1927.840 718.910 1927.900 ;
        RECT 717.670 1885.880 717.990 1885.940 ;
        RECT 718.590 1885.880 718.910 1885.940 ;
        RECT 717.670 1885.740 718.910 1885.880 ;
        RECT 717.670 1885.680 717.990 1885.740 ;
        RECT 718.590 1885.680 718.910 1885.740 ;
        RECT 713.990 1857.320 714.310 1857.380 ;
        RECT 717.670 1857.320 717.990 1857.380 ;
        RECT 713.990 1857.180 717.990 1857.320 ;
        RECT 713.990 1857.120 714.310 1857.180 ;
        RECT 717.670 1857.120 717.990 1857.180 ;
        RECT 713.545 1798.840 713.835 1798.885 ;
        RECT 713.990 1798.840 714.310 1798.900 ;
        RECT 713.545 1798.700 714.310 1798.840 ;
        RECT 713.545 1798.655 713.835 1798.700 ;
        RECT 713.990 1798.640 714.310 1798.700 ;
        RECT 713.530 1766.540 713.850 1766.600 ;
        RECT 713.335 1766.400 713.850 1766.540 ;
        RECT 713.530 1766.340 713.850 1766.400 ;
        RECT 713.530 1653.320 713.850 1653.380 ;
        RECT 713.335 1653.180 713.850 1653.320 ;
        RECT 713.530 1653.120 713.850 1653.180 ;
        RECT 713.545 1637.340 713.835 1637.385 ;
        RECT 713.990 1637.340 714.310 1637.400 ;
        RECT 713.545 1637.200 714.310 1637.340 ;
        RECT 713.545 1637.155 713.835 1637.200 ;
        RECT 713.990 1637.140 714.310 1637.200 ;
        RECT 718.145 1572.400 718.435 1572.445 ;
        RECT 718.590 1572.400 718.910 1572.460 ;
        RECT 718.145 1572.260 718.910 1572.400 ;
        RECT 718.145 1572.215 718.435 1572.260 ;
        RECT 718.590 1572.200 718.910 1572.260 ;
        RECT 718.145 1528.540 718.435 1528.585 ;
        RECT 718.590 1528.540 718.910 1528.600 ;
        RECT 718.145 1528.400 718.910 1528.540 ;
        RECT 718.145 1528.355 718.435 1528.400 ;
        RECT 718.590 1528.340 718.910 1528.400 ;
        RECT 711.690 1480.260 712.010 1480.320 ;
        RECT 718.590 1480.260 718.910 1480.320 ;
        RECT 711.690 1480.120 718.910 1480.260 ;
        RECT 711.690 1480.060 712.010 1480.120 ;
        RECT 718.590 1480.060 718.910 1480.120 ;
        RECT 2070.070 48.180 2070.390 48.240 ;
        RECT 2072.385 48.180 2072.675 48.225 ;
        RECT 2070.070 48.040 2072.675 48.180 ;
        RECT 2070.070 47.980 2070.390 48.040 ;
        RECT 2072.385 47.995 2072.675 48.040 ;
        RECT 2072.370 2.960 2072.690 3.020 ;
        RECT 2072.175 2.820 2072.690 2.960 ;
        RECT 2072.370 2.760 2072.690 2.820 ;
      LAYER via ;
        RECT 717.240 2218.200 717.500 2218.460 ;
        RECT 719.080 2218.200 719.340 2218.460 ;
        RECT 713.100 1946.880 713.360 1947.140 ;
        RECT 718.620 1927.840 718.880 1928.100 ;
        RECT 717.700 1885.680 717.960 1885.940 ;
        RECT 718.620 1885.680 718.880 1885.940 ;
        RECT 714.020 1857.120 714.280 1857.380 ;
        RECT 717.700 1857.120 717.960 1857.380 ;
        RECT 714.020 1798.640 714.280 1798.900 ;
        RECT 713.560 1766.340 713.820 1766.600 ;
        RECT 713.560 1653.120 713.820 1653.380 ;
        RECT 714.020 1637.140 714.280 1637.400 ;
        RECT 718.620 1572.200 718.880 1572.460 ;
        RECT 718.620 1528.340 718.880 1528.600 ;
        RECT 711.720 1480.060 711.980 1480.320 ;
        RECT 718.620 1480.060 718.880 1480.320 ;
        RECT 2070.100 47.980 2070.360 48.240 ;
        RECT 2072.400 2.760 2072.660 3.020 ;
      LAYER met2 ;
        RECT 717.230 2242.795 717.510 2243.165 ;
        RECT 717.300 2218.490 717.440 2242.795 ;
        RECT 717.240 2218.170 717.500 2218.490 ;
        RECT 719.080 2218.170 719.340 2218.490 ;
        RECT 719.140 2160.205 719.280 2218.170 ;
        RECT 719.070 2159.835 719.350 2160.205 ;
        RECT 718.150 2144.195 718.430 2144.565 ;
        RECT 718.220 2128.245 718.360 2144.195 ;
        RECT 718.150 2127.875 718.430 2128.245 ;
        RECT 718.610 2100.675 718.890 2101.045 ;
        RECT 718.680 2084.725 718.820 2100.675 ;
        RECT 718.610 2084.355 718.890 2084.725 ;
        RECT 717.690 2073.475 717.970 2073.845 ;
        RECT 717.760 1990.885 717.900 2073.475 ;
        RECT 717.690 1990.515 717.970 1990.885 ;
        RECT 713.090 1960.595 713.370 1960.965 ;
        RECT 713.160 1947.170 713.300 1960.595 ;
        RECT 713.100 1946.850 713.360 1947.170 ;
        RECT 718.620 1927.810 718.880 1928.130 ;
        RECT 718.680 1885.970 718.820 1927.810 ;
        RECT 717.700 1885.650 717.960 1885.970 ;
        RECT 718.620 1885.650 718.880 1885.970 ;
        RECT 717.760 1857.410 717.900 1885.650 ;
        RECT 714.020 1857.090 714.280 1857.410 ;
        RECT 717.700 1857.090 717.960 1857.410 ;
        RECT 714.080 1798.930 714.220 1857.090 ;
        RECT 714.020 1798.610 714.280 1798.930 ;
        RECT 713.560 1766.310 713.820 1766.630 ;
        RECT 713.620 1653.410 713.760 1766.310 ;
        RECT 713.560 1653.090 713.820 1653.410 ;
        RECT 714.020 1637.110 714.280 1637.430 ;
        RECT 714.080 1576.085 714.220 1637.110 ;
        RECT 714.010 1575.715 714.290 1576.085 ;
        RECT 718.610 1572.315 718.890 1572.685 ;
        RECT 718.620 1572.170 718.880 1572.315 ;
        RECT 718.620 1528.310 718.880 1528.630 ;
        RECT 718.680 1480.350 718.820 1528.310 ;
        RECT 711.720 1480.030 711.980 1480.350 ;
        RECT 718.620 1480.030 718.880 1480.350 ;
        RECT 711.780 1467.285 711.920 1480.030 ;
        RECT 711.710 1466.915 711.990 1467.285 ;
        RECT 704.810 1388.715 705.090 1389.085 ;
        RECT 704.880 1346.925 705.020 1388.715 ;
        RECT 704.810 1346.555 705.090 1346.925 ;
        RECT 721.830 654.995 722.110 655.365 ;
        RECT 721.900 631.565 722.040 654.995 ;
        RECT 721.830 631.195 722.110 631.565 ;
        RECT 2070.090 72.915 2070.370 73.285 ;
        RECT 2070.160 48.270 2070.300 72.915 ;
        RECT 2070.100 47.950 2070.360 48.270 ;
        RECT 2072.400 2.730 2072.660 3.050 ;
        RECT 2072.460 2.400 2072.600 2.730 ;
        RECT 2072.250 -4.800 2072.810 2.400 ;
      LAYER via2 ;
        RECT 717.230 2242.840 717.510 2243.120 ;
        RECT 719.070 2159.880 719.350 2160.160 ;
        RECT 718.150 2144.240 718.430 2144.520 ;
        RECT 718.150 2127.920 718.430 2128.200 ;
        RECT 718.610 2100.720 718.890 2101.000 ;
        RECT 718.610 2084.400 718.890 2084.680 ;
        RECT 717.690 2073.520 717.970 2073.800 ;
        RECT 717.690 1990.560 717.970 1990.840 ;
        RECT 713.090 1960.640 713.370 1960.920 ;
        RECT 714.010 1575.760 714.290 1576.040 ;
        RECT 718.610 1572.360 718.890 1572.640 ;
        RECT 711.710 1466.960 711.990 1467.240 ;
        RECT 704.810 1388.760 705.090 1389.040 ;
        RECT 704.810 1346.600 705.090 1346.880 ;
        RECT 721.830 655.040 722.110 655.320 ;
        RECT 721.830 631.240 722.110 631.520 ;
        RECT 2070.090 72.960 2070.370 73.240 ;
      LAYER met3 ;
        RECT 715.810 2284.695 719.810 2285.295 ;
        RECT 718.830 2282.580 719.130 2284.695 ;
        RECT 718.790 2282.260 719.170 2282.580 ;
        RECT 717.205 2243.130 717.535 2243.145 ;
        RECT 718.790 2243.130 719.170 2243.140 ;
        RECT 717.205 2242.830 719.170 2243.130 ;
        RECT 717.205 2242.815 717.535 2242.830 ;
        RECT 718.790 2242.820 719.170 2242.830 ;
        RECT 719.045 2160.180 719.375 2160.185 ;
        RECT 718.790 2160.170 719.375 2160.180 ;
        RECT 718.590 2159.870 719.375 2160.170 ;
        RECT 718.790 2159.860 719.375 2159.870 ;
        RECT 719.045 2159.855 719.375 2159.860 ;
        RECT 718.125 2144.530 718.455 2144.545 ;
        RECT 718.790 2144.530 719.170 2144.540 ;
        RECT 718.125 2144.230 719.170 2144.530 ;
        RECT 718.125 2144.215 718.455 2144.230 ;
        RECT 718.790 2144.220 719.170 2144.230 ;
        RECT 718.125 2128.210 718.455 2128.225 ;
        RECT 718.790 2128.210 719.170 2128.220 ;
        RECT 718.125 2127.910 719.170 2128.210 ;
        RECT 718.125 2127.895 718.455 2127.910 ;
        RECT 718.790 2127.900 719.170 2127.910 ;
        RECT 718.585 2101.020 718.915 2101.025 ;
        RECT 718.585 2101.010 719.170 2101.020 ;
        RECT 718.360 2100.710 719.170 2101.010 ;
        RECT 718.585 2100.700 719.170 2100.710 ;
        RECT 718.585 2100.695 718.915 2100.700 ;
        RECT 718.585 2084.700 718.915 2084.705 ;
        RECT 718.585 2084.690 719.170 2084.700 ;
        RECT 718.360 2084.390 719.170 2084.690 ;
        RECT 718.585 2084.380 719.170 2084.390 ;
        RECT 718.585 2084.375 718.915 2084.380 ;
        RECT 717.665 2073.810 717.995 2073.825 ;
        RECT 718.790 2073.810 719.170 2073.820 ;
        RECT 717.665 2073.510 719.170 2073.810 ;
        RECT 717.665 2073.495 717.995 2073.510 ;
        RECT 718.790 2073.500 719.170 2073.510 ;
        RECT 717.665 1990.850 717.995 1990.865 ;
        RECT 718.790 1990.850 719.170 1990.860 ;
        RECT 717.665 1990.550 719.170 1990.850 ;
        RECT 717.665 1990.535 717.995 1990.550 ;
        RECT 718.790 1990.540 719.170 1990.550 ;
        RECT 713.065 1960.930 713.395 1960.945 ;
        RECT 718.790 1960.930 719.170 1960.940 ;
        RECT 713.065 1960.630 719.170 1960.930 ;
        RECT 713.065 1960.615 713.395 1960.630 ;
        RECT 718.790 1960.620 719.170 1960.630 ;
        RECT 713.985 1576.050 714.315 1576.065 ;
        RECT 718.790 1576.050 719.170 1576.060 ;
        RECT 713.985 1575.750 719.170 1576.050 ;
        RECT 713.985 1575.735 714.315 1575.750 ;
        RECT 718.790 1575.740 719.170 1575.750 ;
        RECT 718.585 1572.660 718.915 1572.665 ;
        RECT 718.585 1572.650 719.170 1572.660 ;
        RECT 718.585 1572.350 719.370 1572.650 ;
        RECT 718.585 1572.340 719.170 1572.350 ;
        RECT 718.585 1572.335 718.915 1572.340 ;
        RECT 711.685 1467.250 712.015 1467.265 ;
        RECT 718.790 1467.250 719.170 1467.260 ;
        RECT 711.685 1466.950 719.170 1467.250 ;
        RECT 711.685 1466.935 712.015 1466.950 ;
        RECT 718.790 1466.940 719.170 1466.950 ;
        RECT 704.785 1389.050 705.115 1389.065 ;
        RECT 718.790 1389.050 719.170 1389.060 ;
        RECT 704.785 1388.750 719.170 1389.050 ;
        RECT 704.785 1388.735 705.115 1388.750 ;
        RECT 718.790 1388.740 719.170 1388.750 ;
        RECT 704.785 1346.890 705.115 1346.905 ;
        RECT 717.870 1346.890 718.250 1346.900 ;
        RECT 704.785 1346.590 718.250 1346.890 ;
        RECT 704.785 1346.575 705.115 1346.590 ;
        RECT 717.870 1346.580 718.250 1346.590 ;
        RECT 721.805 655.340 722.135 655.345 ;
        RECT 721.550 655.330 722.135 655.340 ;
        RECT 721.550 655.030 722.360 655.330 ;
        RECT 721.550 655.020 722.135 655.030 ;
        RECT 721.805 655.015 722.135 655.020 ;
        RECT 721.805 631.540 722.135 631.545 ;
        RECT 721.550 631.530 722.135 631.540 ;
        RECT 721.350 631.230 722.135 631.530 ;
        RECT 721.550 631.220 722.135 631.230 ;
        RECT 721.805 631.215 722.135 631.220 ;
        RECT 721.550 73.250 721.930 73.260 ;
        RECT 2070.065 73.250 2070.395 73.265 ;
        RECT 721.550 72.950 2070.395 73.250 ;
        RECT 721.550 72.940 721.930 72.950 ;
        RECT 2070.065 72.935 2070.395 72.950 ;
      LAYER via3 ;
        RECT 718.820 2282.260 719.140 2282.580 ;
        RECT 718.820 2242.820 719.140 2243.140 ;
        RECT 718.820 2159.860 719.140 2160.180 ;
        RECT 718.820 2144.220 719.140 2144.540 ;
        RECT 718.820 2127.900 719.140 2128.220 ;
        RECT 718.820 2100.700 719.140 2101.020 ;
        RECT 718.820 2084.380 719.140 2084.700 ;
        RECT 718.820 2073.500 719.140 2073.820 ;
        RECT 718.820 1990.540 719.140 1990.860 ;
        RECT 718.820 1960.620 719.140 1960.940 ;
        RECT 718.820 1575.740 719.140 1576.060 ;
        RECT 718.820 1572.340 719.140 1572.660 ;
        RECT 718.820 1466.940 719.140 1467.260 ;
        RECT 718.820 1388.740 719.140 1389.060 ;
        RECT 717.900 1346.580 718.220 1346.900 ;
        RECT 721.580 655.020 721.900 655.340 ;
        RECT 721.580 631.220 721.900 631.540 ;
        RECT 721.580 72.940 721.900 73.260 ;
      LAYER met4 ;
        RECT 718.815 2282.255 719.145 2282.585 ;
        RECT 718.830 2243.145 719.130 2282.255 ;
        RECT 718.815 2242.815 719.145 2243.145 ;
        RECT 718.815 2159.855 719.145 2160.185 ;
        RECT 718.830 2144.545 719.130 2159.855 ;
        RECT 718.815 2144.215 719.145 2144.545 ;
        RECT 718.815 2127.895 719.145 2128.225 ;
        RECT 718.830 2101.025 719.130 2127.895 ;
        RECT 718.815 2100.695 719.145 2101.025 ;
        RECT 718.815 2084.375 719.145 2084.705 ;
        RECT 718.830 2073.825 719.130 2084.375 ;
        RECT 718.815 2073.495 719.145 2073.825 ;
        RECT 718.815 1990.850 719.145 1990.865 ;
        RECT 718.815 1990.550 720.050 1990.850 ;
        RECT 718.815 1990.535 719.145 1990.550 ;
        RECT 719.750 1962.970 720.050 1990.550 ;
        RECT 718.830 1962.670 720.050 1962.970 ;
        RECT 718.830 1960.945 719.130 1962.670 ;
        RECT 718.815 1960.615 719.145 1960.945 ;
        RECT 718.815 1576.050 719.145 1576.065 ;
        RECT 718.815 1575.750 720.970 1576.050 ;
        RECT 718.815 1575.735 719.145 1575.750 ;
        RECT 718.815 1572.650 719.145 1572.665 ;
        RECT 720.670 1572.650 720.970 1575.750 ;
        RECT 718.815 1572.350 720.970 1572.650 ;
        RECT 718.815 1572.335 719.145 1572.350 ;
        RECT 718.815 1467.250 719.145 1467.265 ;
        RECT 718.815 1466.950 720.050 1467.250 ;
        RECT 718.815 1466.935 719.145 1466.950 ;
        RECT 719.750 1466.570 720.050 1466.950 ;
        RECT 719.750 1466.270 721.890 1466.570 ;
        RECT 721.590 1452.970 721.890 1466.270 ;
        RECT 720.670 1452.670 721.890 1452.970 ;
        RECT 720.670 1433.690 720.970 1452.670 ;
        RECT 720.230 1432.510 721.410 1433.690 ;
        RECT 719.310 1401.910 720.490 1403.090 ;
        RECT 718.815 1389.050 719.145 1389.065 ;
        RECT 719.750 1389.050 720.050 1401.910 ;
        RECT 718.815 1388.750 720.050 1389.050 ;
        RECT 718.815 1388.735 719.145 1388.750 ;
        RECT 717.910 1347.950 721.890 1348.250 ;
        RECT 717.910 1346.905 718.210 1347.950 ;
        RECT 717.895 1346.575 718.225 1346.905 ;
        RECT 721.590 655.345 721.890 1347.950 ;
        RECT 721.575 655.015 721.905 655.345 ;
        RECT 721.575 631.215 721.905 631.545 ;
        RECT 721.590 73.265 721.890 631.215 ;
        RECT 721.575 72.935 721.905 73.265 ;
      LAYER met5 ;
        RECT 718.180 1432.300 721.620 1433.900 ;
        RECT 718.180 1430.500 719.780 1432.300 ;
        RECT 717.260 1428.900 719.780 1430.500 ;
        RECT 717.260 1403.300 718.860 1428.900 ;
        RECT 717.260 1401.700 720.700 1403.300 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 790.370 2381.515 790.650 2381.885 ;
        RECT 790.440 2377.880 790.580 2381.515 ;
        RECT 790.420 2373.880 790.700 2377.880 ;
        RECT 2089.870 19.875 2090.150 20.245 ;
        RECT 2089.940 2.400 2090.080 19.875 ;
        RECT 2089.730 -4.800 2090.290 2.400 ;
      LAYER via2 ;
        RECT 790.370 2381.560 790.650 2381.840 ;
        RECT 2089.870 19.920 2090.150 20.200 ;
      LAYER met3 ;
        RECT 790.345 2381.850 790.675 2381.865 ;
        RECT 1748.270 2381.850 1748.650 2381.860 ;
        RECT 790.345 2381.550 1748.650 2381.850 ;
        RECT 790.345 2381.535 790.675 2381.550 ;
        RECT 1748.270 2381.540 1748.650 2381.550 ;
        RECT 1748.270 20.210 1748.650 20.220 ;
        RECT 2089.845 20.210 2090.175 20.225 ;
        RECT 1748.270 19.910 2090.175 20.210 ;
        RECT 1748.270 19.900 1748.650 19.910 ;
        RECT 2089.845 19.895 2090.175 19.910 ;
      LAYER via3 ;
        RECT 1748.300 2381.540 1748.620 2381.860 ;
        RECT 1748.300 19.900 1748.620 20.220 ;
      LAYER met4 ;
        RECT 1748.295 2381.535 1748.625 2381.865 ;
        RECT 1748.310 20.225 1748.610 2381.535 ;
        RECT 1748.295 19.895 1748.625 20.225 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1772.910 1462.920 1773.230 1462.980 ;
        RECT 2087.090 1462.920 2087.410 1462.980 ;
        RECT 1772.910 1462.780 2087.410 1462.920 ;
        RECT 1772.910 1462.720 1773.230 1462.780 ;
        RECT 2087.090 1462.720 2087.410 1462.780 ;
        RECT 2087.090 20.300 2087.410 20.360 ;
        RECT 2107.790 20.300 2108.110 20.360 ;
        RECT 2087.090 20.160 2108.110 20.300 ;
        RECT 2087.090 20.100 2087.410 20.160 ;
        RECT 2107.790 20.100 2108.110 20.160 ;
      LAYER via ;
        RECT 1772.940 1462.720 1773.200 1462.980 ;
        RECT 2087.120 1462.720 2087.380 1462.980 ;
        RECT 2087.120 20.100 2087.380 20.360 ;
        RECT 2107.820 20.100 2108.080 20.360 ;
      LAYER met2 ;
        RECT 1772.930 1467.595 1773.210 1467.965 ;
        RECT 1773.000 1463.010 1773.140 1467.595 ;
        RECT 1772.940 1462.690 1773.200 1463.010 ;
        RECT 2087.120 1462.690 2087.380 1463.010 ;
        RECT 2087.180 20.390 2087.320 1462.690 ;
        RECT 2087.120 20.070 2087.380 20.390 ;
        RECT 2107.820 20.070 2108.080 20.390 ;
        RECT 2107.880 2.400 2108.020 20.070 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
      LAYER via2 ;
        RECT 1772.930 1467.640 1773.210 1467.920 ;
      LAYER met3 ;
        RECT 1755.835 1467.930 1759.835 1467.935 ;
        RECT 1772.905 1467.930 1773.235 1467.945 ;
        RECT 1755.835 1467.630 1773.235 1467.930 ;
        RECT 1755.835 1467.335 1759.835 1467.630 ;
        RECT 1772.905 1467.615 1773.235 1467.630 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1346.030 2391.460 1346.350 2391.520 ;
        RECT 1758.190 2391.460 1758.510 2391.520 ;
        RECT 1346.030 2391.320 1758.510 2391.460 ;
        RECT 1346.030 2391.260 1346.350 2391.320 ;
        RECT 1758.190 2391.260 1758.510 2391.320 ;
        RECT 1758.190 2321.760 1758.510 2321.820 ;
        RECT 2125.270 2321.760 2125.590 2321.820 ;
        RECT 1758.190 2321.620 2125.590 2321.760 ;
        RECT 1758.190 2321.560 1758.510 2321.620 ;
        RECT 2125.270 2321.560 2125.590 2321.620 ;
      LAYER via ;
        RECT 1346.060 2391.260 1346.320 2391.520 ;
        RECT 1758.220 2391.260 1758.480 2391.520 ;
        RECT 1758.220 2321.560 1758.480 2321.820 ;
        RECT 2125.300 2321.560 2125.560 2321.820 ;
      LAYER met2 ;
        RECT 1346.060 2391.230 1346.320 2391.550 ;
        RECT 1758.220 2391.230 1758.480 2391.550 ;
        RECT 1346.120 2377.880 1346.260 2391.230 ;
        RECT 1346.100 2373.880 1346.380 2377.880 ;
        RECT 1758.280 2321.850 1758.420 2391.230 ;
        RECT 1758.220 2321.530 1758.480 2321.850 ;
        RECT 2125.300 2321.530 2125.560 2321.850 ;
        RECT 2125.360 17.410 2125.500 2321.530 ;
        RECT 2125.360 17.270 2125.960 17.410 ;
        RECT 2125.820 2.400 2125.960 17.270 ;
        RECT 2125.610 -4.800 2126.170 2.400 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 708.010 72.320 708.330 72.380 ;
        RECT 2139.070 72.320 2139.390 72.380 ;
        RECT 708.010 72.180 2139.390 72.320 ;
        RECT 708.010 72.120 708.330 72.180 ;
        RECT 2139.070 72.120 2139.390 72.180 ;
      LAYER via ;
        RECT 708.040 72.120 708.300 72.380 ;
        RECT 2139.100 72.120 2139.360 72.380 ;
      LAYER met2 ;
        RECT 708.030 1507.035 708.310 1507.405 ;
        RECT 708.100 72.410 708.240 1507.035 ;
        RECT 708.040 72.090 708.300 72.410 ;
        RECT 2139.100 72.090 2139.360 72.410 ;
        RECT 2139.160 16.730 2139.300 72.090 ;
        RECT 2139.160 16.590 2143.900 16.730 ;
        RECT 2143.760 2.400 2143.900 16.590 ;
        RECT 2143.550 -4.800 2144.110 2.400 ;
      LAYER via2 ;
        RECT 708.030 1507.080 708.310 1507.360 ;
      LAYER met3 ;
        RECT 708.005 1507.370 708.335 1507.385 ;
        RECT 715.810 1507.370 719.810 1507.375 ;
        RECT 708.005 1507.070 719.810 1507.370 ;
        RECT 708.005 1507.055 708.335 1507.070 ;
        RECT 715.810 1506.775 719.810 1507.070 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1772.910 1608.100 1773.230 1608.160 ;
        RECT 2045.690 1608.100 2046.010 1608.160 ;
        RECT 1772.910 1607.960 2046.010 1608.100 ;
        RECT 1772.910 1607.900 1773.230 1607.960 ;
        RECT 2045.690 1607.900 2046.010 1607.960 ;
        RECT 2045.690 19.620 2046.010 19.680 ;
        RECT 2161.610 19.620 2161.930 19.680 ;
        RECT 2045.690 19.480 2161.930 19.620 ;
        RECT 2045.690 19.420 2046.010 19.480 ;
        RECT 2161.610 19.420 2161.930 19.480 ;
      LAYER via ;
        RECT 1772.940 1607.900 1773.200 1608.160 ;
        RECT 2045.720 1607.900 2045.980 1608.160 ;
        RECT 2045.720 19.420 2045.980 19.680 ;
        RECT 2161.640 19.420 2161.900 19.680 ;
      LAYER met2 ;
        RECT 1772.930 1613.115 1773.210 1613.485 ;
        RECT 1773.000 1608.190 1773.140 1613.115 ;
        RECT 1772.940 1607.870 1773.200 1608.190 ;
        RECT 2045.720 1607.870 2045.980 1608.190 ;
        RECT 2045.780 19.710 2045.920 1607.870 ;
        RECT 2045.720 19.390 2045.980 19.710 ;
        RECT 2161.640 19.390 2161.900 19.710 ;
        RECT 2161.700 2.400 2161.840 19.390 ;
        RECT 2161.490 -4.800 2162.050 2.400 ;
      LAYER via2 ;
        RECT 1772.930 1613.160 1773.210 1613.440 ;
      LAYER met3 ;
        RECT 1755.835 1613.450 1759.835 1613.455 ;
        RECT 1772.905 1613.450 1773.235 1613.465 ;
        RECT 1755.835 1613.150 1773.235 1613.450 ;
        RECT 1755.835 1612.855 1759.835 1613.150 ;
        RECT 1772.905 1613.135 1773.235 1613.150 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1771.990 2166.720 1772.310 2166.780 ;
        RECT 2162.990 2166.720 2163.310 2166.780 ;
        RECT 1771.990 2166.580 2163.310 2166.720 ;
        RECT 1771.990 2166.520 1772.310 2166.580 ;
        RECT 2162.990 2166.520 2163.310 2166.580 ;
        RECT 2162.990 19.620 2163.310 19.680 ;
        RECT 2179.090 19.620 2179.410 19.680 ;
        RECT 2162.990 19.480 2179.410 19.620 ;
        RECT 2162.990 19.420 2163.310 19.480 ;
        RECT 2179.090 19.420 2179.410 19.480 ;
      LAYER via ;
        RECT 1772.020 2166.520 1772.280 2166.780 ;
        RECT 2163.020 2166.520 2163.280 2166.780 ;
        RECT 2163.020 19.420 2163.280 19.680 ;
        RECT 2179.120 19.420 2179.380 19.680 ;
      LAYER met2 ;
        RECT 1772.010 2169.355 1772.290 2169.725 ;
        RECT 1772.080 2166.810 1772.220 2169.355 ;
        RECT 1772.020 2166.490 1772.280 2166.810 ;
        RECT 2163.020 2166.490 2163.280 2166.810 ;
        RECT 2163.080 19.710 2163.220 2166.490 ;
        RECT 2163.020 19.390 2163.280 19.710 ;
        RECT 2179.120 19.390 2179.380 19.710 ;
        RECT 2179.180 2.400 2179.320 19.390 ;
        RECT 2178.970 -4.800 2179.530 2.400 ;
      LAYER via2 ;
        RECT 1772.010 2169.400 1772.290 2169.680 ;
      LAYER met3 ;
        RECT 1755.835 2169.690 1759.835 2169.695 ;
        RECT 1771.985 2169.690 1772.315 2169.705 ;
        RECT 1755.835 2169.390 1772.315 2169.690 ;
        RECT 1755.835 2169.095 1759.835 2169.390 ;
        RECT 1771.985 2169.375 1772.315 2169.390 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1715.870 2388.400 1716.190 2388.460 ;
        RECT 2176.790 2388.400 2177.110 2388.460 ;
        RECT 1715.870 2388.260 2177.110 2388.400 ;
        RECT 1715.870 2388.200 1716.190 2388.260 ;
        RECT 2176.790 2388.200 2177.110 2388.260 ;
        RECT 2176.790 20.300 2177.110 20.360 ;
        RECT 2197.030 20.300 2197.350 20.360 ;
        RECT 2176.790 20.160 2197.350 20.300 ;
        RECT 2176.790 20.100 2177.110 20.160 ;
        RECT 2197.030 20.100 2197.350 20.160 ;
      LAYER via ;
        RECT 1715.900 2388.200 1716.160 2388.460 ;
        RECT 2176.820 2388.200 2177.080 2388.460 ;
        RECT 2176.820 20.100 2177.080 20.360 ;
        RECT 2197.060 20.100 2197.320 20.360 ;
      LAYER met2 ;
        RECT 1715.900 2388.170 1716.160 2388.490 ;
        RECT 2176.820 2388.170 2177.080 2388.490 ;
        RECT 1715.960 2377.880 1716.100 2388.170 ;
        RECT 1715.940 2373.880 1716.220 2377.880 ;
        RECT 2176.880 20.390 2177.020 2388.170 ;
        RECT 2176.820 20.070 2177.080 20.390 ;
        RECT 2197.060 20.070 2197.320 20.390 ;
        RECT 2197.120 2.400 2197.260 20.070 ;
        RECT 2196.910 -4.800 2197.470 2.400 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1768.310 1380.300 1768.630 1380.360 ;
        RECT 2197.490 1380.300 2197.810 1380.360 ;
        RECT 1768.310 1380.160 2197.810 1380.300 ;
        RECT 1768.310 1380.100 1768.630 1380.160 ;
        RECT 2197.490 1380.100 2197.810 1380.160 ;
        RECT 2197.490 20.640 2197.810 20.700 ;
        RECT 2214.970 20.640 2215.290 20.700 ;
        RECT 2197.490 20.500 2215.290 20.640 ;
        RECT 2197.490 20.440 2197.810 20.500 ;
        RECT 2214.970 20.440 2215.290 20.500 ;
      LAYER via ;
        RECT 1768.340 1380.100 1768.600 1380.360 ;
        RECT 2197.520 1380.100 2197.780 1380.360 ;
        RECT 2197.520 20.440 2197.780 20.700 ;
        RECT 2215.000 20.440 2215.260 20.700 ;
      LAYER met2 ;
        RECT 1768.330 1381.915 1768.610 1382.285 ;
        RECT 1768.400 1380.390 1768.540 1381.915 ;
        RECT 1768.340 1380.070 1768.600 1380.390 ;
        RECT 2197.520 1380.070 2197.780 1380.390 ;
        RECT 2197.580 20.730 2197.720 1380.070 ;
        RECT 2197.520 20.410 2197.780 20.730 ;
        RECT 2215.000 20.410 2215.260 20.730 ;
        RECT 2215.060 2.400 2215.200 20.410 ;
        RECT 2214.850 -4.800 2215.410 2.400 ;
      LAYER via2 ;
        RECT 1768.330 1381.960 1768.610 1382.240 ;
      LAYER met3 ;
        RECT 1755.835 1382.250 1759.835 1382.255 ;
        RECT 1768.305 1382.250 1768.635 1382.265 ;
        RECT 1755.835 1381.950 1768.635 1382.250 ;
        RECT 1755.835 1381.655 1759.835 1381.950 ;
        RECT 1768.305 1381.935 1768.635 1381.950 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2228.790 154.515 2229.070 154.885 ;
        RECT 2228.860 16.730 2229.000 154.515 ;
        RECT 2228.860 16.590 2233.140 16.730 ;
        RECT 2233.000 2.400 2233.140 16.590 ;
        RECT 2232.790 -4.800 2233.350 2.400 ;
      LAYER via2 ;
        RECT 2228.790 154.560 2229.070 154.840 ;
      LAYER met3 ;
        RECT 699.470 2071.770 699.850 2071.780 ;
        RECT 715.810 2071.770 719.810 2071.775 ;
        RECT 699.470 2071.470 719.810 2071.770 ;
        RECT 699.470 2071.460 699.850 2071.470 ;
        RECT 715.810 2071.175 719.810 2071.470 ;
        RECT 699.470 154.850 699.850 154.860 ;
        RECT 2228.765 154.850 2229.095 154.865 ;
        RECT 699.470 154.550 2229.095 154.850 ;
        RECT 699.470 154.540 699.850 154.550 ;
        RECT 2228.765 154.535 2229.095 154.550 ;
      LAYER via3 ;
        RECT 699.500 2071.460 699.820 2071.780 ;
        RECT 699.500 154.540 699.820 154.860 ;
      LAYER met4 ;
        RECT 699.495 2071.455 699.825 2071.785 ;
        RECT 699.510 154.865 699.810 2071.455 ;
        RECT 699.495 154.535 699.825 154.865 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 793.110 1301.080 793.430 1301.140 ;
        RECT 1762.790 1301.080 1763.110 1301.140 ;
        RECT 793.110 1300.940 1763.110 1301.080 ;
        RECT 793.110 1300.880 793.430 1300.940 ;
        RECT 1762.790 1300.880 1763.110 1300.940 ;
        RECT 787.590 20.640 787.910 20.700 ;
        RECT 793.110 20.640 793.430 20.700 ;
        RECT 787.590 20.500 793.430 20.640 ;
        RECT 787.590 20.440 787.910 20.500 ;
        RECT 793.110 20.440 793.430 20.500 ;
      LAYER via ;
        RECT 793.140 1300.880 793.400 1301.140 ;
        RECT 1762.820 1300.880 1763.080 1301.140 ;
        RECT 787.620 20.440 787.880 20.700 ;
        RECT 793.140 20.440 793.400 20.700 ;
      LAYER met2 ;
        RECT 1762.810 1347.915 1763.090 1348.285 ;
        RECT 1762.880 1301.170 1763.020 1347.915 ;
        RECT 793.140 1300.850 793.400 1301.170 ;
        RECT 1762.820 1300.850 1763.080 1301.170 ;
        RECT 793.200 20.730 793.340 1300.850 ;
        RECT 787.620 20.410 787.880 20.730 ;
        RECT 793.140 20.410 793.400 20.730 ;
        RECT 787.680 2.400 787.820 20.410 ;
        RECT 787.470 -4.800 788.030 2.400 ;
      LAYER via2 ;
        RECT 1762.810 1347.960 1763.090 1348.240 ;
      LAYER met3 ;
        RECT 1755.835 1348.250 1759.835 1348.255 ;
        RECT 1762.785 1348.250 1763.115 1348.265 ;
        RECT 1755.835 1347.950 1763.115 1348.250 ;
        RECT 1755.835 1347.655 1759.835 1347.950 ;
        RECT 1762.785 1347.935 1763.115 1347.950 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1143.630 2392.140 1143.950 2392.200 ;
        RECT 1634.910 2392.140 1635.230 2392.200 ;
        RECT 1143.630 2392.000 1635.230 2392.140 ;
        RECT 1143.630 2391.940 1143.950 2392.000 ;
        RECT 1634.910 2391.940 1635.230 2392.000 ;
        RECT 1634.910 2385.680 1635.230 2385.740 ;
        RECT 2249.470 2385.680 2249.790 2385.740 ;
        RECT 1634.910 2385.540 2249.790 2385.680 ;
        RECT 1634.910 2385.480 1635.230 2385.540 ;
        RECT 2249.470 2385.480 2249.790 2385.540 ;
      LAYER via ;
        RECT 1143.660 2391.940 1143.920 2392.200 ;
        RECT 1634.940 2391.940 1635.200 2392.200 ;
        RECT 1634.940 2385.480 1635.200 2385.740 ;
        RECT 2249.500 2385.480 2249.760 2385.740 ;
      LAYER met2 ;
        RECT 1143.660 2391.910 1143.920 2392.230 ;
        RECT 1634.940 2391.910 1635.200 2392.230 ;
        RECT 1143.720 2377.880 1143.860 2391.910 ;
        RECT 1635.000 2385.770 1635.140 2391.910 ;
        RECT 1634.940 2385.450 1635.200 2385.770 ;
        RECT 2249.500 2385.450 2249.760 2385.770 ;
        RECT 1143.700 2373.880 1143.980 2377.880 ;
        RECT 2249.560 16.730 2249.700 2385.450 ;
        RECT 2249.560 16.590 2251.080 16.730 ;
        RECT 2250.940 2.400 2251.080 16.590 ;
        RECT 2250.730 -4.800 2251.290 2.400 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1772.910 1421.780 1773.230 1421.840 ;
        RECT 2052.590 1421.780 2052.910 1421.840 ;
        RECT 1772.910 1421.640 2052.910 1421.780 ;
        RECT 1772.910 1421.580 1773.230 1421.640 ;
        RECT 2052.590 1421.580 2052.910 1421.640 ;
        RECT 2052.590 19.280 2052.910 19.340 ;
        RECT 2268.330 19.280 2268.650 19.340 ;
        RECT 2052.590 19.140 2268.650 19.280 ;
        RECT 2052.590 19.080 2052.910 19.140 ;
        RECT 2268.330 19.080 2268.650 19.140 ;
      LAYER via ;
        RECT 1772.940 1421.580 1773.200 1421.840 ;
        RECT 2052.620 1421.580 2052.880 1421.840 ;
        RECT 2052.620 19.080 2052.880 19.340 ;
        RECT 2268.360 19.080 2268.620 19.340 ;
      LAYER met2 ;
        RECT 1772.930 1425.435 1773.210 1425.805 ;
        RECT 1773.000 1421.870 1773.140 1425.435 ;
        RECT 1772.940 1421.550 1773.200 1421.870 ;
        RECT 2052.620 1421.550 2052.880 1421.870 ;
        RECT 2052.680 19.370 2052.820 1421.550 ;
        RECT 2052.620 19.050 2052.880 19.370 ;
        RECT 2268.360 19.050 2268.620 19.370 ;
        RECT 2268.420 2.400 2268.560 19.050 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
      LAYER via2 ;
        RECT 1772.930 1425.480 1773.210 1425.760 ;
      LAYER met3 ;
        RECT 1755.835 1425.770 1759.835 1425.775 ;
        RECT 1772.905 1425.770 1773.235 1425.785 ;
        RECT 1755.835 1425.470 1773.235 1425.770 ;
        RECT 1755.835 1425.175 1759.835 1425.470 ;
        RECT 1772.905 1425.455 1773.235 1425.470 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 932.030 1317.400 932.350 1317.460 ;
        RECT 938.010 1317.400 938.330 1317.460 ;
        RECT 932.030 1317.260 938.330 1317.400 ;
        RECT 932.030 1317.200 932.350 1317.260 ;
        RECT 938.010 1317.200 938.330 1317.260 ;
        RECT 938.010 38.320 938.330 38.380 ;
        RECT 2286.270 38.320 2286.590 38.380 ;
        RECT 938.010 38.180 2286.590 38.320 ;
        RECT 938.010 38.120 938.330 38.180 ;
        RECT 2286.270 38.120 2286.590 38.180 ;
      LAYER via ;
        RECT 932.060 1317.200 932.320 1317.460 ;
        RECT 938.040 1317.200 938.300 1317.460 ;
        RECT 938.040 38.120 938.300 38.380 ;
        RECT 2286.300 38.120 2286.560 38.380 ;
      LAYER met2 ;
        RECT 932.100 1323.135 932.380 1327.135 ;
        RECT 932.120 1317.490 932.260 1323.135 ;
        RECT 932.060 1317.170 932.320 1317.490 ;
        RECT 938.040 1317.170 938.300 1317.490 ;
        RECT 938.100 38.410 938.240 1317.170 ;
        RECT 938.040 38.090 938.300 38.410 ;
        RECT 2286.300 38.090 2286.560 38.410 ;
        RECT 2286.360 2.400 2286.500 38.090 ;
        RECT 2286.150 -4.800 2286.710 2.400 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 696.970 1280.000 697.290 1280.060 ;
        RECT 2298.230 1280.000 2298.550 1280.060 ;
        RECT 696.970 1279.860 2298.550 1280.000 ;
        RECT 696.970 1279.800 697.290 1279.860 ;
        RECT 2298.230 1279.800 2298.550 1279.860 ;
        RECT 2298.230 24.720 2298.550 24.780 ;
        RECT 2304.210 24.720 2304.530 24.780 ;
        RECT 2298.230 24.580 2304.530 24.720 ;
        RECT 2298.230 24.520 2298.550 24.580 ;
        RECT 2304.210 24.520 2304.530 24.580 ;
      LAYER via ;
        RECT 697.000 1279.800 697.260 1280.060 ;
        RECT 2298.260 1279.800 2298.520 1280.060 ;
        RECT 2298.260 24.520 2298.520 24.780 ;
        RECT 2304.240 24.520 2304.500 24.780 ;
      LAYER met2 ;
        RECT 696.990 1806.235 697.270 1806.605 ;
        RECT 697.060 1280.090 697.200 1806.235 ;
        RECT 697.000 1279.770 697.260 1280.090 ;
        RECT 2298.260 1279.770 2298.520 1280.090 ;
        RECT 2298.320 24.810 2298.460 1279.770 ;
        RECT 2298.260 24.490 2298.520 24.810 ;
        RECT 2304.240 24.490 2304.500 24.810 ;
        RECT 2304.300 2.400 2304.440 24.490 ;
        RECT 2304.090 -4.800 2304.650 2.400 ;
      LAYER via2 ;
        RECT 696.990 1806.280 697.270 1806.560 ;
      LAYER met3 ;
        RECT 696.965 1806.570 697.295 1806.585 ;
        RECT 715.810 1806.570 719.810 1806.575 ;
        RECT 696.965 1806.270 719.810 1806.570 ;
        RECT 696.965 1806.255 697.295 1806.270 ;
        RECT 715.810 1805.975 719.810 1806.270 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1530.950 2388.400 1531.270 2388.460 ;
        RECT 1669.870 2388.400 1670.190 2388.460 ;
        RECT 1530.950 2388.260 1670.190 2388.400 ;
        RECT 1530.950 2388.200 1531.270 2388.260 ;
        RECT 1669.870 2388.200 1670.190 2388.260 ;
        RECT 1669.870 2385.340 1670.190 2385.400 ;
        RECT 2318.470 2385.340 2318.790 2385.400 ;
        RECT 1669.870 2385.200 2318.790 2385.340 ;
        RECT 1669.870 2385.140 1670.190 2385.200 ;
        RECT 2318.470 2385.140 2318.790 2385.200 ;
      LAYER via ;
        RECT 1530.980 2388.200 1531.240 2388.460 ;
        RECT 1669.900 2388.200 1670.160 2388.460 ;
        RECT 1669.900 2385.140 1670.160 2385.400 ;
        RECT 2318.500 2385.140 2318.760 2385.400 ;
      LAYER met2 ;
        RECT 1530.980 2388.170 1531.240 2388.490 ;
        RECT 1669.900 2388.170 1670.160 2388.490 ;
        RECT 1531.040 2377.880 1531.180 2388.170 ;
        RECT 1669.960 2385.430 1670.100 2388.170 ;
        RECT 1669.900 2385.110 1670.160 2385.430 ;
        RECT 2318.500 2385.110 2318.760 2385.430 ;
        RECT 1531.020 2373.880 1531.300 2377.880 ;
        RECT 2318.560 16.730 2318.700 2385.110 ;
        RECT 2318.560 16.590 2322.380 16.730 ;
        RECT 2322.240 2.400 2322.380 16.590 ;
        RECT 2322.030 -4.800 2322.590 2.400 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1612.445 17.425 1612.615 18.615 ;
      LAYER mcon ;
        RECT 1612.445 18.445 1612.615 18.615 ;
      LAYER met1 ;
        RECT 1612.385 18.600 1612.675 18.645 ;
        RECT 2339.630 18.600 2339.950 18.660 ;
        RECT 1612.385 18.460 2339.950 18.600 ;
        RECT 1612.385 18.415 1612.675 18.460 ;
        RECT 2339.630 18.400 2339.950 18.460 ;
        RECT 1593.510 17.580 1593.830 17.640 ;
        RECT 1612.385 17.580 1612.675 17.625 ;
        RECT 1593.510 17.440 1612.675 17.580 ;
        RECT 1593.510 17.380 1593.830 17.440 ;
        RECT 1612.385 17.395 1612.675 17.440 ;
      LAYER via ;
        RECT 2339.660 18.400 2339.920 18.660 ;
        RECT 1593.540 17.380 1593.800 17.640 ;
      LAYER met2 ;
        RECT 1591.740 1323.690 1592.020 1327.135 ;
        RECT 1591.740 1323.550 1593.740 1323.690 ;
        RECT 1591.740 1323.135 1592.020 1323.550 ;
        RECT 1593.600 17.670 1593.740 1323.550 ;
        RECT 2339.660 18.370 2339.920 18.690 ;
        RECT 1593.540 17.350 1593.800 17.670 ;
        RECT 2339.720 2.400 2339.860 18.370 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1398.470 2381.940 1398.790 2382.000 ;
        RECT 2352.970 2381.940 2353.290 2382.000 ;
        RECT 1398.470 2381.800 2353.290 2381.940 ;
        RECT 1398.470 2381.740 1398.790 2381.800 ;
        RECT 2352.970 2381.740 2353.290 2381.800 ;
        RECT 2352.970 62.120 2353.290 62.180 ;
        RECT 2357.570 62.120 2357.890 62.180 ;
        RECT 2352.970 61.980 2357.890 62.120 ;
        RECT 2352.970 61.920 2353.290 61.980 ;
        RECT 2357.570 61.920 2357.890 61.980 ;
      LAYER via ;
        RECT 1398.500 2381.740 1398.760 2382.000 ;
        RECT 2353.000 2381.740 2353.260 2382.000 ;
        RECT 2353.000 61.920 2353.260 62.180 ;
        RECT 2357.600 61.920 2357.860 62.180 ;
      LAYER met2 ;
        RECT 1398.500 2381.710 1398.760 2382.030 ;
        RECT 2353.000 2381.710 2353.260 2382.030 ;
        RECT 1398.560 2377.880 1398.700 2381.710 ;
        RECT 1398.540 2373.880 1398.820 2377.880 ;
        RECT 2353.060 62.210 2353.200 2381.710 ;
        RECT 2353.000 61.890 2353.260 62.210 ;
        RECT 2357.600 61.890 2357.860 62.210 ;
        RECT 2357.660 2.400 2357.800 61.890 ;
        RECT 2357.450 -4.800 2358.010 2.400 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1568.670 1311.280 1568.990 1311.340 ;
        RECT 1572.810 1311.280 1573.130 1311.340 ;
        RECT 1568.670 1311.140 1573.130 1311.280 ;
        RECT 1568.670 1311.080 1568.990 1311.140 ;
        RECT 1572.810 1311.080 1573.130 1311.140 ;
        RECT 1572.810 17.920 1573.130 17.980 ;
        RECT 2375.510 17.920 2375.830 17.980 ;
        RECT 1572.810 17.780 2375.830 17.920 ;
        RECT 1572.810 17.720 1573.130 17.780 ;
        RECT 2375.510 17.720 2375.830 17.780 ;
      LAYER via ;
        RECT 1568.700 1311.080 1568.960 1311.340 ;
        RECT 1572.840 1311.080 1573.100 1311.340 ;
        RECT 1572.840 17.720 1573.100 17.980 ;
        RECT 2375.540 17.720 2375.800 17.980 ;
      LAYER met2 ;
        RECT 1568.740 1323.135 1569.020 1327.135 ;
        RECT 1568.760 1311.370 1568.900 1323.135 ;
        RECT 1568.700 1311.050 1568.960 1311.370 ;
        RECT 1572.840 1311.050 1573.100 1311.370 ;
        RECT 1572.900 18.010 1573.040 1311.050 ;
        RECT 1572.840 17.690 1573.100 18.010 ;
        RECT 2375.540 17.690 2375.800 18.010 ;
        RECT 2375.600 2.400 2375.740 17.690 ;
        RECT 2375.390 -4.800 2375.950 2.400 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1744.465 58.225 1744.635 62.475 ;
      LAYER mcon ;
        RECT 1744.465 62.305 1744.635 62.475 ;
      LAYER met1 ;
        RECT 1744.390 62.460 1744.710 62.520 ;
        RECT 1744.195 62.320 1744.710 62.460 ;
        RECT 1744.390 62.260 1744.710 62.320 ;
        RECT 1744.390 58.380 1744.710 58.440 ;
        RECT 1744.195 58.240 1744.710 58.380 ;
        RECT 1744.390 58.180 1744.710 58.240 ;
        RECT 1744.390 18.940 1744.710 19.000 ;
        RECT 2393.450 18.940 2393.770 19.000 ;
        RECT 1744.390 18.800 2393.770 18.940 ;
        RECT 1744.390 18.740 1744.710 18.800 ;
        RECT 2393.450 18.740 2393.770 18.800 ;
      LAYER via ;
        RECT 1744.420 62.260 1744.680 62.520 ;
        RECT 1744.420 58.180 1744.680 58.440 ;
        RECT 1744.420 18.740 1744.680 19.000 ;
        RECT 2393.480 18.740 2393.740 19.000 ;
      LAYER met2 ;
        RECT 1741.700 1323.690 1741.980 1327.135 ;
        RECT 1741.700 1323.550 1744.620 1323.690 ;
        RECT 1741.700 1323.135 1741.980 1323.550 ;
        RECT 1744.480 62.550 1744.620 1323.550 ;
        RECT 1744.420 62.230 1744.680 62.550 ;
        RECT 1744.420 58.150 1744.680 58.470 ;
        RECT 1744.480 19.030 1744.620 58.150 ;
        RECT 1744.420 18.710 1744.680 19.030 ;
        RECT 2393.480 18.710 2393.740 19.030 ;
        RECT 2393.540 2.400 2393.680 18.710 ;
        RECT 2393.330 -4.800 2393.890 2.400 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 718.205 1797.325 718.375 1813.135 ;
        RECT 717.285 1728.305 717.455 1734.935 ;
        RECT 717.745 1656.225 717.915 1696.175 ;
      LAYER mcon ;
        RECT 718.205 1812.965 718.375 1813.135 ;
        RECT 717.285 1734.765 717.455 1734.935 ;
        RECT 717.745 1696.005 717.915 1696.175 ;
      LAYER met1 ;
        RECT 718.145 1813.120 718.435 1813.165 ;
        RECT 718.590 1813.120 718.910 1813.180 ;
        RECT 718.145 1812.980 718.910 1813.120 ;
        RECT 718.145 1812.935 718.435 1812.980 ;
        RECT 718.590 1812.920 718.910 1812.980 ;
        RECT 717.210 1797.480 717.530 1797.540 ;
        RECT 718.145 1797.480 718.435 1797.525 ;
        RECT 717.210 1797.340 718.435 1797.480 ;
        RECT 717.210 1797.280 717.530 1797.340 ;
        RECT 718.145 1797.295 718.435 1797.340 ;
        RECT 717.210 1734.920 717.530 1734.980 ;
        RECT 717.015 1734.780 717.530 1734.920 ;
        RECT 717.210 1734.720 717.530 1734.780 ;
        RECT 717.210 1728.460 717.530 1728.520 ;
        RECT 717.015 1728.320 717.530 1728.460 ;
        RECT 717.210 1728.260 717.530 1728.320 ;
        RECT 717.210 1696.160 717.530 1696.220 ;
        RECT 717.685 1696.160 717.975 1696.205 ;
        RECT 717.210 1696.020 717.975 1696.160 ;
        RECT 717.210 1695.960 717.530 1696.020 ;
        RECT 717.685 1695.975 717.975 1696.020 ;
        RECT 713.990 1656.380 714.310 1656.440 ;
        RECT 717.685 1656.380 717.975 1656.425 ;
        RECT 713.990 1656.240 717.975 1656.380 ;
        RECT 713.990 1656.180 714.310 1656.240 ;
        RECT 717.685 1656.195 717.975 1656.240 ;
        RECT 2408.170 62.120 2408.490 62.180 ;
        RECT 2411.390 62.120 2411.710 62.180 ;
        RECT 2408.170 61.980 2411.710 62.120 ;
        RECT 2408.170 61.920 2408.490 61.980 ;
        RECT 2411.390 61.920 2411.710 61.980 ;
      LAYER via ;
        RECT 718.620 1812.920 718.880 1813.180 ;
        RECT 717.240 1797.280 717.500 1797.540 ;
        RECT 717.240 1734.720 717.500 1734.980 ;
        RECT 717.240 1728.260 717.500 1728.520 ;
        RECT 717.240 1695.960 717.500 1696.220 ;
        RECT 714.020 1656.180 714.280 1656.440 ;
        RECT 2408.200 61.920 2408.460 62.180 ;
        RECT 2411.420 61.920 2411.680 62.180 ;
      LAYER met2 ;
        RECT 713.090 2011.595 713.370 2011.965 ;
        RECT 713.160 1963.005 713.300 2011.595 ;
        RECT 713.090 1962.635 713.370 1963.005 ;
        RECT 718.610 1821.195 718.890 1821.565 ;
        RECT 718.680 1813.210 718.820 1821.195 ;
        RECT 718.620 1812.890 718.880 1813.210 ;
        RECT 717.240 1797.250 717.500 1797.570 ;
        RECT 717.300 1735.010 717.440 1797.250 ;
        RECT 717.240 1734.690 717.500 1735.010 ;
        RECT 717.240 1728.230 717.500 1728.550 ;
        RECT 717.300 1696.250 717.440 1728.230 ;
        RECT 717.240 1695.930 717.500 1696.250 ;
        RECT 714.020 1656.150 714.280 1656.470 ;
        RECT 714.080 1650.205 714.220 1656.150 ;
        RECT 714.010 1649.835 714.290 1650.205 ;
        RECT 722.290 1014.035 722.570 1014.405 ;
        RECT 722.360 967.485 722.500 1014.035 ;
        RECT 722.290 967.115 722.570 967.485 ;
        RECT 722.750 820.235 723.030 820.605 ;
        RECT 722.820 773.685 722.960 820.235 ;
        RECT 722.750 773.315 723.030 773.685 ;
        RECT 722.750 723.675 723.030 724.045 ;
        RECT 722.820 677.125 722.960 723.675 ;
        RECT 722.750 676.755 723.030 677.125 ;
        RECT 722.290 433.995 722.570 434.365 ;
        RECT 722.360 386.765 722.500 433.995 ;
        RECT 722.290 386.395 722.570 386.765 ;
        RECT 722.750 143.635 723.030 144.005 ;
        RECT 722.820 97.765 722.960 143.635 ;
        RECT 722.750 97.395 723.030 97.765 ;
        RECT 2408.190 79.715 2408.470 80.085 ;
        RECT 2408.260 62.210 2408.400 79.715 ;
        RECT 2408.200 61.890 2408.460 62.210 ;
        RECT 2411.420 61.890 2411.680 62.210 ;
        RECT 2411.480 2.400 2411.620 61.890 ;
        RECT 2411.270 -4.800 2411.830 2.400 ;
      LAYER via2 ;
        RECT 713.090 2011.640 713.370 2011.920 ;
        RECT 713.090 1962.680 713.370 1962.960 ;
        RECT 718.610 1821.240 718.890 1821.520 ;
        RECT 714.010 1649.880 714.290 1650.160 ;
        RECT 722.290 1014.080 722.570 1014.360 ;
        RECT 722.290 967.160 722.570 967.440 ;
        RECT 722.750 820.280 723.030 820.560 ;
        RECT 722.750 773.360 723.030 773.640 ;
        RECT 722.750 723.720 723.030 724.000 ;
        RECT 722.750 676.800 723.030 677.080 ;
        RECT 722.290 434.040 722.570 434.320 ;
        RECT 722.290 386.440 722.570 386.720 ;
        RECT 722.750 143.680 723.030 143.960 ;
        RECT 722.750 97.440 723.030 97.720 ;
        RECT 2408.190 79.760 2408.470 80.040 ;
      LAYER met3 ;
        RECT 713.065 2011.930 713.395 2011.945 ;
        RECT 715.810 2011.930 719.810 2011.935 ;
        RECT 713.065 2011.630 719.810 2011.930 ;
        RECT 713.065 2011.615 713.395 2011.630 ;
        RECT 715.810 2011.335 719.810 2011.630 ;
        RECT 713.065 1962.970 713.395 1962.985 ;
        RECT 714.190 1962.970 714.570 1962.980 ;
        RECT 713.065 1962.670 714.570 1962.970 ;
        RECT 713.065 1962.655 713.395 1962.670 ;
        RECT 714.190 1962.660 714.570 1962.670 ;
        RECT 714.190 1905.850 714.570 1905.860 ;
        RECT 714.190 1905.550 719.130 1905.850 ;
        RECT 714.190 1905.540 714.570 1905.550 ;
        RECT 718.830 1904.500 719.130 1905.550 ;
        RECT 718.790 1904.180 719.170 1904.500 ;
        RECT 714.190 1862.330 714.570 1862.340 ;
        RECT 718.790 1862.330 719.170 1862.340 ;
        RECT 714.190 1862.030 719.170 1862.330 ;
        RECT 714.190 1862.020 714.570 1862.030 ;
        RECT 718.790 1862.020 719.170 1862.030 ;
        RECT 714.190 1849.410 714.570 1849.420 ;
        RECT 718.790 1849.410 719.170 1849.420 ;
        RECT 714.190 1849.110 719.170 1849.410 ;
        RECT 714.190 1849.100 714.570 1849.110 ;
        RECT 718.790 1849.100 719.170 1849.110 ;
        RECT 718.585 1821.540 718.915 1821.545 ;
        RECT 718.585 1821.530 719.170 1821.540 ;
        RECT 718.360 1821.230 719.170 1821.530 ;
        RECT 718.585 1821.220 719.170 1821.230 ;
        RECT 718.585 1821.215 718.915 1821.220 ;
        RECT 713.985 1650.170 714.315 1650.185 ;
        RECT 718.790 1650.170 719.170 1650.180 ;
        RECT 713.985 1649.870 719.170 1650.170 ;
        RECT 713.985 1649.855 714.315 1649.870 ;
        RECT 718.790 1649.860 719.170 1649.870 ;
        RECT 718.790 1641.700 719.170 1642.020 ;
        RECT 714.190 1640.650 714.570 1640.660 ;
        RECT 718.830 1640.650 719.130 1641.700 ;
        RECT 714.190 1640.350 719.130 1640.650 ;
        RECT 714.190 1640.340 714.570 1640.350 ;
        RECT 714.190 1622.970 714.570 1622.980 ;
        RECT 716.950 1622.970 717.330 1622.980 ;
        RECT 714.190 1622.670 717.330 1622.970 ;
        RECT 714.190 1622.660 714.570 1622.670 ;
        RECT 716.950 1622.660 717.330 1622.670 ;
        RECT 691.190 1546.810 691.570 1546.820 ;
        RECT 716.950 1546.810 717.330 1546.820 ;
        RECT 691.190 1546.510 717.330 1546.810 ;
        RECT 691.190 1546.500 691.570 1546.510 ;
        RECT 716.950 1546.500 717.330 1546.510 ;
        RECT 717.870 1373.100 718.250 1373.420 ;
        RECT 717.910 1372.050 718.210 1373.100 ;
        RECT 718.790 1372.050 719.170 1372.060 ;
        RECT 717.910 1371.750 719.170 1372.050 ;
        RECT 718.790 1371.740 719.170 1371.750 ;
        RECT 722.265 1014.380 722.595 1014.385 ;
        RECT 722.265 1014.370 722.850 1014.380 ;
        RECT 722.040 1014.070 722.850 1014.370 ;
        RECT 722.265 1014.060 722.850 1014.070 ;
        RECT 722.265 1014.055 722.595 1014.060 ;
        RECT 722.265 967.450 722.595 967.465 ;
        RECT 722.265 967.135 722.810 967.450 ;
        RECT 722.510 966.780 722.810 967.135 ;
        RECT 722.470 966.460 722.850 966.780 ;
        RECT 722.725 820.580 723.055 820.585 ;
        RECT 722.470 820.570 723.055 820.580 ;
        RECT 722.470 820.270 723.280 820.570 ;
        RECT 722.470 820.260 723.055 820.270 ;
        RECT 722.725 820.255 723.055 820.260 ;
        RECT 722.725 773.650 723.055 773.665 ;
        RECT 722.510 773.335 723.055 773.650 ;
        RECT 722.510 772.980 722.810 773.335 ;
        RECT 722.470 772.660 722.850 772.980 ;
        RECT 722.725 724.020 723.055 724.025 ;
        RECT 722.470 724.010 723.055 724.020 ;
        RECT 722.470 723.710 723.280 724.010 ;
        RECT 722.470 723.700 723.055 723.710 ;
        RECT 722.725 723.695 723.055 723.700 ;
        RECT 722.725 677.090 723.055 677.105 ;
        RECT 722.510 676.775 723.055 677.090 ;
        RECT 722.510 676.420 722.810 676.775 ;
        RECT 722.470 676.100 722.850 676.420 ;
        RECT 722.470 485.020 722.850 485.340 ;
        RECT 722.510 483.300 722.810 485.020 ;
        RECT 722.470 482.980 722.850 483.300 ;
        RECT 722.265 434.340 722.595 434.345 ;
        RECT 722.265 434.330 722.850 434.340 ;
        RECT 722.040 434.030 722.850 434.330 ;
        RECT 722.265 434.020 722.850 434.030 ;
        RECT 722.265 434.015 722.595 434.020 ;
        RECT 722.265 386.740 722.595 386.745 ;
        RECT 722.265 386.730 722.850 386.740 ;
        RECT 722.040 386.430 722.850 386.730 ;
        RECT 722.265 386.420 722.850 386.430 ;
        RECT 722.265 386.415 722.595 386.420 ;
        RECT 722.470 193.980 722.850 194.300 ;
        RECT 722.510 193.620 722.810 193.980 ;
        RECT 722.470 193.300 722.850 193.620 ;
        RECT 722.725 143.980 723.055 143.985 ;
        RECT 722.470 143.970 723.055 143.980 ;
        RECT 722.470 143.670 723.280 143.970 ;
        RECT 722.470 143.660 723.055 143.670 ;
        RECT 722.725 143.655 723.055 143.660 ;
        RECT 722.725 97.740 723.055 97.745 ;
        RECT 722.470 97.730 723.055 97.740 ;
        RECT 722.270 97.430 723.055 97.730 ;
        RECT 722.470 97.420 723.055 97.430 ;
        RECT 722.725 97.415 723.055 97.420 ;
        RECT 722.470 80.050 722.850 80.060 ;
        RECT 2408.165 80.050 2408.495 80.065 ;
        RECT 722.470 79.750 2408.495 80.050 ;
        RECT 722.470 79.740 722.850 79.750 ;
        RECT 2408.165 79.735 2408.495 79.750 ;
      LAYER via3 ;
        RECT 714.220 1962.660 714.540 1962.980 ;
        RECT 714.220 1905.540 714.540 1905.860 ;
        RECT 718.820 1904.180 719.140 1904.500 ;
        RECT 714.220 1862.020 714.540 1862.340 ;
        RECT 718.820 1862.020 719.140 1862.340 ;
        RECT 714.220 1849.100 714.540 1849.420 ;
        RECT 718.820 1849.100 719.140 1849.420 ;
        RECT 718.820 1821.220 719.140 1821.540 ;
        RECT 718.820 1649.860 719.140 1650.180 ;
        RECT 718.820 1641.700 719.140 1642.020 ;
        RECT 714.220 1640.340 714.540 1640.660 ;
        RECT 714.220 1622.660 714.540 1622.980 ;
        RECT 716.980 1622.660 717.300 1622.980 ;
        RECT 691.220 1546.500 691.540 1546.820 ;
        RECT 716.980 1546.500 717.300 1546.820 ;
        RECT 717.900 1373.100 718.220 1373.420 ;
        RECT 718.820 1371.740 719.140 1372.060 ;
        RECT 722.500 1014.060 722.820 1014.380 ;
        RECT 722.500 966.460 722.820 966.780 ;
        RECT 722.500 820.260 722.820 820.580 ;
        RECT 722.500 772.660 722.820 772.980 ;
        RECT 722.500 723.700 722.820 724.020 ;
        RECT 722.500 676.100 722.820 676.420 ;
        RECT 722.500 485.020 722.820 485.340 ;
        RECT 722.500 482.980 722.820 483.300 ;
        RECT 722.500 434.020 722.820 434.340 ;
        RECT 722.500 386.420 722.820 386.740 ;
        RECT 722.500 193.980 722.820 194.300 ;
        RECT 722.500 193.300 722.820 193.620 ;
        RECT 722.500 143.660 722.820 143.980 ;
        RECT 722.500 97.420 722.820 97.740 ;
        RECT 722.500 79.740 722.820 80.060 ;
      LAYER met4 ;
        RECT 714.215 1962.655 714.545 1962.985 ;
        RECT 714.230 1905.865 714.530 1962.655 ;
        RECT 714.215 1905.535 714.545 1905.865 ;
        RECT 718.815 1904.175 719.145 1904.505 ;
        RECT 718.830 1862.345 719.130 1904.175 ;
        RECT 714.215 1862.015 714.545 1862.345 ;
        RECT 718.815 1862.015 719.145 1862.345 ;
        RECT 714.230 1849.425 714.530 1862.015 ;
        RECT 714.215 1849.095 714.545 1849.425 ;
        RECT 718.815 1849.095 719.145 1849.425 ;
        RECT 718.830 1821.545 719.130 1849.095 ;
        RECT 718.815 1821.215 719.145 1821.545 ;
        RECT 718.815 1649.855 719.145 1650.185 ;
        RECT 718.830 1642.025 719.130 1649.855 ;
        RECT 718.815 1641.695 719.145 1642.025 ;
        RECT 714.215 1640.335 714.545 1640.665 ;
        RECT 714.230 1622.985 714.530 1640.335 ;
        RECT 714.215 1622.655 714.545 1622.985 ;
        RECT 716.975 1622.655 717.305 1622.985 ;
        RECT 716.990 1546.825 717.290 1622.655 ;
        RECT 691.215 1546.495 691.545 1546.825 ;
        RECT 716.975 1546.495 717.305 1546.825 ;
        RECT 691.230 1505.090 691.530 1546.495 ;
        RECT 690.790 1503.910 691.970 1505.090 ;
        RECT 719.310 1483.510 720.490 1484.690 ;
        RECT 719.750 1470.650 720.050 1483.510 ;
        RECT 719.750 1470.350 722.810 1470.650 ;
        RECT 722.510 1468.610 722.810 1470.350 ;
        RECT 721.590 1468.310 722.810 1468.610 ;
        RECT 721.590 1467.250 721.890 1468.310 ;
        RECT 721.590 1466.950 722.810 1467.250 ;
        RECT 722.510 1429.850 722.810 1466.950 ;
        RECT 717.910 1429.550 722.810 1429.850 ;
        RECT 717.910 1373.425 718.210 1429.550 ;
        RECT 717.895 1373.095 718.225 1373.425 ;
        RECT 718.815 1371.735 719.145 1372.065 ;
        RECT 718.830 1351.650 719.130 1371.735 ;
        RECT 718.830 1351.350 722.810 1351.650 ;
        RECT 722.510 1014.385 722.810 1351.350 ;
        RECT 722.495 1014.055 722.825 1014.385 ;
        RECT 722.495 966.455 722.825 966.785 ;
        RECT 722.510 820.585 722.810 966.455 ;
        RECT 722.495 820.255 722.825 820.585 ;
        RECT 722.495 772.655 722.825 772.985 ;
        RECT 722.510 724.025 722.810 772.655 ;
        RECT 722.495 723.695 722.825 724.025 ;
        RECT 722.495 676.095 722.825 676.425 ;
        RECT 722.510 485.345 722.810 676.095 ;
        RECT 722.495 485.015 722.825 485.345 ;
        RECT 722.495 482.975 722.825 483.305 ;
        RECT 722.510 434.345 722.810 482.975 ;
        RECT 722.495 434.015 722.825 434.345 ;
        RECT 722.495 386.415 722.825 386.745 ;
        RECT 722.510 194.305 722.810 386.415 ;
        RECT 722.495 193.975 722.825 194.305 ;
        RECT 722.495 193.295 722.825 193.625 ;
        RECT 722.510 143.985 722.810 193.295 ;
        RECT 722.495 143.655 722.825 143.985 ;
        RECT 722.495 97.415 722.825 97.745 ;
        RECT 722.510 80.065 722.810 97.415 ;
        RECT 722.495 79.735 722.825 80.065 ;
      LAYER met5 ;
        RECT 690.580 1503.700 705.060 1505.300 ;
        RECT 703.460 1498.500 705.060 1503.700 ;
        RECT 703.460 1496.900 706.900 1498.500 ;
        RECT 705.300 1484.900 706.900 1496.900 ;
        RECT 705.300 1483.300 720.700 1484.900 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 806.910 1312.980 807.230 1313.040 ;
        RECT 1406.750 1312.980 1407.070 1313.040 ;
        RECT 806.910 1312.840 1407.070 1312.980 ;
        RECT 806.910 1312.780 807.230 1312.840 ;
        RECT 1406.750 1312.780 1407.070 1312.840 ;
        RECT 805.530 62.120 805.850 62.180 ;
        RECT 806.910 62.120 807.230 62.180 ;
        RECT 805.530 61.980 807.230 62.120 ;
        RECT 805.530 61.920 805.850 61.980 ;
        RECT 806.910 61.920 807.230 61.980 ;
      LAYER via ;
        RECT 806.940 1312.780 807.200 1313.040 ;
        RECT 1406.780 1312.780 1407.040 1313.040 ;
        RECT 805.560 61.920 805.820 62.180 ;
        RECT 806.940 61.920 807.200 62.180 ;
      LAYER met2 ;
        RECT 1406.820 1323.135 1407.100 1327.135 ;
        RECT 1406.840 1313.070 1406.980 1323.135 ;
        RECT 806.940 1312.750 807.200 1313.070 ;
        RECT 1406.780 1312.750 1407.040 1313.070 ;
        RECT 807.000 62.210 807.140 1312.750 ;
        RECT 805.560 61.890 805.820 62.210 ;
        RECT 806.940 61.890 807.200 62.210 ;
        RECT 805.620 2.400 805.760 61.890 ;
        RECT 805.410 -4.800 805.970 2.400 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2.830 24.040 3.150 24.100 ;
        RECT 1090.270 24.040 1090.590 24.100 ;
        RECT 2.830 23.900 1090.590 24.040 ;
        RECT 2.830 23.840 3.150 23.900 ;
        RECT 1090.270 23.840 1090.590 23.900 ;
      LAYER via ;
        RECT 2.860 23.840 3.120 24.100 ;
        RECT 1090.300 23.840 1090.560 24.100 ;
      LAYER met2 ;
        RECT 1094.020 1323.690 1094.300 1327.135 ;
        RECT 1090.360 1323.550 1094.300 1323.690 ;
        RECT 1090.360 24.130 1090.500 1323.550 ;
        RECT 1094.020 1323.135 1094.300 1323.550 ;
        RECT 2.860 23.810 3.120 24.130 ;
        RECT 1090.300 23.810 1090.560 24.130 ;
        RECT 2.920 2.400 3.060 23.810 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 726.870 2380.240 727.190 2380.300 ;
        RECT 712.700 2380.100 727.190 2380.240 ;
        RECT 13.410 2379.900 13.730 2379.960 ;
        RECT 712.700 2379.900 712.840 2380.100 ;
        RECT 726.870 2380.040 727.190 2380.100 ;
        RECT 13.410 2379.760 712.840 2379.900 ;
        RECT 13.410 2379.700 13.730 2379.760 ;
        RECT 8.350 17.580 8.670 17.640 ;
        RECT 13.410 17.580 13.730 17.640 ;
        RECT 8.350 17.440 13.730 17.580 ;
        RECT 8.350 17.380 8.670 17.440 ;
        RECT 13.410 17.380 13.730 17.440 ;
      LAYER via ;
        RECT 13.440 2379.700 13.700 2379.960 ;
        RECT 726.900 2380.040 727.160 2380.300 ;
        RECT 8.380 17.380 8.640 17.640 ;
        RECT 13.440 17.380 13.700 17.640 ;
      LAYER met2 ;
        RECT 726.900 2380.010 727.160 2380.330 ;
        RECT 13.440 2379.670 13.700 2379.990 ;
        RECT 13.500 17.670 13.640 2379.670 ;
        RECT 726.960 2377.880 727.100 2380.010 ;
        RECT 726.940 2373.880 727.220 2377.880 ;
        RECT 8.380 17.350 8.640 17.670 ;
        RECT 13.440 17.350 13.700 17.670 ;
        RECT 8.440 2.400 8.580 17.350 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 14.330 17.920 14.650 17.980 ;
        RECT 20.310 17.920 20.630 17.980 ;
        RECT 14.330 17.780 20.630 17.920 ;
        RECT 14.330 17.720 14.650 17.780 ;
        RECT 20.310 17.720 20.630 17.780 ;
      LAYER via ;
        RECT 14.360 17.720 14.620 17.980 ;
        RECT 20.340 17.720 20.600 17.980 ;
      LAYER met2 ;
        RECT 20.330 2378.795 20.610 2379.165 ;
        RECT 1147.330 2378.795 1147.610 2379.165 ;
        RECT 20.400 18.010 20.540 2378.795 ;
        RECT 1147.400 2377.690 1147.540 2378.795 ;
        RECT 1149.220 2377.690 1149.500 2377.880 ;
        RECT 1147.400 2377.550 1149.500 2377.690 ;
        RECT 1149.220 2373.880 1149.500 2377.550 ;
        RECT 14.360 17.690 14.620 18.010 ;
        RECT 20.340 17.690 20.600 18.010 ;
        RECT 14.420 2.400 14.560 17.690 ;
        RECT 14.210 -4.800 14.770 2.400 ;
      LAYER via2 ;
        RECT 20.330 2378.840 20.610 2379.120 ;
        RECT 1147.330 2378.840 1147.610 2379.120 ;
      LAYER met3 ;
        RECT 20.305 2379.130 20.635 2379.145 ;
        RECT 1147.305 2379.130 1147.635 2379.145 ;
        RECT 20.305 2378.830 1147.635 2379.130 ;
        RECT 20.305 2378.815 20.635 2378.830 ;
        RECT 1147.305 2378.815 1147.635 2378.830 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 40.550 1842.700 40.870 1842.760 ;
        RECT 692.370 1842.700 692.690 1842.760 ;
        RECT 40.550 1842.560 692.690 1842.700 ;
        RECT 40.550 1842.500 40.870 1842.560 ;
        RECT 692.370 1842.500 692.690 1842.560 ;
        RECT 38.250 17.920 38.570 17.980 ;
        RECT 40.550 17.920 40.870 17.980 ;
        RECT 38.250 17.780 40.870 17.920 ;
        RECT 38.250 17.720 38.570 17.780 ;
        RECT 40.550 17.720 40.870 17.780 ;
      LAYER via ;
        RECT 40.580 1842.500 40.840 1842.760 ;
        RECT 692.400 1842.500 692.660 1842.760 ;
        RECT 38.280 17.720 38.540 17.980 ;
        RECT 40.580 17.720 40.840 17.980 ;
      LAYER met2 ;
        RECT 692.390 1848.395 692.670 1848.765 ;
        RECT 692.460 1842.790 692.600 1848.395 ;
        RECT 40.580 1842.470 40.840 1842.790 ;
        RECT 692.400 1842.470 692.660 1842.790 ;
        RECT 40.640 18.010 40.780 1842.470 ;
        RECT 38.280 17.690 38.540 18.010 ;
        RECT 40.580 17.690 40.840 18.010 ;
        RECT 38.340 2.400 38.480 17.690 ;
        RECT 38.130 -4.800 38.690 2.400 ;
      LAYER via2 ;
        RECT 692.390 1848.440 692.670 1848.720 ;
      LAYER met3 ;
        RECT 692.365 1848.730 692.695 1848.745 ;
        RECT 715.810 1848.730 719.810 1848.735 ;
        RECT 692.365 1848.430 719.810 1848.730 ;
        RECT 692.365 1848.415 692.695 1848.430 ;
        RECT 715.810 1848.135 719.810 1848.430 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 240.670 23.955 240.950 24.325 ;
        RECT 240.740 2.400 240.880 23.955 ;
        RECT 240.530 -4.800 241.090 2.400 ;
      LAYER via2 ;
        RECT 240.670 24.000 240.950 24.280 ;
      LAYER met3 ;
        RECT 1755.835 2237.095 1759.835 2237.695 ;
        RECT 1759.350 2236.340 1759.650 2237.095 ;
        RECT 1759.310 2236.020 1759.690 2236.340 ;
        RECT 240.645 24.290 240.975 24.305 ;
        RECT 1759.310 24.290 1759.690 24.300 ;
        RECT 240.645 23.990 1759.690 24.290 ;
        RECT 240.645 23.975 240.975 23.990 ;
        RECT 1759.310 23.980 1759.690 23.990 ;
      LAYER via3 ;
        RECT 1759.340 2236.020 1759.660 2236.340 ;
        RECT 1759.340 23.980 1759.660 24.300 ;
      LAYER met4 ;
        RECT 1759.335 2236.015 1759.665 2236.345 ;
        RECT 1759.350 24.305 1759.650 2236.015 ;
        RECT 1759.335 23.975 1759.665 24.305 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 265.490 1315.360 265.810 1315.420 ;
        RECT 1302.790 1315.360 1303.110 1315.420 ;
        RECT 265.490 1315.220 1303.110 1315.360 ;
        RECT 265.490 1315.160 265.810 1315.220 ;
        RECT 1302.790 1315.160 1303.110 1315.220 ;
        RECT 258.130 17.240 258.450 17.300 ;
        RECT 265.490 17.240 265.810 17.300 ;
        RECT 258.130 17.100 265.810 17.240 ;
        RECT 258.130 17.040 258.450 17.100 ;
        RECT 265.490 17.040 265.810 17.100 ;
      LAYER via ;
        RECT 265.520 1315.160 265.780 1315.420 ;
        RECT 1302.820 1315.160 1303.080 1315.420 ;
        RECT 258.160 17.040 258.420 17.300 ;
        RECT 265.520 17.040 265.780 17.300 ;
      LAYER met2 ;
        RECT 1302.860 1323.135 1303.140 1327.135 ;
        RECT 1302.880 1315.450 1303.020 1323.135 ;
        RECT 265.520 1315.130 265.780 1315.450 ;
        RECT 1302.820 1315.130 1303.080 1315.450 ;
        RECT 265.580 17.330 265.720 1315.130 ;
        RECT 258.160 17.010 258.420 17.330 ;
        RECT 265.520 17.010 265.780 17.330 ;
        RECT 258.220 2.400 258.360 17.010 ;
        RECT 258.010 -4.800 258.570 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 949.510 1311.960 949.830 1312.020 ;
        RECT 926.600 1311.820 949.830 1311.960 ;
        RECT 282.510 1311.280 282.830 1311.340 ;
        RECT 926.600 1311.280 926.740 1311.820 ;
        RECT 949.510 1311.760 949.830 1311.820 ;
        RECT 282.510 1311.140 926.740 1311.280 ;
        RECT 282.510 1311.080 282.830 1311.140 ;
        RECT 276.070 16.900 276.390 16.960 ;
        RECT 282.510 16.900 282.830 16.960 ;
        RECT 276.070 16.760 282.830 16.900 ;
        RECT 276.070 16.700 276.390 16.760 ;
        RECT 282.510 16.700 282.830 16.760 ;
      LAYER via ;
        RECT 282.540 1311.080 282.800 1311.340 ;
        RECT 949.540 1311.760 949.800 1312.020 ;
        RECT 276.100 16.700 276.360 16.960 ;
        RECT 282.540 16.700 282.800 16.960 ;
      LAYER met2 ;
        RECT 949.580 1323.135 949.860 1327.135 ;
        RECT 949.600 1312.050 949.740 1323.135 ;
        RECT 949.540 1311.730 949.800 1312.050 ;
        RECT 282.540 1311.050 282.800 1311.370 ;
        RECT 282.600 16.990 282.740 1311.050 ;
        RECT 276.100 16.670 276.360 16.990 ;
        RECT 282.540 16.670 282.800 16.990 ;
        RECT 276.160 2.400 276.300 16.670 ;
        RECT 275.950 -4.800 276.510 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 334.490 1316.040 334.810 1316.100 ;
        RECT 1343.270 1316.040 1343.590 1316.100 ;
        RECT 334.490 1315.900 1343.590 1316.040 ;
        RECT 334.490 1315.840 334.810 1315.900 ;
        RECT 1343.270 1315.840 1343.590 1315.900 ;
        RECT 294.010 16.220 294.330 16.280 ;
        RECT 334.490 16.220 334.810 16.280 ;
        RECT 294.010 16.080 334.810 16.220 ;
        RECT 294.010 16.020 294.330 16.080 ;
        RECT 334.490 16.020 334.810 16.080 ;
      LAYER via ;
        RECT 334.520 1315.840 334.780 1316.100 ;
        RECT 1343.300 1315.840 1343.560 1316.100 ;
        RECT 294.040 16.020 294.300 16.280 ;
        RECT 334.520 16.020 334.780 16.280 ;
      LAYER met2 ;
        RECT 1343.340 1323.135 1343.620 1327.135 ;
        RECT 1343.360 1316.130 1343.500 1323.135 ;
        RECT 334.520 1315.810 334.780 1316.130 ;
        RECT 1343.300 1315.810 1343.560 1316.130 ;
        RECT 334.580 16.310 334.720 1315.810 ;
        RECT 294.040 15.990 294.300 16.310 ;
        RECT 334.520 15.990 334.780 16.310 ;
        RECT 294.100 2.400 294.240 15.990 ;
        RECT 293.890 -4.800 294.450 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 317.010 2379.220 317.330 2379.280 ;
        RECT 842.790 2379.220 843.110 2379.280 ;
        RECT 317.010 2379.080 843.110 2379.220 ;
        RECT 317.010 2379.020 317.330 2379.080 ;
        RECT 842.790 2379.020 843.110 2379.080 ;
        RECT 311.950 16.900 312.270 16.960 ;
        RECT 317.010 16.900 317.330 16.960 ;
        RECT 311.950 16.760 317.330 16.900 ;
        RECT 311.950 16.700 312.270 16.760 ;
        RECT 317.010 16.700 317.330 16.760 ;
      LAYER via ;
        RECT 317.040 2379.020 317.300 2379.280 ;
        RECT 842.820 2379.020 843.080 2379.280 ;
        RECT 311.980 16.700 312.240 16.960 ;
        RECT 317.040 16.700 317.300 16.960 ;
      LAYER met2 ;
        RECT 317.040 2378.990 317.300 2379.310 ;
        RECT 842.820 2378.990 843.080 2379.310 ;
        RECT 317.100 16.990 317.240 2378.990 ;
        RECT 842.880 2377.880 843.020 2378.990 ;
        RECT 842.860 2373.880 843.140 2377.880 ;
        RECT 311.980 16.670 312.240 16.990 ;
        RECT 317.040 16.670 317.300 16.990 ;
        RECT 312.040 2.400 312.180 16.670 ;
        RECT 311.830 -4.800 312.390 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 713.145 2377.705 713.315 2379.915 ;
      LAYER mcon ;
        RECT 713.145 2379.745 713.315 2379.915 ;
      LAYER met1 ;
        RECT 713.085 2379.900 713.375 2379.945 ;
        RECT 756.310 2379.900 756.630 2379.960 ;
        RECT 713.085 2379.760 756.630 2379.900 ;
        RECT 713.085 2379.715 713.375 2379.760 ;
        RECT 756.310 2379.700 756.630 2379.760 ;
        RECT 330.810 2377.860 331.130 2377.920 ;
        RECT 713.085 2377.860 713.375 2377.905 ;
        RECT 330.810 2377.720 713.375 2377.860 ;
        RECT 330.810 2377.660 331.130 2377.720 ;
        RECT 713.085 2377.675 713.375 2377.720 ;
      LAYER via ;
        RECT 756.340 2379.700 756.600 2379.960 ;
        RECT 330.840 2377.660 331.100 2377.920 ;
      LAYER met2 ;
        RECT 756.340 2379.670 756.600 2379.990 ;
        RECT 330.840 2377.630 331.100 2377.950 ;
        RECT 756.400 2377.880 756.540 2379.670 ;
        RECT 330.900 16.900 331.040 2377.630 ;
        RECT 756.380 2373.880 756.660 2377.880 ;
        RECT 329.980 16.760 331.040 16.900 ;
        RECT 329.980 2.400 330.120 16.760 ;
        RECT 329.770 -4.800 330.330 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1072.330 2388.400 1072.650 2388.460 ;
        RECT 1277.030 2388.400 1277.350 2388.460 ;
        RECT 1072.330 2388.260 1277.350 2388.400 ;
        RECT 1072.330 2388.200 1072.650 2388.260 ;
        RECT 1277.030 2388.200 1277.350 2388.260 ;
        RECT 347.370 16.900 347.690 16.960 ;
        RECT 351.510 16.900 351.830 16.960 ;
        RECT 347.370 16.760 351.830 16.900 ;
        RECT 347.370 16.700 347.690 16.760 ;
        RECT 351.510 16.700 351.830 16.760 ;
      LAYER via ;
        RECT 1072.360 2388.200 1072.620 2388.460 ;
        RECT 1277.060 2388.200 1277.320 2388.460 ;
        RECT 347.400 16.700 347.660 16.960 ;
        RECT 351.540 16.700 351.800 16.960 ;
      LAYER met2 ;
        RECT 1072.360 2388.170 1072.620 2388.490 ;
        RECT 1277.060 2388.170 1277.320 2388.490 ;
        RECT 1072.420 2380.525 1072.560 2388.170 ;
        RECT 351.530 2380.155 351.810 2380.525 ;
        RECT 1072.350 2380.155 1072.630 2380.525 ;
        RECT 351.600 16.990 351.740 2380.155 ;
        RECT 1277.120 2377.880 1277.260 2388.170 ;
        RECT 1277.100 2373.880 1277.380 2377.880 ;
        RECT 347.400 16.670 347.660 16.990 ;
        RECT 351.540 16.670 351.800 16.990 ;
        RECT 347.460 2.400 347.600 16.670 ;
        RECT 347.250 -4.800 347.810 2.400 ;
      LAYER via2 ;
        RECT 351.530 2380.200 351.810 2380.480 ;
        RECT 1072.350 2380.200 1072.630 2380.480 ;
      LAYER met3 ;
        RECT 351.505 2380.490 351.835 2380.505 ;
        RECT 1072.325 2380.490 1072.655 2380.505 ;
        RECT 351.505 2380.190 1072.655 2380.490 ;
        RECT 351.505 2380.175 351.835 2380.190 ;
        RECT 1072.325 2380.175 1072.655 2380.190 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 365.310 2375.480 365.630 2375.540 ;
        RECT 807.370 2375.480 807.690 2375.540 ;
        RECT 365.310 2375.340 807.690 2375.480 ;
        RECT 365.310 2375.280 365.630 2375.340 ;
        RECT 807.370 2375.280 807.690 2375.340 ;
      LAYER via ;
        RECT 365.340 2375.280 365.600 2375.540 ;
        RECT 807.400 2375.280 807.660 2375.540 ;
      LAYER met2 ;
        RECT 807.900 2375.650 808.180 2377.880 ;
        RECT 807.460 2375.570 808.180 2375.650 ;
        RECT 365.340 2375.250 365.600 2375.570 ;
        RECT 807.400 2375.510 808.180 2375.570 ;
        RECT 807.400 2375.250 807.660 2375.510 ;
        RECT 365.400 2.400 365.540 2375.250 ;
        RECT 807.900 2373.880 808.180 2375.510 ;
        RECT 365.190 -4.800 365.750 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1048.945 2390.965 1049.115 2392.495 ;
        RECT 1096.785 2390.965 1096.955 2392.495 ;
        RECT 1145.545 2390.965 1145.715 2392.495 ;
        RECT 1193.385 2390.965 1193.555 2392.495 ;
        RECT 1242.145 2390.965 1242.315 2392.495 ;
        RECT 1289.985 2390.965 1290.155 2392.495 ;
        RECT 1634.065 2391.985 1635.615 2392.155 ;
        RECT 1338.745 2390.285 1338.915 2391.135 ;
        RECT 1410.965 2390.285 1411.135 2391.135 ;
        RECT 1435.345 2389.945 1435.515 2391.135 ;
        RECT 1483.185 2389.945 1483.355 2391.135 ;
        RECT 1531.945 2389.945 1532.115 2391.135 ;
        RECT 1579.785 2389.605 1579.955 2391.135 ;
        RECT 1634.065 2390.965 1634.235 2391.985 ;
        RECT 727.405 2380.085 727.575 2380.935 ;
      LAYER mcon ;
        RECT 1048.945 2392.325 1049.115 2392.495 ;
        RECT 1096.785 2392.325 1096.955 2392.495 ;
        RECT 1145.545 2392.325 1145.715 2392.495 ;
        RECT 1193.385 2392.325 1193.555 2392.495 ;
        RECT 1242.145 2392.325 1242.315 2392.495 ;
        RECT 1289.985 2392.325 1290.155 2392.495 ;
        RECT 1635.445 2391.985 1635.615 2392.155 ;
        RECT 1338.745 2390.965 1338.915 2391.135 ;
        RECT 1410.965 2390.965 1411.135 2391.135 ;
        RECT 1435.345 2390.965 1435.515 2391.135 ;
        RECT 1483.185 2390.965 1483.355 2391.135 ;
        RECT 1531.945 2390.965 1532.115 2391.135 ;
        RECT 1579.785 2390.965 1579.955 2391.135 ;
        RECT 727.405 2380.765 727.575 2380.935 ;
      LAYER met1 ;
        RECT 1048.885 2392.480 1049.175 2392.525 ;
        RECT 1096.725 2392.480 1097.015 2392.525 ;
        RECT 1048.885 2392.340 1097.015 2392.480 ;
        RECT 1048.885 2392.295 1049.175 2392.340 ;
        RECT 1096.725 2392.295 1097.015 2392.340 ;
        RECT 1145.485 2392.480 1145.775 2392.525 ;
        RECT 1193.325 2392.480 1193.615 2392.525 ;
        RECT 1145.485 2392.340 1193.615 2392.480 ;
        RECT 1145.485 2392.295 1145.775 2392.340 ;
        RECT 1193.325 2392.295 1193.615 2392.340 ;
        RECT 1242.085 2392.480 1242.375 2392.525 ;
        RECT 1289.925 2392.480 1290.215 2392.525 ;
        RECT 1242.085 2392.340 1290.215 2392.480 ;
        RECT 1242.085 2392.295 1242.375 2392.340 ;
        RECT 1289.925 2392.295 1290.215 2392.340 ;
        RECT 1635.385 2392.140 1635.675 2392.185 ;
        RECT 1646.870 2392.140 1647.190 2392.200 ;
        RECT 1635.385 2392.000 1647.190 2392.140 ;
        RECT 1635.385 2391.955 1635.675 2392.000 ;
        RECT 1646.870 2391.940 1647.190 2392.000 ;
        RECT 1035.070 2391.120 1035.390 2391.180 ;
        RECT 1048.885 2391.120 1049.175 2391.165 ;
        RECT 1035.070 2390.980 1049.175 2391.120 ;
        RECT 1035.070 2390.920 1035.390 2390.980 ;
        RECT 1048.885 2390.935 1049.175 2390.980 ;
        RECT 1096.725 2391.120 1097.015 2391.165 ;
        RECT 1145.485 2391.120 1145.775 2391.165 ;
        RECT 1096.725 2390.980 1145.775 2391.120 ;
        RECT 1096.725 2390.935 1097.015 2390.980 ;
        RECT 1145.485 2390.935 1145.775 2390.980 ;
        RECT 1193.325 2391.120 1193.615 2391.165 ;
        RECT 1242.085 2391.120 1242.375 2391.165 ;
        RECT 1193.325 2390.980 1242.375 2391.120 ;
        RECT 1193.325 2390.935 1193.615 2390.980 ;
        RECT 1242.085 2390.935 1242.375 2390.980 ;
        RECT 1289.925 2391.120 1290.215 2391.165 ;
        RECT 1338.685 2391.120 1338.975 2391.165 ;
        RECT 1289.925 2390.980 1338.975 2391.120 ;
        RECT 1289.925 2390.935 1290.215 2390.980 ;
        RECT 1338.685 2390.935 1338.975 2390.980 ;
        RECT 1410.905 2391.120 1411.195 2391.165 ;
        RECT 1435.285 2391.120 1435.575 2391.165 ;
        RECT 1410.905 2390.980 1435.575 2391.120 ;
        RECT 1410.905 2390.935 1411.195 2390.980 ;
        RECT 1435.285 2390.935 1435.575 2390.980 ;
        RECT 1483.125 2391.120 1483.415 2391.165 ;
        RECT 1531.885 2391.120 1532.175 2391.165 ;
        RECT 1483.125 2390.980 1532.175 2391.120 ;
        RECT 1483.125 2390.935 1483.415 2390.980 ;
        RECT 1531.885 2390.935 1532.175 2390.980 ;
        RECT 1579.725 2391.120 1580.015 2391.165 ;
        RECT 1634.005 2391.120 1634.295 2391.165 ;
        RECT 1579.725 2390.980 1634.295 2391.120 ;
        RECT 1579.725 2390.935 1580.015 2390.980 ;
        RECT 1634.005 2390.935 1634.295 2390.980 ;
        RECT 1338.685 2390.440 1338.975 2390.485 ;
        RECT 1410.905 2390.440 1411.195 2390.485 ;
        RECT 1338.685 2390.300 1411.195 2390.440 ;
        RECT 1338.685 2390.255 1338.975 2390.300 ;
        RECT 1410.905 2390.255 1411.195 2390.300 ;
        RECT 1435.285 2390.100 1435.575 2390.145 ;
        RECT 1483.125 2390.100 1483.415 2390.145 ;
        RECT 1435.285 2389.960 1483.415 2390.100 ;
        RECT 1435.285 2389.915 1435.575 2389.960 ;
        RECT 1483.125 2389.915 1483.415 2389.960 ;
        RECT 1531.885 2390.100 1532.175 2390.145 ;
        RECT 1531.885 2389.960 1539.000 2390.100 ;
        RECT 1531.885 2389.915 1532.175 2389.960 ;
        RECT 1538.860 2389.760 1539.000 2389.960 ;
        RECT 1579.725 2389.760 1580.015 2389.805 ;
        RECT 1538.860 2389.620 1580.015 2389.760 ;
        RECT 1579.725 2389.575 1580.015 2389.620 ;
        RECT 718.130 2380.920 718.450 2380.980 ;
        RECT 727.345 2380.920 727.635 2380.965 ;
        RECT 718.130 2380.780 727.635 2380.920 ;
        RECT 718.130 2380.720 718.450 2380.780 ;
        RECT 727.345 2380.735 727.635 2380.780 ;
        RECT 727.345 2380.240 727.635 2380.285 ;
        RECT 1035.070 2380.240 1035.390 2380.300 ;
        RECT 727.345 2380.100 1035.390 2380.240 ;
        RECT 727.345 2380.055 727.635 2380.100 ;
        RECT 1035.070 2380.040 1035.390 2380.100 ;
        RECT 383.250 16.900 383.570 16.960 ;
        RECT 386.010 16.900 386.330 16.960 ;
        RECT 383.250 16.760 386.330 16.900 ;
        RECT 383.250 16.700 383.570 16.760 ;
        RECT 386.010 16.700 386.330 16.760 ;
      LAYER via ;
        RECT 1646.900 2391.940 1647.160 2392.200 ;
        RECT 1035.100 2390.920 1035.360 2391.180 ;
        RECT 718.160 2380.720 718.420 2380.980 ;
        RECT 1035.100 2380.040 1035.360 2380.300 ;
        RECT 383.280 16.700 383.540 16.960 ;
        RECT 386.040 16.700 386.300 16.960 ;
      LAYER met2 ;
        RECT 1646.900 2391.910 1647.160 2392.230 ;
        RECT 1035.100 2390.890 1035.360 2391.210 ;
        RECT 718.160 2380.690 718.420 2381.010 ;
        RECT 718.220 2374.405 718.360 2380.690 ;
        RECT 1035.160 2380.330 1035.300 2390.890 ;
        RECT 1035.100 2380.010 1035.360 2380.330 ;
        RECT 1646.960 2377.880 1647.100 2391.910 ;
        RECT 386.030 2374.035 386.310 2374.405 ;
        RECT 718.150 2374.035 718.430 2374.405 ;
        RECT 386.100 16.990 386.240 2374.035 ;
        RECT 1646.940 2373.880 1647.220 2377.880 ;
        RECT 383.280 16.670 383.540 16.990 ;
        RECT 386.040 16.670 386.300 16.990 ;
        RECT 383.340 2.400 383.480 16.670 ;
        RECT 383.130 -4.800 383.690 2.400 ;
      LAYER via2 ;
        RECT 386.030 2374.080 386.310 2374.360 ;
        RECT 718.150 2374.080 718.430 2374.360 ;
      LAYER met3 ;
        RECT 386.005 2374.370 386.335 2374.385 ;
        RECT 718.125 2374.370 718.455 2374.385 ;
        RECT 386.005 2374.070 718.455 2374.370 ;
        RECT 386.005 2374.055 386.335 2374.070 ;
        RECT 718.125 2374.055 718.455 2374.070 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1024.030 2388.060 1024.350 2388.120 ;
        RECT 1421.470 2388.060 1421.790 2388.120 ;
        RECT 1024.030 2387.920 1421.790 2388.060 ;
        RECT 1024.030 2387.860 1024.350 2387.920 ;
        RECT 1421.470 2387.860 1421.790 2387.920 ;
        RECT 401.190 16.900 401.510 16.960 ;
        RECT 406.710 16.900 407.030 16.960 ;
        RECT 401.190 16.760 407.030 16.900 ;
        RECT 401.190 16.700 401.510 16.760 ;
        RECT 406.710 16.700 407.030 16.760 ;
      LAYER via ;
        RECT 1024.060 2387.860 1024.320 2388.120 ;
        RECT 1421.500 2387.860 1421.760 2388.120 ;
        RECT 401.220 16.700 401.480 16.960 ;
        RECT 406.740 16.700 407.000 16.960 ;
      LAYER met2 ;
        RECT 1024.060 2387.830 1024.320 2388.150 ;
        RECT 1421.500 2387.830 1421.760 2388.150 ;
        RECT 1024.120 2378.485 1024.260 2387.830 ;
        RECT 406.730 2378.115 407.010 2378.485 ;
        RECT 1024.050 2378.115 1024.330 2378.485 ;
        RECT 406.800 16.990 406.940 2378.115 ;
        RECT 1421.560 2377.880 1421.700 2387.830 ;
        RECT 1421.540 2373.880 1421.820 2377.880 ;
        RECT 401.220 16.670 401.480 16.990 ;
        RECT 406.740 16.670 407.000 16.990 ;
        RECT 401.280 2.400 401.420 16.670 ;
        RECT 401.070 -4.800 401.630 2.400 ;
      LAYER via2 ;
        RECT 406.730 2378.160 407.010 2378.440 ;
        RECT 1024.050 2378.160 1024.330 2378.440 ;
      LAYER met3 ;
        RECT 406.705 2378.450 407.035 2378.465 ;
        RECT 1024.025 2378.450 1024.355 2378.465 ;
        RECT 406.705 2378.150 1024.355 2378.450 ;
        RECT 406.705 2378.135 407.035 2378.150 ;
        RECT 1024.025 2378.135 1024.355 2378.150 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 62.170 17.920 62.490 17.980 ;
        RECT 68.610 17.920 68.930 17.980 ;
        RECT 62.170 17.780 68.930 17.920 ;
        RECT 62.170 17.720 62.490 17.780 ;
        RECT 68.610 17.720 68.930 17.780 ;
      LAYER via ;
        RECT 62.200 17.720 62.460 17.980 ;
        RECT 68.640 17.720 68.900 17.980 ;
      LAYER met2 ;
        RECT 68.630 887.555 68.910 887.925 ;
        RECT 68.700 18.010 68.840 887.555 ;
        RECT 62.200 17.690 62.460 18.010 ;
        RECT 68.640 17.690 68.900 18.010 ;
        RECT 62.260 2.400 62.400 17.690 ;
        RECT 62.050 -4.800 62.610 2.400 ;
      LAYER via2 ;
        RECT 68.630 887.600 68.910 887.880 ;
      LAYER met3 ;
        RECT 1755.835 1561.770 1759.835 1561.775 ;
        RECT 1771.270 1561.770 1771.650 1561.780 ;
        RECT 1755.835 1561.470 1771.650 1561.770 ;
        RECT 1755.835 1561.175 1759.835 1561.470 ;
        RECT 1771.270 1561.460 1771.650 1561.470 ;
        RECT 68.605 887.890 68.935 887.905 ;
        RECT 1771.270 887.890 1771.650 887.900 ;
        RECT 68.605 887.590 1771.650 887.890 ;
        RECT 68.605 887.575 68.935 887.590 ;
        RECT 1771.270 887.580 1771.650 887.590 ;
      LAYER via3 ;
        RECT 1771.300 1561.460 1771.620 1561.780 ;
        RECT 1771.300 887.580 1771.620 887.900 ;
      LAYER met4 ;
        RECT 1771.295 1561.455 1771.625 1561.785 ;
        RECT 1771.310 887.905 1771.610 1561.455 ;
        RECT 1771.295 887.575 1771.625 887.905 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 420.510 1313.660 420.830 1313.720 ;
        RECT 1070.950 1313.660 1071.270 1313.720 ;
        RECT 420.510 1313.520 1071.270 1313.660 ;
        RECT 420.510 1313.460 420.830 1313.520 ;
        RECT 1070.950 1313.460 1071.270 1313.520 ;
      LAYER via ;
        RECT 420.540 1313.460 420.800 1313.720 ;
        RECT 1070.980 1313.460 1071.240 1313.720 ;
      LAYER met2 ;
        RECT 1071.020 1323.135 1071.300 1327.135 ;
        RECT 1071.040 1313.750 1071.180 1323.135 ;
        RECT 420.540 1313.430 420.800 1313.750 ;
        RECT 1070.980 1313.430 1071.240 1313.750 ;
        RECT 420.600 17.410 420.740 1313.430 ;
        RECT 419.220 17.270 420.740 17.410 ;
        RECT 419.220 2.400 419.360 17.270 ;
        RECT 419.010 -4.800 419.570 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 441.210 1794.080 441.530 1794.140 ;
        RECT 705.250 1794.080 705.570 1794.140 ;
        RECT 441.210 1793.940 705.570 1794.080 ;
        RECT 441.210 1793.880 441.530 1793.940 ;
        RECT 705.250 1793.880 705.570 1793.940 ;
        RECT 436.610 16.900 436.930 16.960 ;
        RECT 441.210 16.900 441.530 16.960 ;
        RECT 436.610 16.760 441.530 16.900 ;
        RECT 436.610 16.700 436.930 16.760 ;
        RECT 441.210 16.700 441.530 16.760 ;
      LAYER via ;
        RECT 441.240 1793.880 441.500 1794.140 ;
        RECT 705.280 1793.880 705.540 1794.140 ;
        RECT 436.640 16.700 436.900 16.960 ;
        RECT 441.240 16.700 441.500 16.960 ;
      LAYER met2 ;
        RECT 705.270 1796.715 705.550 1797.085 ;
        RECT 705.340 1794.170 705.480 1796.715 ;
        RECT 441.240 1793.850 441.500 1794.170 ;
        RECT 705.280 1793.850 705.540 1794.170 ;
        RECT 441.300 16.990 441.440 1793.850 ;
        RECT 436.640 16.670 436.900 16.990 ;
        RECT 441.240 16.670 441.500 16.990 ;
        RECT 436.700 2.400 436.840 16.670 ;
        RECT 436.490 -4.800 437.050 2.400 ;
      LAYER via2 ;
        RECT 705.270 1796.760 705.550 1797.040 ;
      LAYER met3 ;
        RECT 705.245 1797.050 705.575 1797.065 ;
        RECT 715.810 1797.050 719.810 1797.055 ;
        RECT 705.245 1796.750 719.810 1797.050 ;
        RECT 705.245 1796.735 705.575 1796.750 ;
        RECT 715.810 1796.455 719.810 1796.750 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 454.550 1911.380 454.870 1911.440 ;
        RECT 706.170 1911.380 706.490 1911.440 ;
        RECT 454.550 1911.240 706.490 1911.380 ;
        RECT 454.550 1911.180 454.870 1911.240 ;
        RECT 706.170 1911.180 706.490 1911.240 ;
      LAYER via ;
        RECT 454.580 1911.180 454.840 1911.440 ;
        RECT 706.200 1911.180 706.460 1911.440 ;
      LAYER met2 ;
        RECT 706.190 1916.395 706.470 1916.765 ;
        RECT 706.260 1911.470 706.400 1916.395 ;
        RECT 454.580 1911.150 454.840 1911.470 ;
        RECT 706.200 1911.150 706.460 1911.470 ;
        RECT 454.640 2.400 454.780 1911.150 ;
        RECT 454.430 -4.800 454.990 2.400 ;
      LAYER via2 ;
        RECT 706.190 1916.440 706.470 1916.720 ;
      LAYER met3 ;
        RECT 706.165 1916.730 706.495 1916.745 ;
        RECT 715.810 1916.730 719.810 1916.735 ;
        RECT 706.165 1916.430 719.810 1916.730 ;
        RECT 706.165 1916.415 706.495 1916.430 ;
        RECT 715.810 1916.135 719.810 1916.430 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 475.710 1711.460 476.030 1711.520 ;
        RECT 710.310 1711.460 710.630 1711.520 ;
        RECT 475.710 1711.320 710.630 1711.460 ;
        RECT 475.710 1711.260 476.030 1711.320 ;
        RECT 710.310 1711.260 710.630 1711.320 ;
        RECT 472.490 16.900 472.810 16.960 ;
        RECT 475.710 16.900 476.030 16.960 ;
        RECT 472.490 16.760 476.030 16.900 ;
        RECT 472.490 16.700 472.810 16.760 ;
        RECT 475.710 16.700 476.030 16.760 ;
      LAYER via ;
        RECT 475.740 1711.260 476.000 1711.520 ;
        RECT 710.340 1711.260 710.600 1711.520 ;
        RECT 472.520 16.700 472.780 16.960 ;
        RECT 475.740 16.700 476.000 16.960 ;
      LAYER met2 ;
        RECT 475.740 1711.230 476.000 1711.550 ;
        RECT 710.340 1711.405 710.600 1711.550 ;
        RECT 475.800 16.990 475.940 1711.230 ;
        RECT 710.330 1711.035 710.610 1711.405 ;
        RECT 472.520 16.670 472.780 16.990 ;
        RECT 475.740 16.670 476.000 16.990 ;
        RECT 472.580 2.400 472.720 16.670 ;
        RECT 472.370 -4.800 472.930 2.400 ;
      LAYER via2 ;
        RECT 710.330 1711.080 710.610 1711.360 ;
      LAYER met3 ;
        RECT 710.305 1711.370 710.635 1711.385 ;
        RECT 715.810 1711.370 719.810 1711.375 ;
        RECT 710.305 1711.070 719.810 1711.370 ;
        RECT 710.305 1711.055 710.635 1711.070 ;
        RECT 715.810 1710.775 719.810 1711.070 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 976.265 2388.245 976.435 2394.195 ;
      LAYER mcon ;
        RECT 976.265 2394.025 976.435 2394.195 ;
      LAYER met1 ;
        RECT 976.205 2394.180 976.495 2394.225 ;
        RECT 1230.110 2394.180 1230.430 2394.240 ;
        RECT 976.205 2394.040 1230.430 2394.180 ;
        RECT 976.205 2393.995 976.495 2394.040 ;
        RECT 1230.110 2393.980 1230.430 2394.040 ;
        RECT 931.570 2388.400 931.890 2388.460 ;
        RECT 976.205 2388.400 976.495 2388.445 ;
        RECT 931.570 2388.260 976.495 2388.400 ;
        RECT 931.570 2388.200 931.890 2388.260 ;
        RECT 976.205 2388.215 976.495 2388.260 ;
        RECT 579.670 2378.200 579.990 2378.260 ;
        RECT 627.510 2378.200 627.830 2378.260 ;
        RECT 579.670 2378.060 627.830 2378.200 ;
        RECT 579.670 2378.000 579.990 2378.060 ;
        RECT 627.510 2378.000 627.830 2378.060 ;
        RECT 855.670 2377.520 855.990 2377.580 ;
        RECT 884.650 2377.520 884.970 2377.580 ;
        RECT 855.670 2377.380 884.970 2377.520 ;
        RECT 855.670 2377.320 855.990 2377.380 ;
        RECT 884.650 2377.320 884.970 2377.380 ;
        RECT 927.430 2377.180 927.750 2377.240 ;
        RECT 931.570 2377.180 931.890 2377.240 ;
        RECT 927.430 2377.040 931.890 2377.180 ;
        RECT 927.430 2376.980 927.750 2377.040 ;
        RECT 931.570 2376.980 931.890 2377.040 ;
        RECT 782.990 2375.140 783.310 2375.200 ;
        RECT 786.670 2375.140 786.990 2375.200 ;
        RECT 782.990 2375.000 786.990 2375.140 ;
        RECT 782.990 2374.940 783.310 2375.000 ;
        RECT 786.670 2374.940 786.990 2375.000 ;
        RECT 490.430 16.900 490.750 16.960 ;
        RECT 496.410 16.900 496.730 16.960 ;
        RECT 490.430 16.760 496.730 16.900 ;
        RECT 490.430 16.700 490.750 16.760 ;
        RECT 496.410 16.700 496.730 16.760 ;
      LAYER via ;
        RECT 1230.140 2393.980 1230.400 2394.240 ;
        RECT 931.600 2388.200 931.860 2388.460 ;
        RECT 579.700 2378.000 579.960 2378.260 ;
        RECT 627.540 2378.000 627.800 2378.260 ;
        RECT 855.700 2377.320 855.960 2377.580 ;
        RECT 884.680 2377.320 884.940 2377.580 ;
        RECT 927.460 2376.980 927.720 2377.240 ;
        RECT 931.600 2376.980 931.860 2377.240 ;
        RECT 783.020 2374.940 783.280 2375.200 ;
        RECT 786.700 2374.940 786.960 2375.200 ;
        RECT 490.460 16.700 490.720 16.960 ;
        RECT 496.440 16.700 496.700 16.960 ;
      LAYER met2 ;
        RECT 1230.140 2393.950 1230.400 2394.270 ;
        RECT 931.600 2388.170 931.860 2388.490 ;
        RECT 579.700 2377.970 579.960 2378.290 ;
        RECT 627.540 2377.970 627.800 2378.290 ;
        RECT 579.760 2377.805 579.900 2377.970 ;
        RECT 496.430 2377.435 496.710 2377.805 ;
        RECT 579.690 2377.435 579.970 2377.805 ;
        RECT 496.500 16.990 496.640 2377.435 ;
        RECT 544.730 2377.010 545.010 2377.125 ;
        RECT 544.730 2376.870 545.400 2377.010 ;
        RECT 544.730 2376.755 545.010 2376.870 ;
        RECT 545.260 2376.445 545.400 2376.870 ;
        RECT 627.600 2376.445 627.740 2377.970 ;
        RECT 855.700 2377.290 855.960 2377.610 ;
        RECT 884.680 2377.290 884.940 2377.610 ;
        RECT 855.760 2377.125 855.900 2377.290 ;
        RECT 884.740 2377.125 884.880 2377.290 ;
        RECT 931.660 2377.270 931.800 2388.170 ;
        RECT 1230.200 2377.880 1230.340 2393.950 ;
        RECT 927.460 2377.125 927.720 2377.270 ;
        RECT 783.010 2376.755 783.290 2377.125 ;
        RECT 786.690 2376.755 786.970 2377.125 ;
        RECT 855.690 2376.755 855.970 2377.125 ;
        RECT 884.670 2376.755 884.950 2377.125 ;
        RECT 927.450 2376.755 927.730 2377.125 ;
        RECT 931.600 2376.950 931.860 2377.270 ;
        RECT 545.190 2376.075 545.470 2376.445 ;
        RECT 627.530 2376.075 627.810 2376.445 ;
        RECT 783.080 2375.230 783.220 2376.755 ;
        RECT 786.760 2375.230 786.900 2376.755 ;
        RECT 783.020 2374.910 783.280 2375.230 ;
        RECT 786.700 2374.910 786.960 2375.230 ;
        RECT 1230.180 2373.880 1230.460 2377.880 ;
        RECT 490.460 16.670 490.720 16.990 ;
        RECT 496.440 16.670 496.700 16.990 ;
        RECT 490.520 2.400 490.660 16.670 ;
        RECT 490.310 -4.800 490.870 2.400 ;
      LAYER via2 ;
        RECT 496.430 2377.480 496.710 2377.760 ;
        RECT 579.690 2377.480 579.970 2377.760 ;
        RECT 544.730 2376.800 545.010 2377.080 ;
        RECT 783.010 2376.800 783.290 2377.080 ;
        RECT 786.690 2376.800 786.970 2377.080 ;
        RECT 855.690 2376.800 855.970 2377.080 ;
        RECT 884.670 2376.800 884.950 2377.080 ;
        RECT 927.450 2376.800 927.730 2377.080 ;
        RECT 545.190 2376.120 545.470 2376.400 ;
        RECT 627.530 2376.120 627.810 2376.400 ;
      LAYER met3 ;
        RECT 496.405 2377.770 496.735 2377.785 ;
        RECT 579.665 2377.770 579.995 2377.785 ;
        RECT 496.405 2377.470 497.410 2377.770 ;
        RECT 496.405 2377.455 496.735 2377.470 ;
        RECT 497.110 2377.090 497.410 2377.470 ;
        RECT 578.990 2377.470 579.995 2377.770 ;
        RECT 544.705 2377.090 545.035 2377.105 ;
        RECT 497.110 2376.790 545.035 2377.090 ;
        RECT 544.705 2376.775 545.035 2376.790 ;
        RECT 545.165 2376.410 545.495 2376.425 ;
        RECT 578.990 2376.410 579.290 2377.470 ;
        RECT 579.665 2377.455 579.995 2377.470 ;
        RECT 782.985 2377.090 783.315 2377.105 ;
        RECT 716.990 2376.790 783.315 2377.090 ;
        RECT 545.165 2376.110 579.290 2376.410 ;
        RECT 627.505 2376.410 627.835 2376.425 ;
        RECT 716.990 2376.410 717.290 2376.790 ;
        RECT 782.985 2376.775 783.315 2376.790 ;
        RECT 786.665 2377.090 786.995 2377.105 ;
        RECT 820.910 2377.090 821.290 2377.100 ;
        RECT 786.665 2376.790 821.290 2377.090 ;
        RECT 786.665 2376.775 786.995 2376.790 ;
        RECT 820.910 2376.780 821.290 2376.790 ;
        RECT 822.750 2377.090 823.130 2377.100 ;
        RECT 855.665 2377.090 855.995 2377.105 ;
        RECT 822.750 2376.790 855.995 2377.090 ;
        RECT 822.750 2376.780 823.130 2376.790 ;
        RECT 855.665 2376.775 855.995 2376.790 ;
        RECT 884.645 2377.090 884.975 2377.105 ;
        RECT 927.425 2377.090 927.755 2377.105 ;
        RECT 884.645 2376.790 927.755 2377.090 ;
        RECT 884.645 2376.775 884.975 2376.790 ;
        RECT 927.425 2376.775 927.755 2376.790 ;
        RECT 627.505 2376.110 717.290 2376.410 ;
        RECT 545.165 2376.095 545.495 2376.110 ;
        RECT 627.505 2376.095 627.835 2376.110 ;
      LAYER via3 ;
        RECT 820.940 2376.780 821.260 2377.100 ;
        RECT 822.780 2376.780 823.100 2377.100 ;
      LAYER met4 ;
        RECT 820.950 2378.150 823.090 2378.450 ;
        RECT 820.950 2377.105 821.250 2378.150 ;
        RECT 822.790 2377.105 823.090 2378.150 ;
        RECT 820.935 2376.775 821.265 2377.105 ;
        RECT 822.775 2376.775 823.105 2377.105 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 510.210 2382.280 510.530 2382.340 ;
        RECT 1675.390 2382.280 1675.710 2382.340 ;
        RECT 510.210 2382.140 1675.710 2382.280 ;
        RECT 510.210 2382.080 510.530 2382.140 ;
        RECT 1675.390 2382.080 1675.710 2382.140 ;
        RECT 507.910 16.900 508.230 16.960 ;
        RECT 510.210 16.900 510.530 16.960 ;
        RECT 507.910 16.760 510.530 16.900 ;
        RECT 507.910 16.700 508.230 16.760 ;
        RECT 510.210 16.700 510.530 16.760 ;
      LAYER via ;
        RECT 510.240 2382.080 510.500 2382.340 ;
        RECT 1675.420 2382.080 1675.680 2382.340 ;
        RECT 507.940 16.700 508.200 16.960 ;
        RECT 510.240 16.700 510.500 16.960 ;
      LAYER met2 ;
        RECT 510.240 2382.050 510.500 2382.370 ;
        RECT 1675.420 2382.050 1675.680 2382.370 ;
        RECT 510.300 16.990 510.440 2382.050 ;
        RECT 1675.480 2377.880 1675.620 2382.050 ;
        RECT 1675.460 2373.880 1675.740 2377.880 ;
        RECT 507.940 16.670 508.200 16.990 ;
        RECT 510.240 16.670 510.500 16.990 ;
        RECT 508.000 2.400 508.140 16.670 ;
        RECT 507.790 -4.800 508.350 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 530.450 1960.000 530.770 1960.060 ;
        RECT 710.310 1960.000 710.630 1960.060 ;
        RECT 530.450 1959.860 710.630 1960.000 ;
        RECT 530.450 1959.800 530.770 1959.860 ;
        RECT 710.310 1959.800 710.630 1959.860 ;
        RECT 525.850 17.240 526.170 17.300 ;
        RECT 530.450 17.240 530.770 17.300 ;
        RECT 525.850 17.100 530.770 17.240 ;
        RECT 525.850 17.040 526.170 17.100 ;
        RECT 530.450 17.040 530.770 17.100 ;
      LAYER via ;
        RECT 530.480 1959.800 530.740 1960.060 ;
        RECT 710.340 1959.800 710.600 1960.060 ;
        RECT 525.880 17.040 526.140 17.300 ;
        RECT 530.480 17.040 530.740 17.300 ;
      LAYER met2 ;
        RECT 530.480 1959.770 530.740 1960.090 ;
        RECT 710.330 1959.915 710.610 1960.285 ;
        RECT 710.340 1959.770 710.600 1959.915 ;
        RECT 530.540 17.330 530.680 1959.770 ;
        RECT 525.880 17.010 526.140 17.330 ;
        RECT 530.480 17.010 530.740 17.330 ;
        RECT 525.940 2.400 526.080 17.010 ;
        RECT 525.730 -4.800 526.290 2.400 ;
      LAYER via2 ;
        RECT 710.330 1959.960 710.610 1960.240 ;
      LAYER met3 ;
        RECT 710.305 1960.250 710.635 1960.265 ;
        RECT 715.810 1960.250 719.810 1960.255 ;
        RECT 710.305 1959.950 719.810 1960.250 ;
        RECT 710.305 1959.935 710.635 1959.950 ;
        RECT 715.810 1959.655 719.810 1959.950 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 544.710 1359.560 545.030 1359.620 ;
        RECT 701.570 1359.560 701.890 1359.620 ;
        RECT 544.710 1359.420 701.890 1359.560 ;
        RECT 544.710 1359.360 545.030 1359.420 ;
        RECT 701.570 1359.360 701.890 1359.420 ;
      LAYER via ;
        RECT 544.740 1359.360 545.000 1359.620 ;
        RECT 701.600 1359.360 701.860 1359.620 ;
      LAYER met2 ;
        RECT 701.590 1361.515 701.870 1361.885 ;
        RECT 701.660 1359.650 701.800 1361.515 ;
        RECT 544.740 1359.330 545.000 1359.650 ;
        RECT 701.600 1359.330 701.860 1359.650 ;
        RECT 544.800 16.900 544.940 1359.330 ;
        RECT 543.880 16.760 544.940 16.900 ;
        RECT 543.880 2.400 544.020 16.760 ;
        RECT 543.670 -4.800 544.230 2.400 ;
      LAYER via2 ;
        RECT 701.590 1361.560 701.870 1361.840 ;
      LAYER met3 ;
        RECT 701.565 1361.850 701.895 1361.865 ;
        RECT 715.810 1361.850 719.810 1361.855 ;
        RECT 701.565 1361.550 719.810 1361.850 ;
        RECT 701.565 1361.535 701.895 1361.550 ;
        RECT 715.810 1361.255 719.810 1361.550 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 561.730 39.680 562.050 39.740 ;
        RECT 1768.310 39.680 1768.630 39.740 ;
        RECT 561.730 39.540 1768.630 39.680 ;
        RECT 561.730 39.480 562.050 39.540 ;
        RECT 1768.310 39.480 1768.630 39.540 ;
      LAYER via ;
        RECT 561.760 39.480 562.020 39.740 ;
        RECT 1768.340 39.480 1768.600 39.740 ;
      LAYER met2 ;
        RECT 1768.330 1365.595 1768.610 1365.965 ;
        RECT 1768.400 39.770 1768.540 1365.595 ;
        RECT 561.760 39.450 562.020 39.770 ;
        RECT 1768.340 39.450 1768.600 39.770 ;
        RECT 561.820 2.400 561.960 39.450 ;
        RECT 561.610 -4.800 562.170 2.400 ;
      LAYER via2 ;
        RECT 1768.330 1365.640 1768.610 1365.920 ;
      LAYER met3 ;
        RECT 1755.835 1365.930 1759.835 1365.935 ;
        RECT 1768.305 1365.930 1768.635 1365.945 ;
        RECT 1755.835 1365.630 1768.635 1365.930 ;
        RECT 1755.835 1365.335 1759.835 1365.630 ;
        RECT 1768.305 1365.615 1768.635 1365.630 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 579.670 18.260 579.990 18.320 ;
        RECT 585.650 18.260 585.970 18.320 ;
        RECT 579.670 18.120 585.970 18.260 ;
        RECT 579.670 18.060 579.990 18.120 ;
        RECT 585.650 18.060 585.970 18.120 ;
      LAYER via ;
        RECT 579.700 18.060 579.960 18.320 ;
        RECT 585.680 18.060 585.940 18.320 ;
      LAYER met2 ;
        RECT 585.670 81.075 585.950 81.445 ;
        RECT 585.740 18.350 585.880 81.075 ;
        RECT 579.700 18.030 579.960 18.350 ;
        RECT 585.680 18.030 585.940 18.350 ;
        RECT 579.760 2.400 579.900 18.030 ;
        RECT 579.550 -4.800 580.110 2.400 ;
      LAYER via2 ;
        RECT 585.670 81.120 585.950 81.400 ;
      LAYER met3 ;
        RECT 1755.835 2040.490 1759.835 2040.495 ;
        RECT 1760.230 2040.490 1760.610 2040.500 ;
        RECT 1755.835 2040.190 1760.610 2040.490 ;
        RECT 1755.835 2039.895 1759.835 2040.190 ;
        RECT 1760.230 2040.180 1760.610 2040.190 ;
        RECT 585.645 81.410 585.975 81.425 ;
        RECT 1760.230 81.410 1760.610 81.420 ;
        RECT 585.645 81.110 1760.610 81.410 ;
        RECT 585.645 81.095 585.975 81.110 ;
        RECT 1760.230 81.100 1760.610 81.110 ;
      LAYER via3 ;
        RECT 1760.260 2040.180 1760.580 2040.500 ;
        RECT 1760.260 81.100 1760.580 81.420 ;
      LAYER met4 ;
        RECT 1760.255 2040.175 1760.585 2040.505 ;
        RECT 1760.270 81.425 1760.570 2040.175 ;
        RECT 1760.255 81.095 1760.585 81.425 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 868.550 2387.720 868.870 2387.780 ;
        RECT 1212.630 2387.720 1212.950 2387.780 ;
        RECT 868.550 2387.580 1212.950 2387.720 ;
        RECT 868.550 2387.520 868.870 2387.580 ;
        RECT 1212.630 2387.520 1212.950 2387.580 ;
        RECT 89.310 2384.660 89.630 2384.720 ;
        RECT 868.550 2384.660 868.870 2384.720 ;
        RECT 89.310 2384.520 868.870 2384.660 ;
        RECT 89.310 2384.460 89.630 2384.520 ;
        RECT 868.550 2384.460 868.870 2384.520 ;
        RECT 86.090 17.920 86.410 17.980 ;
        RECT 89.310 17.920 89.630 17.980 ;
        RECT 86.090 17.780 89.630 17.920 ;
        RECT 86.090 17.720 86.410 17.780 ;
        RECT 89.310 17.720 89.630 17.780 ;
      LAYER via ;
        RECT 868.580 2387.520 868.840 2387.780 ;
        RECT 1212.660 2387.520 1212.920 2387.780 ;
        RECT 89.340 2384.460 89.600 2384.720 ;
        RECT 868.580 2384.460 868.840 2384.720 ;
        RECT 86.120 17.720 86.380 17.980 ;
        RECT 89.340 17.720 89.600 17.980 ;
      LAYER met2 ;
        RECT 868.580 2387.490 868.840 2387.810 ;
        RECT 1212.660 2387.490 1212.920 2387.810 ;
        RECT 868.640 2384.750 868.780 2387.490 ;
        RECT 89.340 2384.430 89.600 2384.750 ;
        RECT 868.580 2384.430 868.840 2384.750 ;
        RECT 89.400 18.010 89.540 2384.430 ;
        RECT 1212.720 2377.880 1212.860 2387.490 ;
        RECT 1212.700 2373.880 1212.980 2377.880 ;
        RECT 86.120 17.690 86.380 18.010 ;
        RECT 89.340 17.690 89.600 18.010 ;
        RECT 86.180 2.400 86.320 17.690 ;
        RECT 85.970 -4.800 86.530 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 599.910 2391.120 600.230 2391.180 ;
        RECT 1033.230 2391.120 1033.550 2391.180 ;
        RECT 599.910 2390.980 1033.550 2391.120 ;
        RECT 599.910 2390.920 600.230 2390.980 ;
        RECT 1033.230 2390.920 1033.550 2390.980 ;
        RECT 597.150 17.240 597.470 17.300 ;
        RECT 599.910 17.240 600.230 17.300 ;
        RECT 597.150 17.100 600.230 17.240 ;
        RECT 597.150 17.040 597.470 17.100 ;
        RECT 599.910 17.040 600.230 17.100 ;
      LAYER via ;
        RECT 599.940 2390.920 600.200 2391.180 ;
        RECT 1033.260 2390.920 1033.520 2391.180 ;
        RECT 597.180 17.040 597.440 17.300 ;
        RECT 599.940 17.040 600.200 17.300 ;
      LAYER met2 ;
        RECT 599.940 2390.890 600.200 2391.210 ;
        RECT 1033.260 2390.890 1033.520 2391.210 ;
        RECT 600.000 17.330 600.140 2390.890 ;
        RECT 1033.320 2377.880 1033.460 2390.890 ;
        RECT 1033.300 2373.880 1033.580 2377.880 ;
        RECT 597.180 17.010 597.440 17.330 ;
        RECT 599.940 17.010 600.200 17.330 ;
        RECT 597.240 2.400 597.380 17.010 ;
        RECT 597.030 -4.800 597.590 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 615.090 15.200 615.410 15.260 ;
        RECT 620.610 15.200 620.930 15.260 ;
        RECT 615.090 15.060 620.930 15.200 ;
        RECT 615.090 15.000 615.410 15.060 ;
        RECT 620.610 15.000 620.930 15.060 ;
      LAYER via ;
        RECT 615.120 15.000 615.380 15.260 ;
        RECT 620.640 15.000 620.900 15.260 ;
      LAYER met2 ;
        RECT 620.630 81.755 620.910 82.125 ;
        RECT 620.700 15.290 620.840 81.755 ;
        RECT 615.120 14.970 615.380 15.290 ;
        RECT 620.640 14.970 620.900 15.290 ;
        RECT 615.180 2.400 615.320 14.970 ;
        RECT 614.970 -4.800 615.530 2.400 ;
      LAYER via2 ;
        RECT 620.630 81.800 620.910 82.080 ;
      LAYER met3 ;
        RECT 1755.835 2032.330 1759.835 2032.335 ;
        RECT 1766.670 2032.330 1767.050 2032.340 ;
        RECT 1755.835 2032.030 1767.050 2032.330 ;
        RECT 1755.835 2031.735 1759.835 2032.030 ;
        RECT 1766.670 2032.020 1767.050 2032.030 ;
        RECT 620.605 82.090 620.935 82.105 ;
        RECT 1766.670 82.090 1767.050 82.100 ;
        RECT 620.605 81.790 1767.050 82.090 ;
        RECT 620.605 81.775 620.935 81.790 ;
        RECT 1766.670 81.780 1767.050 81.790 ;
      LAYER via3 ;
        RECT 1766.700 2032.020 1767.020 2032.340 ;
        RECT 1766.700 81.780 1767.020 82.100 ;
      LAYER met4 ;
        RECT 1766.695 2032.015 1767.025 2032.345 ;
        RECT 1766.710 82.105 1767.010 2032.015 ;
        RECT 1766.695 81.775 1767.025 82.105 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 109.550 18.260 109.870 18.320 ;
        RECT 175.790 18.260 176.110 18.320 ;
        RECT 109.550 18.120 176.110 18.260 ;
        RECT 109.550 18.060 109.870 18.120 ;
        RECT 175.790 18.060 176.110 18.120 ;
      LAYER via ;
        RECT 109.580 18.060 109.840 18.320 ;
        RECT 175.820 18.060 176.080 18.320 ;
      LAYER met2 ;
        RECT 1447.300 1323.135 1447.580 1327.135 ;
        RECT 1447.320 1314.285 1447.460 1323.135 ;
        RECT 175.810 1313.915 176.090 1314.285 ;
        RECT 1447.250 1313.915 1447.530 1314.285 ;
        RECT 175.880 18.350 176.020 1313.915 ;
        RECT 109.580 18.030 109.840 18.350 ;
        RECT 175.820 18.030 176.080 18.350 ;
        RECT 109.640 2.400 109.780 18.030 ;
        RECT 109.430 -4.800 109.990 2.400 ;
      LAYER via2 ;
        RECT 175.810 1313.960 176.090 1314.240 ;
        RECT 1447.250 1313.960 1447.530 1314.240 ;
      LAYER met3 ;
        RECT 175.785 1314.250 176.115 1314.265 ;
        RECT 1447.225 1314.250 1447.555 1314.265 ;
        RECT 175.785 1313.950 1447.555 1314.250 ;
        RECT 175.785 1313.935 176.115 1313.950 ;
        RECT 1447.225 1313.935 1447.555 1313.950 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 158.845 1315.205 159.015 1316.055 ;
        RECT 227.845 1313.845 228.015 1315.375 ;
        RECT 275.685 1313.845 275.855 1315.035 ;
        RECT 276.145 1314.865 276.315 1316.055 ;
        RECT 323.985 1314.865 324.155 1316.055 ;
        RECT 372.745 1313.505 372.915 1315.035 ;
        RECT 420.585 1313.675 420.755 1315.035 ;
        RECT 420.125 1313.505 420.755 1313.675 ;
        RECT 469.345 1312.485 469.515 1315.035 ;
        RECT 517.185 1312.485 517.355 1315.035 ;
        RECT 565.945 1314.865 566.115 1317.755 ;
        RECT 613.785 1314.865 613.955 1317.755 ;
        RECT 662.545 1311.465 662.715 1315.035 ;
        RECT 726.025 1311.465 726.195 1315.035 ;
        RECT 759.145 1312.825 759.315 1315.035 ;
        RECT 806.985 1312.995 807.155 1315.035 ;
        RECT 855.745 1314.865 855.915 1317.415 ;
        RECT 903.585 1314.865 903.755 1317.415 ;
        RECT 931.645 1314.865 931.815 1315.715 ;
        RECT 806.525 1312.825 807.155 1312.995 ;
      LAYER mcon ;
        RECT 565.945 1317.585 566.115 1317.755 ;
        RECT 158.845 1315.885 159.015 1316.055 ;
        RECT 276.145 1315.885 276.315 1316.055 ;
        RECT 227.845 1315.205 228.015 1315.375 ;
        RECT 275.685 1314.865 275.855 1315.035 ;
        RECT 323.985 1315.885 324.155 1316.055 ;
        RECT 372.745 1314.865 372.915 1315.035 ;
        RECT 420.585 1314.865 420.755 1315.035 ;
        RECT 469.345 1314.865 469.515 1315.035 ;
        RECT 517.185 1314.865 517.355 1315.035 ;
        RECT 613.785 1317.585 613.955 1317.755 ;
        RECT 855.745 1317.245 855.915 1317.415 ;
        RECT 662.545 1314.865 662.715 1315.035 ;
        RECT 726.025 1314.865 726.195 1315.035 ;
        RECT 759.145 1314.865 759.315 1315.035 ;
        RECT 806.985 1314.865 807.155 1315.035 ;
        RECT 903.585 1317.245 903.755 1317.415 ;
        RECT 931.645 1315.545 931.815 1315.715 ;
      LAYER met1 ;
        RECT 565.885 1317.740 566.175 1317.785 ;
        RECT 613.725 1317.740 614.015 1317.785 ;
        RECT 565.885 1317.600 614.015 1317.740 ;
        RECT 565.885 1317.555 566.175 1317.600 ;
        RECT 613.725 1317.555 614.015 1317.600 ;
        RECT 855.685 1317.400 855.975 1317.445 ;
        RECT 903.525 1317.400 903.815 1317.445 ;
        RECT 855.685 1317.260 903.815 1317.400 ;
        RECT 855.685 1317.215 855.975 1317.260 ;
        RECT 903.525 1317.215 903.815 1317.260 ;
        RECT 137.610 1316.040 137.930 1316.100 ;
        RECT 158.785 1316.040 159.075 1316.085 ;
        RECT 137.610 1315.900 159.075 1316.040 ;
        RECT 137.610 1315.840 137.930 1315.900 ;
        RECT 158.785 1315.855 159.075 1315.900 ;
        RECT 276.085 1316.040 276.375 1316.085 ;
        RECT 323.925 1316.040 324.215 1316.085 ;
        RECT 276.085 1315.900 324.215 1316.040 ;
        RECT 276.085 1315.855 276.375 1315.900 ;
        RECT 323.925 1315.855 324.215 1315.900 ;
        RECT 931.585 1315.700 931.875 1315.745 ;
        RECT 1012.990 1315.700 1013.310 1315.760 ;
        RECT 931.585 1315.560 1013.310 1315.700 ;
        RECT 931.585 1315.515 931.875 1315.560 ;
        RECT 1012.990 1315.500 1013.310 1315.560 ;
        RECT 158.785 1315.360 159.075 1315.405 ;
        RECT 227.785 1315.360 228.075 1315.405 ;
        RECT 158.785 1315.220 228.075 1315.360 ;
        RECT 158.785 1315.175 159.075 1315.220 ;
        RECT 227.785 1315.175 228.075 1315.220 ;
        RECT 275.625 1315.020 275.915 1315.065 ;
        RECT 276.085 1315.020 276.375 1315.065 ;
        RECT 275.625 1314.880 276.375 1315.020 ;
        RECT 275.625 1314.835 275.915 1314.880 ;
        RECT 276.085 1314.835 276.375 1314.880 ;
        RECT 323.925 1315.020 324.215 1315.065 ;
        RECT 372.685 1315.020 372.975 1315.065 ;
        RECT 323.925 1314.880 372.975 1315.020 ;
        RECT 323.925 1314.835 324.215 1314.880 ;
        RECT 372.685 1314.835 372.975 1314.880 ;
        RECT 420.525 1315.020 420.815 1315.065 ;
        RECT 469.285 1315.020 469.575 1315.065 ;
        RECT 420.525 1314.880 469.575 1315.020 ;
        RECT 420.525 1314.835 420.815 1314.880 ;
        RECT 469.285 1314.835 469.575 1314.880 ;
        RECT 517.125 1315.020 517.415 1315.065 ;
        RECT 565.885 1315.020 566.175 1315.065 ;
        RECT 517.125 1314.880 566.175 1315.020 ;
        RECT 517.125 1314.835 517.415 1314.880 ;
        RECT 565.885 1314.835 566.175 1314.880 ;
        RECT 613.725 1315.020 614.015 1315.065 ;
        RECT 662.485 1315.020 662.775 1315.065 ;
        RECT 613.725 1314.880 662.775 1315.020 ;
        RECT 613.725 1314.835 614.015 1314.880 ;
        RECT 662.485 1314.835 662.775 1314.880 ;
        RECT 725.965 1315.020 726.255 1315.065 ;
        RECT 759.085 1315.020 759.375 1315.065 ;
        RECT 725.965 1314.880 759.375 1315.020 ;
        RECT 725.965 1314.835 726.255 1314.880 ;
        RECT 759.085 1314.835 759.375 1314.880 ;
        RECT 806.925 1315.020 807.215 1315.065 ;
        RECT 855.685 1315.020 855.975 1315.065 ;
        RECT 806.925 1314.880 855.975 1315.020 ;
        RECT 806.925 1314.835 807.215 1314.880 ;
        RECT 855.685 1314.835 855.975 1314.880 ;
        RECT 903.525 1315.020 903.815 1315.065 ;
        RECT 931.585 1315.020 931.875 1315.065 ;
        RECT 903.525 1314.880 931.875 1315.020 ;
        RECT 903.525 1314.835 903.815 1314.880 ;
        RECT 931.585 1314.835 931.875 1314.880 ;
        RECT 227.785 1314.000 228.075 1314.045 ;
        RECT 275.625 1314.000 275.915 1314.045 ;
        RECT 227.785 1313.860 275.915 1314.000 ;
        RECT 227.785 1313.815 228.075 1313.860 ;
        RECT 275.625 1313.815 275.915 1313.860 ;
        RECT 372.685 1313.660 372.975 1313.705 ;
        RECT 420.065 1313.660 420.355 1313.705 ;
        RECT 372.685 1313.520 420.355 1313.660 ;
        RECT 372.685 1313.475 372.975 1313.520 ;
        RECT 420.065 1313.475 420.355 1313.520 ;
        RECT 759.085 1312.980 759.375 1313.025 ;
        RECT 806.465 1312.980 806.755 1313.025 ;
        RECT 759.085 1312.840 806.755 1312.980 ;
        RECT 759.085 1312.795 759.375 1312.840 ;
        RECT 806.465 1312.795 806.755 1312.840 ;
        RECT 469.285 1312.640 469.575 1312.685 ;
        RECT 517.125 1312.640 517.415 1312.685 ;
        RECT 469.285 1312.500 517.415 1312.640 ;
        RECT 469.285 1312.455 469.575 1312.500 ;
        RECT 517.125 1312.455 517.415 1312.500 ;
        RECT 662.485 1311.620 662.775 1311.665 ;
        RECT 725.965 1311.620 726.255 1311.665 ;
        RECT 662.485 1311.480 726.255 1311.620 ;
        RECT 662.485 1311.435 662.775 1311.480 ;
        RECT 725.965 1311.435 726.255 1311.480 ;
        RECT 133.470 17.240 133.790 17.300 ;
        RECT 137.610 17.240 137.930 17.300 ;
        RECT 133.470 17.100 137.930 17.240 ;
        RECT 133.470 17.040 133.790 17.100 ;
        RECT 137.610 17.040 137.930 17.100 ;
      LAYER via ;
        RECT 137.640 1315.840 137.900 1316.100 ;
        RECT 1013.020 1315.500 1013.280 1315.760 ;
        RECT 133.500 17.040 133.760 17.300 ;
        RECT 137.640 17.040 137.900 17.300 ;
      LAYER met2 ;
        RECT 1013.060 1323.135 1013.340 1327.135 ;
        RECT 137.640 1315.810 137.900 1316.130 ;
        RECT 137.700 17.330 137.840 1315.810 ;
        RECT 1013.080 1315.790 1013.220 1323.135 ;
        RECT 1013.020 1315.470 1013.280 1315.790 ;
        RECT 133.500 17.010 133.760 17.330 ;
        RECT 137.640 17.010 137.900 17.330 ;
        RECT 133.560 2.400 133.700 17.010 ;
        RECT 133.350 -4.800 133.910 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 151.410 1338.820 151.730 1338.880 ;
        RECT 706.630 1338.820 706.950 1338.880 ;
        RECT 151.410 1338.680 706.950 1338.820 ;
        RECT 151.410 1338.620 151.730 1338.680 ;
        RECT 706.630 1338.620 706.950 1338.680 ;
      LAYER via ;
        RECT 151.440 1338.620 151.700 1338.880 ;
        RECT 706.660 1338.620 706.920 1338.880 ;
      LAYER met2 ;
        RECT 706.650 1343.835 706.930 1344.205 ;
        RECT 706.720 1338.910 706.860 1343.835 ;
        RECT 151.440 1338.590 151.700 1338.910 ;
        RECT 706.660 1338.590 706.920 1338.910 ;
        RECT 151.500 2.400 151.640 1338.590 ;
        RECT 151.290 -4.800 151.850 2.400 ;
      LAYER via2 ;
        RECT 706.650 1343.880 706.930 1344.160 ;
      LAYER met3 ;
        RECT 706.625 1344.170 706.955 1344.185 ;
        RECT 715.810 1344.170 719.810 1344.175 ;
        RECT 706.625 1343.870 719.810 1344.170 ;
        RECT 706.625 1343.855 706.955 1343.870 ;
        RECT 715.810 1343.575 719.810 1343.870 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 172.110 1314.680 172.430 1314.740 ;
        RECT 1082.910 1314.680 1083.230 1314.740 ;
        RECT 172.110 1314.540 1083.230 1314.680 ;
        RECT 172.110 1314.480 172.430 1314.540 ;
        RECT 1082.910 1314.480 1083.230 1314.540 ;
        RECT 169.350 17.240 169.670 17.300 ;
        RECT 172.110 17.240 172.430 17.300 ;
        RECT 169.350 17.100 172.430 17.240 ;
        RECT 169.350 17.040 169.670 17.100 ;
        RECT 172.110 17.040 172.430 17.100 ;
      LAYER via ;
        RECT 172.140 1314.480 172.400 1314.740 ;
        RECT 1082.940 1314.480 1083.200 1314.740 ;
        RECT 169.380 17.040 169.640 17.300 ;
        RECT 172.140 17.040 172.400 17.300 ;
      LAYER met2 ;
        RECT 1082.980 1323.135 1083.260 1327.135 ;
        RECT 1083.000 1314.770 1083.140 1323.135 ;
        RECT 172.140 1314.450 172.400 1314.770 ;
        RECT 1082.940 1314.450 1083.200 1314.770 ;
        RECT 172.200 17.330 172.340 1314.450 ;
        RECT 169.380 17.010 169.640 17.330 ;
        RECT 172.140 17.010 172.400 17.330 ;
        RECT 169.440 2.400 169.580 17.010 ;
        RECT 169.230 -4.800 169.790 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 186.830 17.240 187.150 17.300 ;
        RECT 203.390 17.240 203.710 17.300 ;
        RECT 186.830 17.100 203.710 17.240 ;
        RECT 186.830 17.040 187.150 17.100 ;
        RECT 203.390 17.040 203.710 17.100 ;
      LAYER via ;
        RECT 186.860 17.040 187.120 17.300 ;
        RECT 203.420 17.040 203.680 17.300 ;
      LAYER met2 ;
        RECT 203.410 2388.995 203.690 2389.365 ;
        RECT 1253.130 2388.995 1253.410 2389.365 ;
        RECT 203.480 17.330 203.620 2388.995 ;
        RECT 1253.200 2377.880 1253.340 2388.995 ;
        RECT 1253.180 2373.880 1253.460 2377.880 ;
        RECT 186.860 17.010 187.120 17.330 ;
        RECT 203.420 17.010 203.680 17.330 ;
        RECT 186.920 2.400 187.060 17.010 ;
        RECT 186.710 -4.800 187.270 2.400 ;
      LAYER via2 ;
        RECT 203.410 2389.040 203.690 2389.320 ;
        RECT 1253.130 2389.040 1253.410 2389.320 ;
      LAYER met3 ;
        RECT 203.385 2389.330 203.715 2389.345 ;
        RECT 1253.105 2389.330 1253.435 2389.345 ;
        RECT 203.385 2389.030 1253.435 2389.330 ;
        RECT 203.385 2389.015 203.715 2389.030 ;
        RECT 1253.105 2389.015 1253.435 2389.030 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1546.130 1306.860 1546.450 1306.920 ;
        RECT 1549.350 1306.860 1549.670 1306.920 ;
        RECT 1546.130 1306.720 1549.670 1306.860 ;
        RECT 1546.130 1306.660 1546.450 1306.720 ;
        RECT 1549.350 1306.660 1549.670 1306.720 ;
        RECT 204.770 38.660 205.090 38.720 ;
        RECT 1546.130 38.660 1546.450 38.720 ;
        RECT 204.770 38.520 1546.450 38.660 ;
        RECT 204.770 38.460 205.090 38.520 ;
        RECT 1546.130 38.460 1546.450 38.520 ;
      LAYER via ;
        RECT 1546.160 1306.660 1546.420 1306.920 ;
        RECT 1549.380 1306.660 1549.640 1306.920 ;
        RECT 204.800 38.460 205.060 38.720 ;
        RECT 1546.160 38.460 1546.420 38.720 ;
      LAYER met2 ;
        RECT 1551.260 1323.690 1551.540 1327.135 ;
        RECT 1549.440 1323.550 1551.540 1323.690 ;
        RECT 1549.440 1306.950 1549.580 1323.550 ;
        RECT 1551.260 1323.135 1551.540 1323.550 ;
        RECT 1546.160 1306.630 1546.420 1306.950 ;
        RECT 1549.380 1306.630 1549.640 1306.950 ;
        RECT 1546.220 38.750 1546.360 1306.630 ;
        RECT 204.800 38.430 205.060 38.750 ;
        RECT 1546.160 38.430 1546.420 38.750 ;
        RECT 204.860 2.400 205.000 38.430 ;
        RECT 204.650 -4.800 205.210 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 222.730 30.755 223.010 31.125 ;
        RECT 222.800 2.400 222.940 30.755 ;
        RECT 222.590 -4.800 223.150 2.400 ;
      LAYER via2 ;
        RECT 222.730 30.800 223.010 31.080 ;
      LAYER met3 ;
        RECT 1755.835 1681.450 1759.835 1681.455 ;
        RECT 1762.070 1681.450 1762.450 1681.460 ;
        RECT 1755.835 1681.150 1762.450 1681.450 ;
        RECT 1755.835 1680.855 1759.835 1681.150 ;
        RECT 1762.070 1681.140 1762.450 1681.150 ;
        RECT 222.705 31.090 223.035 31.105 ;
        RECT 1762.070 31.090 1762.450 31.100 ;
        RECT 222.705 30.790 1762.450 31.090 ;
        RECT 222.705 30.775 223.035 30.790 ;
        RECT 1762.070 30.780 1762.450 30.790 ;
      LAYER via3 ;
        RECT 1762.100 1681.140 1762.420 1681.460 ;
        RECT 1762.100 30.780 1762.420 31.100 ;
      LAYER met4 ;
        RECT 1762.095 1681.135 1762.425 1681.465 ;
        RECT 1762.110 31.105 1762.410 1681.135 ;
        RECT 1762.095 30.775 1762.425 31.105 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 19.850 1428.580 20.170 1428.640 ;
        RECT 712.610 1428.580 712.930 1428.640 ;
        RECT 19.850 1428.440 712.930 1428.580 ;
        RECT 19.850 1428.380 20.170 1428.440 ;
        RECT 712.610 1428.380 712.930 1428.440 ;
      LAYER via ;
        RECT 19.880 1428.380 20.140 1428.640 ;
        RECT 712.640 1428.380 712.900 1428.640 ;
      LAYER met2 ;
        RECT 712.630 1429.515 712.910 1429.885 ;
        RECT 712.700 1428.670 712.840 1429.515 ;
        RECT 19.880 1428.350 20.140 1428.670 ;
        RECT 712.640 1428.350 712.900 1428.670 ;
        RECT 19.940 17.410 20.080 1428.350 ;
        RECT 19.940 17.270 20.540 17.410 ;
        RECT 20.400 2.400 20.540 17.270 ;
        RECT 20.190 -4.800 20.750 2.400 ;
      LAYER via2 ;
        RECT 712.630 1429.560 712.910 1429.840 ;
      LAYER met3 ;
        RECT 712.605 1429.850 712.935 1429.865 ;
        RECT 715.810 1429.850 719.810 1429.855 ;
        RECT 712.605 1429.550 719.810 1429.850 ;
        RECT 712.605 1429.535 712.935 1429.550 ;
        RECT 715.810 1429.255 719.810 1429.550 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 44.230 31.860 44.550 31.920 ;
        RECT 1359.370 31.860 1359.690 31.920 ;
        RECT 44.230 31.720 1359.690 31.860 ;
        RECT 44.230 31.660 44.550 31.720 ;
        RECT 1359.370 31.660 1359.690 31.720 ;
      LAYER via ;
        RECT 44.260 31.660 44.520 31.920 ;
        RECT 1359.400 31.660 1359.660 31.920 ;
      LAYER met2 ;
        RECT 1359.900 1323.690 1360.180 1327.135 ;
        RECT 1359.460 1323.550 1360.180 1323.690 ;
        RECT 1359.460 31.950 1359.600 1323.550 ;
        RECT 1359.900 1323.135 1360.180 1323.550 ;
        RECT 44.260 31.630 44.520 31.950 ;
        RECT 1359.400 31.630 1359.660 31.950 ;
        RECT 44.320 2.400 44.460 31.630 ;
        RECT 44.110 -4.800 44.670 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 266.040 17.100 519.640 17.240 ;
        RECT 246.630 16.900 246.950 16.960 ;
        RECT 266.040 16.900 266.180 17.100 ;
        RECT 246.630 16.760 266.180 16.900 ;
        RECT 246.630 16.700 246.950 16.760 ;
        RECT 519.500 15.880 519.640 17.100 ;
        RECT 562.190 15.880 562.510 15.940 ;
        RECT 519.500 15.740 562.510 15.880 ;
        RECT 562.190 15.680 562.510 15.740 ;
      LAYER via ;
        RECT 246.660 16.700 246.920 16.960 ;
        RECT 562.220 15.680 562.480 15.940 ;
      LAYER met2 ;
        RECT 562.210 2388.315 562.490 2388.685 ;
        RECT 1178.610 2388.315 1178.890 2388.685 ;
        RECT 246.660 16.670 246.920 16.990 ;
        RECT 246.720 2.400 246.860 16.670 ;
        RECT 562.280 15.970 562.420 2388.315 ;
        RECT 1178.680 2377.880 1178.820 2388.315 ;
        RECT 1178.660 2373.880 1178.940 2377.880 ;
        RECT 562.220 15.650 562.480 15.970 ;
        RECT 246.510 -4.800 247.070 2.400 ;
      LAYER via2 ;
        RECT 562.210 2388.360 562.490 2388.640 ;
        RECT 1178.610 2388.360 1178.890 2388.640 ;
      LAYER met3 ;
        RECT 562.185 2388.650 562.515 2388.665 ;
        RECT 1178.585 2388.650 1178.915 2388.665 ;
        RECT 562.185 2388.350 1178.915 2388.650 ;
        RECT 562.185 2388.335 562.515 2388.350 ;
        RECT 1178.585 2388.335 1178.915 2388.350 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 264.110 33.560 264.430 33.620 ;
        RECT 1256.330 33.560 1256.650 33.620 ;
        RECT 264.110 33.420 1256.650 33.560 ;
        RECT 264.110 33.360 264.430 33.420 ;
        RECT 1256.330 33.360 1256.650 33.420 ;
      LAYER via ;
        RECT 264.140 33.360 264.400 33.620 ;
        RECT 1256.360 33.360 1256.620 33.620 ;
      LAYER met2 ;
        RECT 1262.380 1323.690 1262.660 1327.135 ;
        RECT 1256.420 1323.550 1262.660 1323.690 ;
        RECT 1256.420 33.650 1256.560 1323.550 ;
        RECT 1262.380 1323.135 1262.660 1323.550 ;
        RECT 264.140 33.330 264.400 33.650 ;
        RECT 1256.360 33.330 1256.620 33.650 ;
        RECT 264.200 2.400 264.340 33.330 ;
        RECT 263.990 -4.800 264.550 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 282.050 33.220 282.370 33.280 ;
        RECT 1345.570 33.220 1345.890 33.280 ;
        RECT 282.050 33.080 1345.890 33.220 ;
        RECT 282.050 33.020 282.370 33.080 ;
        RECT 1345.570 33.020 1345.890 33.080 ;
      LAYER via ;
        RECT 282.080 33.020 282.340 33.280 ;
        RECT 1345.600 33.020 1345.860 33.280 ;
      LAYER met2 ;
        RECT 1348.860 1323.690 1349.140 1327.135 ;
        RECT 1345.660 1323.550 1349.140 1323.690 ;
        RECT 1345.660 33.310 1345.800 1323.550 ;
        RECT 1348.860 1323.135 1349.140 1323.550 ;
        RECT 282.080 32.990 282.340 33.310 ;
        RECT 1345.600 32.990 1345.860 33.310 ;
        RECT 282.140 2.400 282.280 32.990 ;
        RECT 281.930 -4.800 282.490 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 303.210 1314.000 303.530 1314.060 ;
        RECT 886.030 1314.000 886.350 1314.060 ;
        RECT 303.210 1313.860 886.350 1314.000 ;
        RECT 303.210 1313.800 303.530 1313.860 ;
        RECT 886.030 1313.800 886.350 1313.860 ;
        RECT 299.990 14.520 300.310 14.580 ;
        RECT 303.210 14.520 303.530 14.580 ;
        RECT 299.990 14.380 303.530 14.520 ;
        RECT 299.990 14.320 300.310 14.380 ;
        RECT 303.210 14.320 303.530 14.380 ;
      LAYER via ;
        RECT 303.240 1313.800 303.500 1314.060 ;
        RECT 886.060 1313.800 886.320 1314.060 ;
        RECT 300.020 14.320 300.280 14.580 ;
        RECT 303.240 14.320 303.500 14.580 ;
      LAYER met2 ;
        RECT 886.100 1323.135 886.380 1327.135 ;
        RECT 886.120 1314.090 886.260 1323.135 ;
        RECT 303.240 1313.770 303.500 1314.090 ;
        RECT 886.060 1313.770 886.320 1314.090 ;
        RECT 303.300 14.610 303.440 1313.770 ;
        RECT 300.020 14.290 300.280 14.610 ;
        RECT 303.240 14.290 303.500 14.610 ;
        RECT 300.080 2.400 300.220 14.290 ;
        RECT 299.870 -4.800 300.430 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 323.450 1566.620 323.770 1566.680 ;
        RECT 710.310 1566.620 710.630 1566.680 ;
        RECT 323.450 1566.480 710.630 1566.620 ;
        RECT 323.450 1566.420 323.770 1566.480 ;
        RECT 710.310 1566.420 710.630 1566.480 ;
        RECT 317.930 16.900 318.250 16.960 ;
        RECT 323.450 16.900 323.770 16.960 ;
        RECT 317.930 16.760 323.770 16.900 ;
        RECT 317.930 16.700 318.250 16.760 ;
        RECT 323.450 16.700 323.770 16.760 ;
      LAYER via ;
        RECT 323.480 1566.420 323.740 1566.680 ;
        RECT 710.340 1566.420 710.600 1566.680 ;
        RECT 317.960 16.700 318.220 16.960 ;
        RECT 323.480 16.700 323.740 16.960 ;
      LAYER met2 ;
        RECT 710.330 1566.875 710.610 1567.245 ;
        RECT 710.400 1566.710 710.540 1566.875 ;
        RECT 323.480 1566.390 323.740 1566.710 ;
        RECT 710.340 1566.390 710.600 1566.710 ;
        RECT 323.540 16.990 323.680 1566.390 ;
        RECT 317.960 16.670 318.220 16.990 ;
        RECT 323.480 16.670 323.740 16.990 ;
        RECT 318.020 2.400 318.160 16.670 ;
        RECT 317.810 -4.800 318.370 2.400 ;
      LAYER via2 ;
        RECT 710.330 1566.920 710.610 1567.200 ;
      LAYER met3 ;
        RECT 710.305 1567.210 710.635 1567.225 ;
        RECT 715.810 1567.210 719.810 1567.215 ;
        RECT 710.305 1566.910 719.810 1567.210 ;
        RECT 710.305 1566.895 710.635 1566.910 ;
        RECT 715.810 1566.615 719.810 1566.910 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 335.870 32.200 336.190 32.260 ;
        RECT 1476.670 32.200 1476.990 32.260 ;
        RECT 335.870 32.060 1476.990 32.200 ;
        RECT 335.870 32.000 336.190 32.060 ;
        RECT 1476.670 32.000 1476.990 32.060 ;
      LAYER via ;
        RECT 335.900 32.000 336.160 32.260 ;
        RECT 1476.700 32.000 1476.960 32.260 ;
      LAYER met2 ;
        RECT 1482.260 1323.690 1482.540 1327.135 ;
        RECT 1476.760 1323.550 1482.540 1323.690 ;
        RECT 1476.760 32.290 1476.900 1323.550 ;
        RECT 1482.260 1323.135 1482.540 1323.550 ;
        RECT 335.900 31.970 336.160 32.290 ;
        RECT 1476.700 31.970 1476.960 32.290 ;
        RECT 335.960 2.400 336.100 31.970 ;
        RECT 335.750 -4.800 336.310 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 362.090 2389.760 362.410 2389.820 ;
        RECT 871.310 2389.760 871.630 2389.820 ;
        RECT 362.090 2389.620 871.630 2389.760 ;
        RECT 362.090 2389.560 362.410 2389.620 ;
        RECT 871.310 2389.560 871.630 2389.620 ;
        RECT 353.350 16.900 353.670 16.960 ;
        RECT 362.090 16.900 362.410 16.960 ;
        RECT 353.350 16.760 362.410 16.900 ;
        RECT 353.350 16.700 353.670 16.760 ;
        RECT 362.090 16.700 362.410 16.760 ;
      LAYER via ;
        RECT 362.120 2389.560 362.380 2389.820 ;
        RECT 871.340 2389.560 871.600 2389.820 ;
        RECT 353.380 16.700 353.640 16.960 ;
        RECT 362.120 16.700 362.380 16.960 ;
      LAYER met2 ;
        RECT 362.120 2389.530 362.380 2389.850 ;
        RECT 871.340 2389.530 871.600 2389.850 ;
        RECT 362.180 16.990 362.320 2389.530 ;
        RECT 871.400 2377.880 871.540 2389.530 ;
        RECT 871.380 2373.880 871.660 2377.880 ;
        RECT 353.380 16.670 353.640 16.990 ;
        RECT 362.120 16.670 362.380 16.990 ;
        RECT 353.440 2.400 353.580 16.670 ;
        RECT 353.230 -4.800 353.790 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 372.210 1316.720 372.530 1316.780 ;
        RECT 1174.910 1316.720 1175.230 1316.780 ;
        RECT 372.210 1316.580 1175.230 1316.720 ;
        RECT 372.210 1316.520 372.530 1316.580 ;
        RECT 1174.910 1316.520 1175.230 1316.580 ;
      LAYER via ;
        RECT 372.240 1316.520 372.500 1316.780 ;
        RECT 1174.940 1316.520 1175.200 1316.780 ;
      LAYER met2 ;
        RECT 1174.980 1323.135 1175.260 1327.135 ;
        RECT 1175.000 1316.810 1175.140 1323.135 ;
        RECT 372.240 1316.490 372.500 1316.810 ;
        RECT 1174.940 1316.490 1175.200 1316.810 ;
        RECT 372.300 16.900 372.440 1316.490 ;
        RECT 371.380 16.760 372.440 16.900 ;
        RECT 371.380 2.400 371.520 16.760 ;
        RECT 371.170 -4.800 371.730 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 392.910 1877.040 393.230 1877.100 ;
        RECT 704.330 1877.040 704.650 1877.100 ;
        RECT 392.910 1876.900 704.650 1877.040 ;
        RECT 392.910 1876.840 393.230 1876.900 ;
        RECT 704.330 1876.840 704.650 1876.900 ;
        RECT 389.230 16.900 389.550 16.960 ;
        RECT 392.910 16.900 393.230 16.960 ;
        RECT 389.230 16.760 393.230 16.900 ;
        RECT 389.230 16.700 389.550 16.760 ;
        RECT 392.910 16.700 393.230 16.760 ;
      LAYER via ;
        RECT 392.940 1876.840 393.200 1877.100 ;
        RECT 704.360 1876.840 704.620 1877.100 ;
        RECT 389.260 16.700 389.520 16.960 ;
        RECT 392.940 16.700 393.200 16.960 ;
      LAYER met2 ;
        RECT 704.350 1882.395 704.630 1882.765 ;
        RECT 704.420 1877.130 704.560 1882.395 ;
        RECT 392.940 1876.810 393.200 1877.130 ;
        RECT 704.360 1876.810 704.620 1877.130 ;
        RECT 393.000 16.990 393.140 1876.810 ;
        RECT 389.260 16.670 389.520 16.990 ;
        RECT 392.940 16.670 393.200 16.990 ;
        RECT 389.320 2.400 389.460 16.670 ;
        RECT 389.110 -4.800 389.670 2.400 ;
      LAYER via2 ;
        RECT 704.350 1882.440 704.630 1882.720 ;
      LAYER met3 ;
        RECT 704.325 1882.730 704.655 1882.745 ;
        RECT 715.810 1882.730 719.810 1882.735 ;
        RECT 704.325 1882.430 719.810 1882.730 ;
        RECT 704.325 1882.415 704.655 1882.430 ;
        RECT 715.810 1882.135 719.810 1882.430 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 407.170 19.960 407.490 20.020 ;
        RECT 444.890 19.960 445.210 20.020 ;
        RECT 407.170 19.820 445.210 19.960 ;
        RECT 407.170 19.760 407.490 19.820 ;
        RECT 444.890 19.760 445.210 19.820 ;
      LAYER via ;
        RECT 407.200 19.760 407.460 20.020 ;
        RECT 444.920 19.760 445.180 20.020 ;
      LAYER met2 ;
        RECT 444.910 2389.675 445.190 2390.045 ;
        RECT 1658.850 2389.675 1659.130 2390.045 ;
        RECT 444.980 20.050 445.120 2389.675 ;
        RECT 1658.920 2377.880 1659.060 2389.675 ;
        RECT 1658.900 2373.880 1659.180 2377.880 ;
        RECT 407.200 19.730 407.460 20.050 ;
        RECT 444.920 19.730 445.180 20.050 ;
        RECT 407.260 2.400 407.400 19.730 ;
        RECT 407.050 -4.800 407.610 2.400 ;
      LAYER via2 ;
        RECT 444.910 2389.720 445.190 2390.000 ;
        RECT 1658.850 2389.720 1659.130 2390.000 ;
      LAYER met3 ;
        RECT 444.885 2390.010 445.215 2390.025 ;
        RECT 1658.825 2390.010 1659.155 2390.025 ;
        RECT 444.885 2389.710 1659.155 2390.010 ;
        RECT 444.885 2389.695 445.215 2389.710 ;
        RECT 1658.825 2389.695 1659.155 2389.710 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 68.150 18.600 68.470 18.660 ;
        RECT 106.790 18.600 107.110 18.660 ;
        RECT 68.150 18.460 107.110 18.600 ;
        RECT 68.150 18.400 68.470 18.460 ;
        RECT 106.790 18.400 107.110 18.460 ;
      LAYER via ;
        RECT 68.180 18.400 68.440 18.660 ;
        RECT 106.820 18.400 107.080 18.660 ;
      LAYER met2 ;
        RECT 1267.900 1323.135 1268.180 1327.135 ;
        RECT 1267.920 1314.965 1268.060 1323.135 ;
        RECT 106.810 1314.595 107.090 1314.965 ;
        RECT 1267.850 1314.595 1268.130 1314.965 ;
        RECT 106.880 18.690 107.020 1314.595 ;
        RECT 68.180 18.370 68.440 18.690 ;
        RECT 106.820 18.370 107.080 18.690 ;
        RECT 68.240 2.400 68.380 18.370 ;
        RECT 68.030 -4.800 68.590 2.400 ;
      LAYER via2 ;
        RECT 106.810 1314.640 107.090 1314.920 ;
        RECT 1267.850 1314.640 1268.130 1314.920 ;
      LAYER met3 ;
        RECT 106.785 1314.930 107.115 1314.945 ;
        RECT 1267.825 1314.930 1268.155 1314.945 ;
        RECT 106.785 1314.630 1268.155 1314.930 ;
        RECT 106.785 1314.615 107.115 1314.630 ;
        RECT 1267.825 1314.615 1268.155 1314.630 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1459.190 2387.720 1459.510 2387.780 ;
        RECT 1652.390 2387.720 1652.710 2387.780 ;
        RECT 1459.190 2387.580 1652.710 2387.720 ;
        RECT 1459.190 2387.520 1459.510 2387.580 ;
        RECT 1652.390 2387.520 1652.710 2387.580 ;
        RECT 424.650 16.900 424.970 16.960 ;
        RECT 427.410 16.900 427.730 16.960 ;
        RECT 424.650 16.760 427.730 16.900 ;
        RECT 424.650 16.700 424.970 16.760 ;
        RECT 427.410 16.700 427.730 16.760 ;
      LAYER via ;
        RECT 1459.220 2387.520 1459.480 2387.780 ;
        RECT 1652.420 2387.520 1652.680 2387.780 ;
        RECT 424.680 16.700 424.940 16.960 ;
        RECT 427.440 16.700 427.700 16.960 ;
      LAYER met2 ;
        RECT 1459.220 2387.490 1459.480 2387.810 ;
        RECT 1652.420 2387.490 1652.680 2387.810 ;
        RECT 1459.280 2380.525 1459.420 2387.490 ;
        RECT 1459.210 2380.155 1459.490 2380.525 ;
        RECT 427.430 2379.475 427.710 2379.845 ;
        RECT 427.500 16.990 427.640 2379.475 ;
        RECT 1652.480 2377.880 1652.620 2387.490 ;
        RECT 1652.460 2373.880 1652.740 2377.880 ;
        RECT 424.680 16.670 424.940 16.990 ;
        RECT 427.440 16.670 427.700 16.990 ;
        RECT 424.740 2.400 424.880 16.670 ;
        RECT 424.530 -4.800 425.090 2.400 ;
      LAYER via2 ;
        RECT 1459.210 2380.200 1459.490 2380.480 ;
        RECT 427.430 2379.520 427.710 2379.800 ;
      LAYER met3 ;
        RECT 1459.185 2380.490 1459.515 2380.505 ;
        RECT 1438.270 2380.190 1459.515 2380.490 ;
        RECT 427.405 2379.810 427.735 2379.825 ;
        RECT 1438.270 2379.810 1438.570 2380.190 ;
        RECT 1459.185 2380.175 1459.515 2380.190 ;
        RECT 427.405 2379.510 1438.570 2379.810 ;
        RECT 427.405 2379.495 427.735 2379.510 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1749.010 2374.290 1749.290 2374.405 ;
        RECT 1750.900 2374.290 1751.180 2377.880 ;
        RECT 1749.010 2374.150 1751.180 2374.290 ;
        RECT 1749.010 2374.035 1749.290 2374.150 ;
        RECT 1750.900 2373.880 1751.180 2374.150 ;
        RECT 442.610 45.715 442.890 46.085 ;
        RECT 442.680 2.400 442.820 45.715 ;
        RECT 442.470 -4.800 443.030 2.400 ;
      LAYER via2 ;
        RECT 1749.010 2374.080 1749.290 2374.360 ;
        RECT 442.610 45.760 442.890 46.040 ;
      LAYER met3 ;
        RECT 1746.430 2374.370 1746.810 2374.380 ;
        RECT 1748.985 2374.370 1749.315 2374.385 ;
        RECT 1746.430 2374.070 1749.315 2374.370 ;
        RECT 1746.430 2374.060 1746.810 2374.070 ;
        RECT 1748.985 2374.055 1749.315 2374.070 ;
        RECT 442.585 46.050 442.915 46.065 ;
        RECT 1746.430 46.050 1746.810 46.060 ;
        RECT 442.585 45.750 1746.810 46.050 ;
        RECT 442.585 45.735 442.915 45.750 ;
        RECT 1746.430 45.740 1746.810 45.750 ;
      LAYER via3 ;
        RECT 1746.460 2374.060 1746.780 2374.380 ;
        RECT 1746.460 45.740 1746.780 46.060 ;
      LAYER met4 ;
        RECT 1746.455 2374.055 1746.785 2374.385 ;
        RECT 1746.470 46.065 1746.770 2374.055 ;
        RECT 1746.455 45.735 1746.785 46.065 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 460.530 20.300 460.850 20.360 ;
        RECT 638.090 20.300 638.410 20.360 ;
        RECT 460.530 20.160 638.410 20.300 ;
        RECT 460.530 20.100 460.850 20.160 ;
        RECT 638.090 20.100 638.410 20.160 ;
      LAYER via ;
        RECT 460.560 20.100 460.820 20.360 ;
        RECT 638.120 20.100 638.380 20.360 ;
      LAYER met2 ;
        RECT 638.110 2391.035 638.390 2391.405 ;
        RECT 1531.430 2391.035 1531.710 2391.405 ;
        RECT 638.180 20.390 638.320 2391.035 ;
        RECT 1531.500 2389.250 1531.640 2391.035 ;
        RECT 1531.500 2389.110 1532.560 2389.250 ;
        RECT 1532.420 2377.690 1532.560 2389.110 ;
        RECT 1537.460 2377.690 1537.740 2377.880 ;
        RECT 1532.420 2377.550 1537.740 2377.690 ;
        RECT 1537.460 2373.880 1537.740 2377.550 ;
        RECT 460.560 20.070 460.820 20.390 ;
        RECT 638.120 20.070 638.380 20.390 ;
        RECT 460.620 2.400 460.760 20.070 ;
        RECT 460.410 -4.800 460.970 2.400 ;
      LAYER via2 ;
        RECT 638.110 2391.080 638.390 2391.360 ;
        RECT 1531.430 2391.080 1531.710 2391.360 ;
      LAYER met3 ;
        RECT 638.085 2391.370 638.415 2391.385 ;
        RECT 1531.405 2391.370 1531.735 2391.385 ;
        RECT 638.085 2391.070 1531.735 2391.370 ;
        RECT 638.085 2391.055 638.415 2391.070 ;
        RECT 1531.405 2391.055 1531.735 2391.070 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 482.610 1313.320 482.930 1313.380 ;
        RECT 1088.430 1313.320 1088.750 1313.380 ;
        RECT 482.610 1313.180 1088.750 1313.320 ;
        RECT 482.610 1313.120 482.930 1313.180 ;
        RECT 1088.430 1313.120 1088.750 1313.180 ;
        RECT 478.470 16.900 478.790 16.960 ;
        RECT 482.610 16.900 482.930 16.960 ;
        RECT 478.470 16.760 482.930 16.900 ;
        RECT 478.470 16.700 478.790 16.760 ;
        RECT 482.610 16.700 482.930 16.760 ;
      LAYER via ;
        RECT 482.640 1313.120 482.900 1313.380 ;
        RECT 1088.460 1313.120 1088.720 1313.380 ;
        RECT 478.500 16.700 478.760 16.960 ;
        RECT 482.640 16.700 482.900 16.960 ;
      LAYER met2 ;
        RECT 1088.500 1323.135 1088.780 1327.135 ;
        RECT 1088.520 1313.410 1088.660 1323.135 ;
        RECT 482.640 1313.090 482.900 1313.410 ;
        RECT 1088.460 1313.090 1088.720 1313.410 ;
        RECT 482.700 16.990 482.840 1313.090 ;
        RECT 478.500 16.670 478.760 16.990 ;
        RECT 482.640 16.670 482.900 16.990 ;
        RECT 478.560 2.400 478.700 16.670 ;
        RECT 478.350 -4.800 478.910 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 686.390 2387.720 686.710 2387.780 ;
        RECT 848.310 2387.720 848.630 2387.780 ;
        RECT 686.390 2387.580 848.630 2387.720 ;
        RECT 686.390 2387.520 686.710 2387.580 ;
        RECT 848.310 2387.520 848.630 2387.580 ;
        RECT 495.950 19.960 496.270 20.020 ;
        RECT 686.390 19.960 686.710 20.020 ;
        RECT 495.950 19.820 686.710 19.960 ;
        RECT 495.950 19.760 496.270 19.820 ;
        RECT 686.390 19.760 686.710 19.820 ;
      LAYER via ;
        RECT 686.420 2387.520 686.680 2387.780 ;
        RECT 848.340 2387.520 848.600 2387.780 ;
        RECT 495.980 19.760 496.240 20.020 ;
        RECT 686.420 19.760 686.680 20.020 ;
      LAYER met2 ;
        RECT 686.420 2387.490 686.680 2387.810 ;
        RECT 848.340 2387.490 848.600 2387.810 ;
        RECT 686.480 20.050 686.620 2387.490 ;
        RECT 848.400 2377.880 848.540 2387.490 ;
        RECT 848.380 2373.880 848.660 2377.880 ;
        RECT 495.980 19.730 496.240 20.050 ;
        RECT 686.420 19.730 686.680 20.050 ;
        RECT 496.040 9.930 496.180 19.730 ;
        RECT 496.040 9.790 496.640 9.930 ;
        RECT 496.500 2.400 496.640 9.790 ;
        RECT 496.290 -4.800 496.850 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 517.110 2173.860 517.430 2173.920 ;
        RECT 709.390 2173.860 709.710 2173.920 ;
        RECT 517.110 2173.720 709.710 2173.860 ;
        RECT 517.110 2173.660 517.430 2173.720 ;
        RECT 709.390 2173.660 709.710 2173.720 ;
        RECT 513.890 16.900 514.210 16.960 ;
        RECT 517.110 16.900 517.430 16.960 ;
        RECT 513.890 16.760 517.430 16.900 ;
        RECT 513.890 16.700 514.210 16.760 ;
        RECT 517.110 16.700 517.430 16.760 ;
      LAYER via ;
        RECT 517.140 2173.660 517.400 2173.920 ;
        RECT 709.420 2173.660 709.680 2173.920 ;
        RECT 513.920 16.700 514.180 16.960 ;
        RECT 517.140 16.700 517.400 16.960 ;
      LAYER met2 ;
        RECT 517.140 2173.630 517.400 2173.950 ;
        RECT 709.420 2173.805 709.680 2173.950 ;
        RECT 517.200 16.990 517.340 2173.630 ;
        RECT 709.410 2173.435 709.690 2173.805 ;
        RECT 513.920 16.670 514.180 16.990 ;
        RECT 517.140 16.670 517.400 16.990 ;
        RECT 513.980 2.400 514.120 16.670 ;
        RECT 513.770 -4.800 514.330 2.400 ;
      LAYER via2 ;
        RECT 709.410 2173.480 709.690 2173.760 ;
      LAYER met3 ;
        RECT 709.385 2173.770 709.715 2173.785 ;
        RECT 715.810 2173.770 719.810 2173.775 ;
        RECT 709.385 2173.470 719.810 2173.770 ;
        RECT 709.385 2173.455 709.715 2173.470 ;
        RECT 715.810 2173.175 719.810 2173.470 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 693.290 2391.460 693.610 2391.520 ;
        RECT 1293.590 2391.460 1293.910 2391.520 ;
        RECT 693.290 2391.320 1293.910 2391.460 ;
        RECT 693.290 2391.260 693.610 2391.320 ;
        RECT 1293.590 2391.260 1293.910 2391.320 ;
        RECT 531.830 20.640 532.150 20.700 ;
        RECT 693.290 20.640 693.610 20.700 ;
        RECT 531.830 20.500 693.610 20.640 ;
        RECT 531.830 20.440 532.150 20.500 ;
        RECT 693.290 20.440 693.610 20.500 ;
      LAYER via ;
        RECT 693.320 2391.260 693.580 2391.520 ;
        RECT 1293.620 2391.260 1293.880 2391.520 ;
        RECT 531.860 20.440 532.120 20.700 ;
        RECT 693.320 20.440 693.580 20.700 ;
      LAYER met2 ;
        RECT 693.320 2391.230 693.580 2391.550 ;
        RECT 1293.620 2391.230 1293.880 2391.550 ;
        RECT 693.380 20.730 693.520 2391.230 ;
        RECT 1293.680 2377.880 1293.820 2391.230 ;
        RECT 1293.660 2373.880 1293.940 2377.880 ;
        RECT 531.860 20.410 532.120 20.730 ;
        RECT 693.320 20.410 693.580 20.730 ;
        RECT 531.920 2.400 532.060 20.410 ;
        RECT 531.710 -4.800 532.270 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 549.790 38.235 550.070 38.605 ;
        RECT 549.860 2.400 550.000 38.235 ;
        RECT 549.650 -4.800 550.210 2.400 ;
      LAYER via2 ;
        RECT 549.790 38.280 550.070 38.560 ;
      LAYER met3 ;
        RECT 1755.835 1980.650 1759.835 1980.655 ;
        RECT 1761.150 1980.650 1761.530 1980.660 ;
        RECT 1755.835 1980.350 1761.530 1980.650 ;
        RECT 1755.835 1980.055 1759.835 1980.350 ;
        RECT 1761.150 1980.340 1761.530 1980.350 ;
        RECT 549.765 38.570 550.095 38.585 ;
        RECT 1761.150 38.570 1761.530 38.580 ;
        RECT 549.765 38.270 1761.530 38.570 ;
        RECT 549.765 38.255 550.095 38.270 ;
        RECT 1761.150 38.260 1761.530 38.270 ;
      LAYER via3 ;
        RECT 1761.180 1980.340 1761.500 1980.660 ;
        RECT 1761.180 38.260 1761.500 38.580 ;
      LAYER met4 ;
        RECT 1761.175 1980.335 1761.505 1980.665 ;
        RECT 1761.190 38.585 1761.490 1980.335 ;
        RECT 1761.175 38.255 1761.505 38.585 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 572.310 80.140 572.630 80.200 ;
        RECT 1760.950 80.140 1761.270 80.200 ;
        RECT 572.310 80.000 1761.270 80.140 ;
        RECT 572.310 79.940 572.630 80.000 ;
        RECT 1760.950 79.940 1761.270 80.000 ;
        RECT 567.710 15.540 568.030 15.600 ;
        RECT 572.310 15.540 572.630 15.600 ;
        RECT 567.710 15.400 572.630 15.540 ;
        RECT 567.710 15.340 568.030 15.400 ;
        RECT 572.310 15.340 572.630 15.400 ;
      LAYER via ;
        RECT 572.340 79.940 572.600 80.200 ;
        RECT 1760.980 79.940 1761.240 80.200 ;
        RECT 567.740 15.340 568.000 15.600 ;
        RECT 572.340 15.340 572.600 15.600 ;
      LAYER met2 ;
        RECT 1760.970 1997.995 1761.250 1998.365 ;
        RECT 1761.040 80.230 1761.180 1997.995 ;
        RECT 572.340 79.910 572.600 80.230 ;
        RECT 1760.980 79.910 1761.240 80.230 ;
        RECT 572.400 15.630 572.540 79.910 ;
        RECT 567.740 15.310 568.000 15.630 ;
        RECT 572.340 15.310 572.600 15.630 ;
        RECT 567.800 2.400 567.940 15.310 ;
        RECT 567.590 -4.800 568.150 2.400 ;
      LAYER via2 ;
        RECT 1760.970 1998.040 1761.250 1998.320 ;
      LAYER met3 ;
        RECT 1755.835 1998.330 1759.835 1998.335 ;
        RECT 1760.945 1998.330 1761.275 1998.345 ;
        RECT 1755.835 1998.030 1761.275 1998.330 ;
        RECT 1755.835 1997.735 1759.835 1998.030 ;
        RECT 1760.945 1998.015 1761.275 1998.030 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 783.065 2389.265 784.155 2389.435 ;
        RECT 783.985 2388.925 784.155 2389.265 ;
      LAYER met1 ;
        RECT 586.110 2389.420 586.430 2389.480 ;
        RECT 783.005 2389.420 783.295 2389.465 ;
        RECT 586.110 2389.280 783.295 2389.420 ;
        RECT 586.110 2389.220 586.430 2389.280 ;
        RECT 783.005 2389.235 783.295 2389.280 ;
        RECT 783.925 2389.080 784.215 2389.125 ;
        RECT 819.790 2389.080 820.110 2389.140 ;
        RECT 783.925 2388.940 820.110 2389.080 ;
        RECT 783.925 2388.895 784.215 2388.940 ;
        RECT 819.790 2388.880 820.110 2388.940 ;
      LAYER via ;
        RECT 586.140 2389.220 586.400 2389.480 ;
        RECT 819.820 2388.880 820.080 2389.140 ;
      LAYER met2 ;
        RECT 586.140 2389.190 586.400 2389.510 ;
        RECT 586.200 17.410 586.340 2389.190 ;
        RECT 819.820 2388.850 820.080 2389.170 ;
        RECT 819.880 2377.880 820.020 2388.850 ;
        RECT 819.860 2373.880 820.140 2377.880 ;
        RECT 585.740 17.270 586.340 17.410 ;
        RECT 585.740 2.400 585.880 17.270 ;
        RECT 585.530 -4.800 586.090 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 96.210 1314.340 96.530 1314.400 ;
        RECT 1024.950 1314.340 1025.270 1314.400 ;
        RECT 96.210 1314.200 1025.270 1314.340 ;
        RECT 96.210 1314.140 96.530 1314.200 ;
        RECT 1024.950 1314.140 1025.270 1314.200 ;
        RECT 91.610 17.920 91.930 17.980 ;
        RECT 96.210 17.920 96.530 17.980 ;
        RECT 91.610 17.780 96.530 17.920 ;
        RECT 91.610 17.720 91.930 17.780 ;
        RECT 96.210 17.720 96.530 17.780 ;
      LAYER via ;
        RECT 96.240 1314.140 96.500 1314.400 ;
        RECT 1024.980 1314.140 1025.240 1314.400 ;
        RECT 91.640 17.720 91.900 17.980 ;
        RECT 96.240 17.720 96.500 17.980 ;
      LAYER met2 ;
        RECT 1025.020 1323.135 1025.300 1327.135 ;
        RECT 1025.040 1314.430 1025.180 1323.135 ;
        RECT 96.240 1314.110 96.500 1314.430 ;
        RECT 1024.980 1314.110 1025.240 1314.430 ;
        RECT 96.300 18.010 96.440 1314.110 ;
        RECT 91.640 17.690 91.900 18.010 ;
        RECT 96.240 17.690 96.500 18.010 ;
        RECT 91.700 2.400 91.840 17.690 ;
        RECT 91.490 -4.800 92.050 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 606.810 80.480 607.130 80.540 ;
        RECT 1766.010 80.480 1766.330 80.540 ;
        RECT 606.810 80.340 1766.330 80.480 ;
        RECT 606.810 80.280 607.130 80.340 ;
        RECT 1766.010 80.280 1766.330 80.340 ;
        RECT 603.130 17.240 603.450 17.300 ;
        RECT 606.810 17.240 607.130 17.300 ;
        RECT 603.130 17.100 607.130 17.240 ;
        RECT 603.130 17.040 603.450 17.100 ;
        RECT 606.810 17.040 607.130 17.100 ;
      LAYER via ;
        RECT 606.840 80.280 607.100 80.540 ;
        RECT 1766.040 80.280 1766.300 80.540 ;
        RECT 603.160 17.040 603.420 17.300 ;
        RECT 606.840 17.040 607.100 17.300 ;
      LAYER met2 ;
        RECT 1766.030 1405.035 1766.310 1405.405 ;
        RECT 1766.100 80.570 1766.240 1405.035 ;
        RECT 606.840 80.250 607.100 80.570 ;
        RECT 1766.040 80.250 1766.300 80.570 ;
        RECT 606.900 17.330 607.040 80.250 ;
        RECT 603.160 17.010 603.420 17.330 ;
        RECT 606.840 17.010 607.100 17.330 ;
        RECT 603.220 2.400 603.360 17.010 ;
        RECT 603.010 -4.800 603.570 2.400 ;
      LAYER via2 ;
        RECT 1766.030 1405.080 1766.310 1405.360 ;
      LAYER met3 ;
        RECT 1755.835 1407.495 1759.835 1408.095 ;
        RECT 1759.350 1405.370 1759.650 1407.495 ;
        RECT 1766.005 1405.370 1766.335 1405.385 ;
        RECT 1759.350 1405.070 1766.335 1405.370 ;
        RECT 1766.005 1405.055 1766.335 1405.070 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 627.050 886.960 627.370 887.020 ;
        RECT 1771.530 886.960 1771.850 887.020 ;
        RECT 627.050 886.820 1771.850 886.960 ;
        RECT 627.050 886.760 627.370 886.820 ;
        RECT 1771.530 886.760 1771.850 886.820 ;
        RECT 621.070 18.260 621.390 18.320 ;
        RECT 627.050 18.260 627.370 18.320 ;
        RECT 621.070 18.120 627.370 18.260 ;
        RECT 621.070 18.060 621.390 18.120 ;
        RECT 627.050 18.060 627.370 18.120 ;
      LAYER via ;
        RECT 627.080 886.760 627.340 887.020 ;
        RECT 1771.560 886.760 1771.820 887.020 ;
        RECT 621.100 18.060 621.360 18.320 ;
        RECT 627.080 18.060 627.340 18.320 ;
      LAYER met2 ;
        RECT 1771.550 1449.915 1771.830 1450.285 ;
        RECT 1771.620 887.050 1771.760 1449.915 ;
        RECT 627.080 886.730 627.340 887.050 ;
        RECT 1771.560 886.730 1771.820 887.050 ;
        RECT 627.140 18.350 627.280 886.730 ;
        RECT 621.100 18.030 621.360 18.350 ;
        RECT 627.080 18.030 627.340 18.350 ;
        RECT 621.160 2.400 621.300 18.030 ;
        RECT 620.950 -4.800 621.510 2.400 ;
      LAYER via2 ;
        RECT 1771.550 1449.960 1771.830 1450.240 ;
      LAYER met3 ;
        RECT 1755.835 1450.250 1759.835 1450.255 ;
        RECT 1771.525 1450.250 1771.855 1450.265 ;
        RECT 1755.835 1449.950 1771.855 1450.250 ;
        RECT 1755.835 1449.655 1759.835 1449.950 ;
        RECT 1771.525 1449.935 1771.855 1449.950 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1504.805 1173.085 1504.975 1207.255 ;
        RECT 1505.725 338.045 1505.895 386.155 ;
        RECT 1505.265 289.765 1505.435 303.875 ;
      LAYER mcon ;
        RECT 1504.805 1207.085 1504.975 1207.255 ;
        RECT 1505.725 385.985 1505.895 386.155 ;
        RECT 1505.265 303.705 1505.435 303.875 ;
      LAYER met1 ;
        RECT 1505.650 1304.480 1505.970 1304.540 ;
        RECT 1510.710 1304.480 1511.030 1304.540 ;
        RECT 1505.650 1304.340 1511.030 1304.480 ;
        RECT 1505.650 1304.280 1505.970 1304.340 ;
        RECT 1510.710 1304.280 1511.030 1304.340 ;
        RECT 1504.730 1293.940 1505.050 1294.000 ;
        RECT 1505.650 1293.940 1505.970 1294.000 ;
        RECT 1504.730 1293.800 1505.970 1293.940 ;
        RECT 1504.730 1293.740 1505.050 1293.800 ;
        RECT 1505.650 1293.740 1505.970 1293.800 ;
        RECT 1504.730 1207.240 1505.050 1207.300 ;
        RECT 1504.535 1207.100 1505.050 1207.240 ;
        RECT 1504.730 1207.040 1505.050 1207.100 ;
        RECT 1504.745 1173.240 1505.035 1173.285 ;
        RECT 1505.650 1173.240 1505.970 1173.300 ;
        RECT 1504.745 1173.100 1505.970 1173.240 ;
        RECT 1504.745 1173.055 1505.035 1173.100 ;
        RECT 1505.650 1173.040 1505.970 1173.100 ;
        RECT 1504.730 1111.020 1505.050 1111.080 ;
        RECT 1506.110 1111.020 1506.430 1111.080 ;
        RECT 1504.730 1110.880 1506.430 1111.020 ;
        RECT 1504.730 1110.820 1505.050 1110.880 ;
        RECT 1506.110 1110.820 1506.430 1110.880 ;
        RECT 1506.110 1077.020 1506.430 1077.080 ;
        RECT 1505.740 1076.880 1506.430 1077.020 ;
        RECT 1505.740 1076.400 1505.880 1076.880 ;
        RECT 1506.110 1076.820 1506.430 1076.880 ;
        RECT 1505.650 1076.140 1505.970 1076.400 ;
        RECT 1504.730 1014.460 1505.050 1014.520 ;
        RECT 1506.110 1014.460 1506.430 1014.520 ;
        RECT 1504.730 1014.320 1506.430 1014.460 ;
        RECT 1504.730 1014.260 1505.050 1014.320 ;
        RECT 1506.110 1014.260 1506.430 1014.320 ;
        RECT 1506.110 980.460 1506.430 980.520 ;
        RECT 1505.740 980.320 1506.430 980.460 ;
        RECT 1505.740 979.840 1505.880 980.320 ;
        RECT 1506.110 980.260 1506.430 980.320 ;
        RECT 1505.650 979.580 1505.970 979.840 ;
        RECT 1504.730 917.900 1505.050 917.960 ;
        RECT 1506.110 917.900 1506.430 917.960 ;
        RECT 1504.730 917.760 1506.430 917.900 ;
        RECT 1504.730 917.700 1505.050 917.760 ;
        RECT 1506.110 917.700 1506.430 917.760 ;
        RECT 1505.190 869.620 1505.510 869.680 ;
        RECT 1506.110 869.620 1506.430 869.680 ;
        RECT 1505.190 869.480 1506.430 869.620 ;
        RECT 1505.190 869.420 1505.510 869.480 ;
        RECT 1506.110 869.420 1506.430 869.480 ;
        RECT 1504.270 759.120 1504.590 759.180 ;
        RECT 1505.190 759.120 1505.510 759.180 ;
        RECT 1504.270 758.980 1505.510 759.120 ;
        RECT 1504.270 758.920 1504.590 758.980 ;
        RECT 1505.190 758.920 1505.510 758.980 ;
        RECT 1505.190 652.020 1505.510 652.080 ;
        RECT 1506.110 652.020 1506.430 652.080 ;
        RECT 1505.190 651.880 1506.430 652.020 ;
        RECT 1505.190 651.820 1505.510 651.880 ;
        RECT 1506.110 651.820 1506.430 651.880 ;
        RECT 1505.190 593.340 1505.510 593.600 ;
        RECT 1505.280 593.200 1505.420 593.340 ;
        RECT 1505.650 593.200 1505.970 593.260 ;
        RECT 1505.280 593.060 1505.970 593.200 ;
        RECT 1505.650 593.000 1505.970 593.060 ;
        RECT 1504.730 545.260 1505.050 545.320 ;
        RECT 1505.650 545.260 1505.970 545.320 ;
        RECT 1504.730 545.120 1505.970 545.260 ;
        RECT 1504.730 545.060 1505.050 545.120 ;
        RECT 1505.650 545.060 1505.970 545.120 ;
        RECT 1505.190 458.900 1505.510 458.960 ;
        RECT 1506.110 458.900 1506.430 458.960 ;
        RECT 1505.190 458.760 1506.430 458.900 ;
        RECT 1505.190 458.700 1505.510 458.760 ;
        RECT 1506.110 458.700 1506.430 458.760 ;
        RECT 1505.190 400.220 1505.510 400.480 ;
        RECT 1505.280 399.740 1505.420 400.220 ;
        RECT 1505.650 399.740 1505.970 399.800 ;
        RECT 1505.280 399.600 1505.970 399.740 ;
        RECT 1505.650 399.540 1505.970 399.600 ;
        RECT 1505.650 386.140 1505.970 386.200 ;
        RECT 1505.455 386.000 1505.970 386.140 ;
        RECT 1505.650 385.940 1505.970 386.000 ;
        RECT 1505.665 338.200 1505.955 338.245 ;
        RECT 1506.110 338.200 1506.430 338.260 ;
        RECT 1505.665 338.060 1506.430 338.200 ;
        RECT 1505.665 338.015 1505.955 338.060 ;
        RECT 1506.110 338.000 1506.430 338.060 ;
        RECT 1505.205 303.860 1505.495 303.905 ;
        RECT 1506.110 303.860 1506.430 303.920 ;
        RECT 1505.205 303.720 1506.430 303.860 ;
        RECT 1505.205 303.675 1505.495 303.720 ;
        RECT 1506.110 303.660 1506.430 303.720 ;
        RECT 1505.190 289.920 1505.510 289.980 ;
        RECT 1504.995 289.780 1505.510 289.920 ;
        RECT 1505.190 289.720 1505.510 289.780 ;
        RECT 1504.270 276.320 1504.590 276.380 ;
        RECT 1505.190 276.320 1505.510 276.380 ;
        RECT 1504.270 276.180 1505.510 276.320 ;
        RECT 1504.270 276.120 1504.590 276.180 ;
        RECT 1505.190 276.120 1505.510 276.180 ;
        RECT 1504.270 179.760 1504.590 179.820 ;
        RECT 1505.190 179.760 1505.510 179.820 ;
        RECT 1504.270 179.620 1505.510 179.760 ;
        RECT 1504.270 179.560 1504.590 179.620 ;
        RECT 1505.190 179.560 1505.510 179.620 ;
        RECT 1504.270 83.200 1504.590 83.260 ;
        RECT 1505.190 83.200 1505.510 83.260 ;
        RECT 1504.270 83.060 1505.510 83.200 ;
        RECT 1504.270 83.000 1504.590 83.060 ;
        RECT 1505.190 83.000 1505.510 83.060 ;
        RECT 115.530 31.520 115.850 31.580 ;
        RECT 1504.730 31.520 1505.050 31.580 ;
        RECT 115.530 31.380 1505.050 31.520 ;
        RECT 115.530 31.320 115.850 31.380 ;
        RECT 1504.730 31.320 1505.050 31.380 ;
      LAYER via ;
        RECT 1505.680 1304.280 1505.940 1304.540 ;
        RECT 1510.740 1304.280 1511.000 1304.540 ;
        RECT 1504.760 1293.740 1505.020 1294.000 ;
        RECT 1505.680 1293.740 1505.940 1294.000 ;
        RECT 1504.760 1207.040 1505.020 1207.300 ;
        RECT 1505.680 1173.040 1505.940 1173.300 ;
        RECT 1504.760 1110.820 1505.020 1111.080 ;
        RECT 1506.140 1110.820 1506.400 1111.080 ;
        RECT 1506.140 1076.820 1506.400 1077.080 ;
        RECT 1505.680 1076.140 1505.940 1076.400 ;
        RECT 1504.760 1014.260 1505.020 1014.520 ;
        RECT 1506.140 1014.260 1506.400 1014.520 ;
        RECT 1506.140 980.260 1506.400 980.520 ;
        RECT 1505.680 979.580 1505.940 979.840 ;
        RECT 1504.760 917.700 1505.020 917.960 ;
        RECT 1506.140 917.700 1506.400 917.960 ;
        RECT 1505.220 869.420 1505.480 869.680 ;
        RECT 1506.140 869.420 1506.400 869.680 ;
        RECT 1504.300 758.920 1504.560 759.180 ;
        RECT 1505.220 758.920 1505.480 759.180 ;
        RECT 1505.220 651.820 1505.480 652.080 ;
        RECT 1506.140 651.820 1506.400 652.080 ;
        RECT 1505.220 593.340 1505.480 593.600 ;
        RECT 1505.680 593.000 1505.940 593.260 ;
        RECT 1504.760 545.060 1505.020 545.320 ;
        RECT 1505.680 545.060 1505.940 545.320 ;
        RECT 1505.220 458.700 1505.480 458.960 ;
        RECT 1506.140 458.700 1506.400 458.960 ;
        RECT 1505.220 400.220 1505.480 400.480 ;
        RECT 1505.680 399.540 1505.940 399.800 ;
        RECT 1505.680 385.940 1505.940 386.200 ;
        RECT 1506.140 338.000 1506.400 338.260 ;
        RECT 1506.140 303.660 1506.400 303.920 ;
        RECT 1505.220 289.720 1505.480 289.980 ;
        RECT 1504.300 276.120 1504.560 276.380 ;
        RECT 1505.220 276.120 1505.480 276.380 ;
        RECT 1504.300 179.560 1504.560 179.820 ;
        RECT 1505.220 179.560 1505.480 179.820 ;
        RECT 1504.300 83.000 1504.560 83.260 ;
        RECT 1505.220 83.000 1505.480 83.260 ;
        RECT 115.560 31.320 115.820 31.580 ;
        RECT 1504.760 31.320 1505.020 31.580 ;
      LAYER met2 ;
        RECT 1510.780 1323.135 1511.060 1327.135 ;
        RECT 1510.800 1304.570 1510.940 1323.135 ;
        RECT 1505.680 1304.250 1505.940 1304.570 ;
        RECT 1510.740 1304.250 1511.000 1304.570 ;
        RECT 1505.740 1294.030 1505.880 1304.250 ;
        RECT 1504.760 1293.710 1505.020 1294.030 ;
        RECT 1505.680 1293.710 1505.940 1294.030 ;
        RECT 1504.820 1280.170 1504.960 1293.710 ;
        RECT 1504.360 1280.030 1504.960 1280.170 ;
        RECT 1504.360 1221.010 1504.500 1280.030 ;
        RECT 1504.360 1220.870 1504.960 1221.010 ;
        RECT 1504.820 1207.330 1504.960 1220.870 ;
        RECT 1504.760 1207.010 1505.020 1207.330 ;
        RECT 1505.680 1173.010 1505.940 1173.330 ;
        RECT 1505.740 1159.245 1505.880 1173.010 ;
        RECT 1504.750 1158.875 1505.030 1159.245 ;
        RECT 1505.670 1158.875 1505.950 1159.245 ;
        RECT 1504.820 1111.110 1504.960 1158.875 ;
        RECT 1504.760 1110.790 1505.020 1111.110 ;
        RECT 1506.140 1110.790 1506.400 1111.110 ;
        RECT 1506.200 1077.110 1506.340 1110.790 ;
        RECT 1506.140 1076.790 1506.400 1077.110 ;
        RECT 1505.680 1076.110 1505.940 1076.430 ;
        RECT 1505.740 1062.685 1505.880 1076.110 ;
        RECT 1504.750 1062.315 1505.030 1062.685 ;
        RECT 1505.670 1062.315 1505.950 1062.685 ;
        RECT 1504.820 1014.550 1504.960 1062.315 ;
        RECT 1504.760 1014.230 1505.020 1014.550 ;
        RECT 1506.140 1014.230 1506.400 1014.550 ;
        RECT 1506.200 980.550 1506.340 1014.230 ;
        RECT 1506.140 980.230 1506.400 980.550 ;
        RECT 1505.680 979.550 1505.940 979.870 ;
        RECT 1505.740 966.125 1505.880 979.550 ;
        RECT 1504.750 965.755 1505.030 966.125 ;
        RECT 1505.670 965.755 1505.950 966.125 ;
        RECT 1504.820 917.990 1504.960 965.755 ;
        RECT 1504.760 917.670 1505.020 917.990 ;
        RECT 1506.140 917.670 1506.400 917.990 ;
        RECT 1506.200 869.710 1506.340 917.670 ;
        RECT 1505.220 869.565 1505.480 869.710 ;
        RECT 1505.210 869.195 1505.490 869.565 ;
        RECT 1506.140 869.390 1506.400 869.710 ;
        RECT 1504.750 820.915 1505.030 821.285 ;
        RECT 1504.820 807.570 1504.960 820.915 ;
        RECT 1504.820 807.430 1505.420 807.570 ;
        RECT 1505.280 759.210 1505.420 807.430 ;
        RECT 1504.300 758.890 1504.560 759.210 ;
        RECT 1505.220 758.890 1505.480 759.210 ;
        RECT 1504.360 758.610 1504.500 758.890 ;
        RECT 1504.360 758.470 1504.960 758.610 ;
        RECT 1504.820 711.010 1504.960 758.470 ;
        RECT 1504.820 710.870 1505.420 711.010 ;
        RECT 1505.280 652.110 1505.420 710.870 ;
        RECT 1505.220 651.790 1505.480 652.110 ;
        RECT 1506.140 651.790 1506.400 652.110 ;
        RECT 1506.200 628.165 1506.340 651.790 ;
        RECT 1505.210 627.795 1505.490 628.165 ;
        RECT 1506.130 627.795 1506.410 628.165 ;
        RECT 1505.280 593.630 1505.420 627.795 ;
        RECT 1505.220 593.310 1505.480 593.630 ;
        RECT 1505.680 592.970 1505.940 593.290 ;
        RECT 1505.740 545.350 1505.880 592.970 ;
        RECT 1504.760 545.030 1505.020 545.350 ;
        RECT 1505.680 545.030 1505.940 545.350 ;
        RECT 1504.820 517.890 1504.960 545.030 ;
        RECT 1504.820 517.750 1505.420 517.890 ;
        RECT 1505.280 458.990 1505.420 517.750 ;
        RECT 1505.220 458.670 1505.480 458.990 ;
        RECT 1506.140 458.670 1506.400 458.990 ;
        RECT 1506.200 435.045 1506.340 458.670 ;
        RECT 1505.210 434.675 1505.490 435.045 ;
        RECT 1506.130 434.675 1506.410 435.045 ;
        RECT 1505.280 400.510 1505.420 434.675 ;
        RECT 1505.220 400.190 1505.480 400.510 ;
        RECT 1505.680 399.510 1505.940 399.830 ;
        RECT 1505.740 386.230 1505.880 399.510 ;
        RECT 1505.680 385.910 1505.940 386.230 ;
        RECT 1506.140 337.970 1506.400 338.290 ;
        RECT 1506.200 303.950 1506.340 337.970 ;
        RECT 1506.140 303.630 1506.400 303.950 ;
        RECT 1505.220 289.690 1505.480 290.010 ;
        RECT 1505.280 276.410 1505.420 289.690 ;
        RECT 1504.300 276.090 1504.560 276.410 ;
        RECT 1505.220 276.090 1505.480 276.410 ;
        RECT 1504.360 275.810 1504.500 276.090 ;
        RECT 1504.360 275.670 1504.960 275.810 ;
        RECT 1504.820 228.210 1504.960 275.670 ;
        RECT 1504.820 228.070 1505.420 228.210 ;
        RECT 1505.280 179.850 1505.420 228.070 ;
        RECT 1504.300 179.530 1504.560 179.850 ;
        RECT 1505.220 179.530 1505.480 179.850 ;
        RECT 1504.360 130.970 1504.500 179.530 ;
        RECT 1504.360 130.830 1505.420 130.970 ;
        RECT 1505.280 83.290 1505.420 130.830 ;
        RECT 1504.300 82.970 1504.560 83.290 ;
        RECT 1505.220 82.970 1505.480 83.290 ;
        RECT 1504.360 82.690 1504.500 82.970 ;
        RECT 1504.360 82.550 1504.960 82.690 ;
        RECT 1504.820 31.610 1504.960 82.550 ;
        RECT 115.560 31.290 115.820 31.610 ;
        RECT 1504.760 31.290 1505.020 31.610 ;
        RECT 115.620 2.400 115.760 31.290 ;
        RECT 115.410 -4.800 115.970 2.400 ;
      LAYER via2 ;
        RECT 1504.750 1158.920 1505.030 1159.200 ;
        RECT 1505.670 1158.920 1505.950 1159.200 ;
        RECT 1504.750 1062.360 1505.030 1062.640 ;
        RECT 1505.670 1062.360 1505.950 1062.640 ;
        RECT 1504.750 965.800 1505.030 966.080 ;
        RECT 1505.670 965.800 1505.950 966.080 ;
        RECT 1505.210 869.240 1505.490 869.520 ;
        RECT 1504.750 820.960 1505.030 821.240 ;
        RECT 1505.210 627.840 1505.490 628.120 ;
        RECT 1506.130 627.840 1506.410 628.120 ;
        RECT 1505.210 434.720 1505.490 435.000 ;
        RECT 1506.130 434.720 1506.410 435.000 ;
      LAYER met3 ;
        RECT 1504.725 1159.210 1505.055 1159.225 ;
        RECT 1505.645 1159.210 1505.975 1159.225 ;
        RECT 1504.725 1158.910 1505.975 1159.210 ;
        RECT 1504.725 1158.895 1505.055 1158.910 ;
        RECT 1505.645 1158.895 1505.975 1158.910 ;
        RECT 1504.725 1062.650 1505.055 1062.665 ;
        RECT 1505.645 1062.650 1505.975 1062.665 ;
        RECT 1504.725 1062.350 1505.975 1062.650 ;
        RECT 1504.725 1062.335 1505.055 1062.350 ;
        RECT 1505.645 1062.335 1505.975 1062.350 ;
        RECT 1504.725 966.090 1505.055 966.105 ;
        RECT 1505.645 966.090 1505.975 966.105 ;
        RECT 1504.725 965.790 1505.975 966.090 ;
        RECT 1504.725 965.775 1505.055 965.790 ;
        RECT 1505.645 965.775 1505.975 965.790 ;
        RECT 1504.470 869.530 1504.850 869.540 ;
        RECT 1505.185 869.530 1505.515 869.545 ;
        RECT 1504.470 869.230 1505.515 869.530 ;
        RECT 1504.470 869.220 1504.850 869.230 ;
        RECT 1505.185 869.215 1505.515 869.230 ;
        RECT 1504.725 821.260 1505.055 821.265 ;
        RECT 1504.470 821.250 1505.055 821.260 ;
        RECT 1504.470 820.950 1505.280 821.250 ;
        RECT 1504.470 820.940 1505.055 820.950 ;
        RECT 1504.725 820.935 1505.055 820.940 ;
        RECT 1505.185 628.130 1505.515 628.145 ;
        RECT 1506.105 628.130 1506.435 628.145 ;
        RECT 1505.185 627.830 1506.435 628.130 ;
        RECT 1505.185 627.815 1505.515 627.830 ;
        RECT 1506.105 627.815 1506.435 627.830 ;
        RECT 1505.185 435.010 1505.515 435.025 ;
        RECT 1506.105 435.010 1506.435 435.025 ;
        RECT 1505.185 434.710 1506.435 435.010 ;
        RECT 1505.185 434.695 1505.515 434.710 ;
        RECT 1506.105 434.695 1506.435 434.710 ;
      LAYER via3 ;
        RECT 1504.500 869.220 1504.820 869.540 ;
        RECT 1504.500 820.940 1504.820 821.260 ;
      LAYER met4 ;
        RECT 1504.495 869.215 1504.825 869.545 ;
        RECT 1504.510 821.265 1504.810 869.215 ;
        RECT 1504.495 820.935 1504.825 821.265 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 144.510 1317.400 144.830 1317.460 ;
        RECT 840.030 1317.400 840.350 1317.460 ;
        RECT 144.510 1317.260 840.350 1317.400 ;
        RECT 144.510 1317.200 144.830 1317.260 ;
        RECT 840.030 1317.200 840.350 1317.260 ;
        RECT 139.450 16.220 139.770 16.280 ;
        RECT 144.510 16.220 144.830 16.280 ;
        RECT 139.450 16.080 144.830 16.220 ;
        RECT 139.450 16.020 139.770 16.080 ;
        RECT 144.510 16.020 144.830 16.080 ;
      LAYER via ;
        RECT 144.540 1317.200 144.800 1317.460 ;
        RECT 840.060 1317.200 840.320 1317.460 ;
        RECT 139.480 16.020 139.740 16.280 ;
        RECT 144.540 16.020 144.800 16.280 ;
      LAYER met2 ;
        RECT 840.100 1323.135 840.380 1327.135 ;
        RECT 840.120 1317.490 840.260 1323.135 ;
        RECT 144.540 1317.170 144.800 1317.490 ;
        RECT 840.060 1317.170 840.320 1317.490 ;
        RECT 144.600 16.310 144.740 1317.170 ;
        RECT 139.480 15.990 139.740 16.310 ;
        RECT 144.540 15.990 144.800 16.310 ;
        RECT 139.540 2.400 139.680 15.990 ;
        RECT 139.330 -4.800 139.890 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1768.330 1886.475 1768.610 1886.845 ;
        RECT 1768.400 1573.365 1768.540 1886.475 ;
        RECT 1768.330 1572.995 1768.610 1573.365 ;
        RECT 157.410 17.835 157.690 18.205 ;
        RECT 157.480 2.400 157.620 17.835 ;
        RECT 157.270 -4.800 157.830 2.400 ;
      LAYER via2 ;
        RECT 1768.330 1886.520 1768.610 1886.800 ;
        RECT 1768.330 1573.040 1768.610 1573.320 ;
        RECT 157.410 17.880 157.690 18.160 ;
      LAYER met3 ;
        RECT 1755.835 1886.810 1759.835 1886.815 ;
        RECT 1768.305 1886.810 1768.635 1886.825 ;
        RECT 1755.835 1886.510 1768.635 1886.810 ;
        RECT 1755.835 1886.215 1759.835 1886.510 ;
        RECT 1768.305 1886.495 1768.635 1886.510 ;
        RECT 1762.990 1573.330 1763.370 1573.340 ;
        RECT 1768.305 1573.330 1768.635 1573.345 ;
        RECT 1762.990 1573.030 1768.635 1573.330 ;
        RECT 1762.990 1573.020 1763.370 1573.030 ;
        RECT 1768.305 1573.015 1768.635 1573.030 ;
        RECT 157.385 18.170 157.715 18.185 ;
        RECT 1762.990 18.170 1763.370 18.180 ;
        RECT 157.385 17.870 1763.370 18.170 ;
        RECT 157.385 17.855 157.715 17.870 ;
        RECT 1762.990 17.860 1763.370 17.870 ;
      LAYER via3 ;
        RECT 1763.020 1573.020 1763.340 1573.340 ;
        RECT 1763.020 17.860 1763.340 18.180 ;
      LAYER met4 ;
        RECT 1763.015 1573.015 1763.345 1573.345 ;
        RECT 1763.030 18.185 1763.330 1573.015 ;
        RECT 1763.015 17.855 1763.345 18.185 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 174.870 32.540 175.190 32.600 ;
        RECT 1311.070 32.540 1311.390 32.600 ;
        RECT 174.870 32.400 1311.390 32.540 ;
        RECT 174.870 32.340 175.190 32.400 ;
        RECT 1311.070 32.340 1311.390 32.400 ;
      LAYER via ;
        RECT 174.900 32.340 175.160 32.600 ;
        RECT 1311.100 32.340 1311.360 32.600 ;
      LAYER met2 ;
        RECT 1313.900 1323.690 1314.180 1327.135 ;
        RECT 1311.160 1323.550 1314.180 1323.690 ;
        RECT 1311.160 32.630 1311.300 1323.550 ;
        RECT 1313.900 1323.135 1314.180 1323.550 ;
        RECT 174.900 32.310 175.160 32.630 ;
        RECT 1311.100 32.310 1311.360 32.630 ;
        RECT 174.960 2.400 175.100 32.310 ;
        RECT 174.750 -4.800 175.310 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 192.810 24.380 193.130 24.440 ;
        RECT 1131.670 24.380 1131.990 24.440 ;
        RECT 192.810 24.240 1131.990 24.380 ;
        RECT 192.810 24.180 193.130 24.240 ;
        RECT 1131.670 24.180 1131.990 24.240 ;
      LAYER via ;
        RECT 192.840 24.180 193.100 24.440 ;
        RECT 1131.700 24.180 1131.960 24.440 ;
      LAYER met2 ;
        RECT 1134.500 1323.690 1134.780 1327.135 ;
        RECT 1131.760 1323.550 1134.780 1323.690 ;
        RECT 1131.760 24.470 1131.900 1323.550 ;
        RECT 1134.500 1323.135 1134.780 1323.550 ;
        RECT 192.840 24.150 193.100 24.470 ;
        RECT 1131.700 24.150 1131.960 24.470 ;
        RECT 192.900 2.400 193.040 24.150 ;
        RECT 192.690 -4.800 193.250 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 210.750 32.880 211.070 32.940 ;
        RECT 1317.970 32.880 1318.290 32.940 ;
        RECT 210.750 32.740 1318.290 32.880 ;
        RECT 210.750 32.680 211.070 32.740 ;
        RECT 1317.970 32.680 1318.290 32.740 ;
      LAYER via ;
        RECT 210.780 32.680 211.040 32.940 ;
        RECT 1318.000 32.680 1318.260 32.940 ;
      LAYER met2 ;
        RECT 1319.420 1323.690 1319.700 1327.135 ;
        RECT 1318.060 1323.550 1319.700 1323.690 ;
        RECT 1318.060 32.970 1318.200 1323.550 ;
        RECT 1319.420 1323.135 1319.700 1323.550 ;
        RECT 210.780 32.650 211.040 32.970 ;
        RECT 1318.000 32.650 1318.260 32.970 ;
        RECT 210.840 2.400 210.980 32.650 ;
        RECT 210.630 -4.800 211.190 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 234.210 2111.640 234.530 2111.700 ;
        RECT 696.970 2111.640 697.290 2111.700 ;
        RECT 234.210 2111.500 697.290 2111.640 ;
        RECT 234.210 2111.440 234.530 2111.500 ;
        RECT 696.970 2111.440 697.290 2111.500 ;
        RECT 228.690 17.240 229.010 17.300 ;
        RECT 234.210 17.240 234.530 17.300 ;
        RECT 228.690 17.100 234.530 17.240 ;
        RECT 228.690 17.040 229.010 17.100 ;
        RECT 234.210 17.040 234.530 17.100 ;
      LAYER via ;
        RECT 234.240 2111.440 234.500 2111.700 ;
        RECT 697.000 2111.440 697.260 2111.700 ;
        RECT 228.720 17.040 228.980 17.300 ;
        RECT 234.240 17.040 234.500 17.300 ;
      LAYER met2 ;
        RECT 696.990 2113.595 697.270 2113.965 ;
        RECT 697.060 2111.730 697.200 2113.595 ;
        RECT 234.240 2111.410 234.500 2111.730 ;
        RECT 697.000 2111.410 697.260 2111.730 ;
        RECT 234.300 17.330 234.440 2111.410 ;
        RECT 228.720 17.010 228.980 17.330 ;
        RECT 234.240 17.010 234.500 17.330 ;
        RECT 228.780 2.400 228.920 17.010 ;
        RECT 228.570 -4.800 229.130 2.400 ;
      LAYER via2 ;
        RECT 696.990 2113.640 697.270 2113.920 ;
      LAYER met3 ;
        RECT 696.965 2113.930 697.295 2113.945 ;
        RECT 715.810 2113.930 719.810 2113.935 ;
        RECT 696.965 2113.630 719.810 2113.930 ;
        RECT 696.965 2113.615 697.295 2113.630 ;
        RECT 715.810 2113.335 719.810 2113.630 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 50.210 37.980 50.530 38.040 ;
        RECT 1580.170 37.980 1580.490 38.040 ;
        RECT 50.210 37.840 1580.490 37.980 ;
        RECT 50.210 37.780 50.530 37.840 ;
        RECT 1580.170 37.780 1580.490 37.840 ;
      LAYER via ;
        RECT 50.240 37.780 50.500 38.040 ;
        RECT 1580.200 37.780 1580.460 38.040 ;
      LAYER met2 ;
        RECT 1586.220 1323.690 1586.500 1327.135 ;
        RECT 1580.260 1323.550 1586.500 1323.690 ;
        RECT 1580.260 38.070 1580.400 1323.550 ;
        RECT 1586.220 1323.135 1586.500 1323.550 ;
        RECT 50.240 37.750 50.500 38.070 ;
        RECT 1580.200 37.750 1580.460 38.070 ;
        RECT 50.300 2.400 50.440 37.750 ;
        RECT 50.090 -4.800 50.650 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 252.610 18.260 252.930 18.320 ;
        RECT 548.390 18.260 548.710 18.320 ;
        RECT 252.610 18.120 548.710 18.260 ;
        RECT 252.610 18.060 252.930 18.120 ;
        RECT 548.390 18.060 548.710 18.120 ;
      LAYER via ;
        RECT 252.640 18.060 252.900 18.320 ;
        RECT 548.420 18.060 548.680 18.320 ;
      LAYER met2 ;
        RECT 548.410 2390.355 548.690 2390.725 ;
        RECT 1300.050 2390.355 1300.330 2390.725 ;
        RECT 548.480 18.350 548.620 2390.355 ;
        RECT 1300.120 2377.880 1300.260 2390.355 ;
        RECT 1300.100 2373.880 1300.380 2377.880 ;
        RECT 252.640 18.030 252.900 18.350 ;
        RECT 548.420 18.030 548.680 18.350 ;
        RECT 252.700 2.400 252.840 18.030 ;
        RECT 252.490 -4.800 253.050 2.400 ;
      LAYER via2 ;
        RECT 548.410 2390.400 548.690 2390.680 ;
        RECT 1300.050 2390.400 1300.330 2390.680 ;
      LAYER met3 ;
        RECT 548.385 2390.690 548.715 2390.705 ;
        RECT 1300.025 2390.690 1300.355 2390.705 ;
        RECT 548.385 2390.390 1300.355 2390.690 ;
        RECT 548.385 2390.375 548.715 2390.390 ;
        RECT 1300.025 2390.375 1300.355 2390.390 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 275.610 1316.380 275.930 1316.440 ;
        RECT 989.990 1316.380 990.310 1316.440 ;
        RECT 275.610 1316.240 990.310 1316.380 ;
        RECT 275.610 1316.180 275.930 1316.240 ;
        RECT 989.990 1316.180 990.310 1316.240 ;
        RECT 270.090 16.900 270.410 16.960 ;
        RECT 275.610 16.900 275.930 16.960 ;
        RECT 270.090 16.760 275.930 16.900 ;
        RECT 270.090 16.700 270.410 16.760 ;
        RECT 275.610 16.700 275.930 16.760 ;
      LAYER via ;
        RECT 275.640 1316.180 275.900 1316.440 ;
        RECT 990.020 1316.180 990.280 1316.440 ;
        RECT 270.120 16.700 270.380 16.960 ;
        RECT 275.640 16.700 275.900 16.960 ;
      LAYER met2 ;
        RECT 990.060 1323.135 990.340 1327.135 ;
        RECT 990.080 1316.470 990.220 1323.135 ;
        RECT 275.640 1316.150 275.900 1316.470 ;
        RECT 990.020 1316.150 990.280 1316.470 ;
        RECT 275.700 16.990 275.840 1316.150 ;
        RECT 270.120 16.670 270.380 16.990 ;
        RECT 275.640 16.670 275.900 16.990 ;
        RECT 270.180 2.400 270.320 16.670 ;
        RECT 269.970 -4.800 270.530 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 697.965 2387.225 698.135 2390.455 ;
        RECT 726.025 2387.225 726.195 2390.795 ;
        RECT 759.145 2387.225 759.315 2390.795 ;
        RECT 786.745 2387.225 786.915 2390.795 ;
        RECT 952.345 2387.905 952.515 2390.795 ;
        RECT 976.725 2388.075 976.895 2388.415 ;
        RECT 1000.185 2388.245 1000.355 2390.795 ;
        RECT 1049.405 2390.625 1049.575 2392.835 ;
        RECT 1096.325 2390.625 1096.495 2392.835 ;
        RECT 974.885 2387.905 976.895 2388.075 ;
        RECT 541.565 16.065 541.735 19.295 ;
      LAYER mcon ;
        RECT 1049.405 2392.665 1049.575 2392.835 ;
        RECT 726.025 2390.625 726.195 2390.795 ;
        RECT 697.965 2390.285 698.135 2390.455 ;
        RECT 759.145 2390.625 759.315 2390.795 ;
        RECT 786.745 2390.625 786.915 2390.795 ;
        RECT 952.345 2390.625 952.515 2390.795 ;
        RECT 1000.185 2390.625 1000.355 2390.795 ;
        RECT 1096.325 2392.665 1096.495 2392.835 ;
        RECT 976.725 2388.245 976.895 2388.415 ;
        RECT 541.565 19.125 541.735 19.295 ;
      LAYER met1 ;
        RECT 1049.345 2392.820 1049.635 2392.865 ;
        RECT 1096.265 2392.820 1096.555 2392.865 ;
        RECT 1049.345 2392.680 1096.555 2392.820 ;
        RECT 1049.345 2392.635 1049.635 2392.680 ;
        RECT 1096.265 2392.635 1096.555 2392.680 ;
        RECT 569.090 2390.780 569.410 2390.840 ;
        RECT 725.965 2390.780 726.255 2390.825 ;
        RECT 759.085 2390.780 759.375 2390.825 ;
        RECT 569.090 2390.640 614.400 2390.780 ;
        RECT 569.090 2390.580 569.410 2390.640 ;
        RECT 614.260 2390.440 614.400 2390.640 ;
        RECT 725.965 2390.640 759.375 2390.780 ;
        RECT 725.965 2390.595 726.255 2390.640 ;
        RECT 759.085 2390.595 759.375 2390.640 ;
        RECT 786.685 2390.780 786.975 2390.825 ;
        RECT 855.670 2390.780 855.990 2390.840 ;
        RECT 786.685 2390.640 855.990 2390.780 ;
        RECT 786.685 2390.595 786.975 2390.640 ;
        RECT 855.670 2390.580 855.990 2390.640 ;
        RECT 903.510 2390.780 903.830 2390.840 ;
        RECT 952.285 2390.780 952.575 2390.825 ;
        RECT 903.510 2390.640 952.575 2390.780 ;
        RECT 903.510 2390.580 903.830 2390.640 ;
        RECT 952.285 2390.595 952.575 2390.640 ;
        RECT 1000.125 2390.780 1000.415 2390.825 ;
        RECT 1049.345 2390.780 1049.635 2390.825 ;
        RECT 1000.125 2390.640 1049.635 2390.780 ;
        RECT 1000.125 2390.595 1000.415 2390.640 ;
        RECT 1049.345 2390.595 1049.635 2390.640 ;
        RECT 1096.265 2390.780 1096.555 2390.825 ;
        RECT 1120.630 2390.780 1120.950 2390.840 ;
        RECT 1096.265 2390.640 1120.950 2390.780 ;
        RECT 1096.265 2390.595 1096.555 2390.640 ;
        RECT 1120.630 2390.580 1120.950 2390.640 ;
        RECT 697.905 2390.440 698.195 2390.485 ;
        RECT 614.260 2390.300 698.195 2390.440 ;
        RECT 697.905 2390.255 698.195 2390.300 ;
        RECT 976.665 2388.400 976.955 2388.445 ;
        RECT 1000.125 2388.400 1000.415 2388.445 ;
        RECT 976.665 2388.260 1000.415 2388.400 ;
        RECT 976.665 2388.215 976.955 2388.260 ;
        RECT 1000.125 2388.215 1000.415 2388.260 ;
        RECT 855.670 2388.060 855.990 2388.120 ;
        RECT 903.510 2388.060 903.830 2388.120 ;
        RECT 855.670 2387.920 903.830 2388.060 ;
        RECT 855.670 2387.860 855.990 2387.920 ;
        RECT 903.510 2387.860 903.830 2387.920 ;
        RECT 952.285 2388.060 952.575 2388.105 ;
        RECT 974.825 2388.060 975.115 2388.105 ;
        RECT 952.285 2387.920 975.115 2388.060 ;
        RECT 952.285 2387.875 952.575 2387.920 ;
        RECT 974.825 2387.875 975.115 2387.920 ;
        RECT 697.905 2387.380 698.195 2387.425 ;
        RECT 725.965 2387.380 726.255 2387.425 ;
        RECT 697.905 2387.240 726.255 2387.380 ;
        RECT 697.905 2387.195 698.195 2387.240 ;
        RECT 725.965 2387.195 726.255 2387.240 ;
        RECT 759.085 2387.380 759.375 2387.425 ;
        RECT 786.685 2387.380 786.975 2387.425 ;
        RECT 759.085 2387.240 786.975 2387.380 ;
        RECT 759.085 2387.195 759.375 2387.240 ;
        RECT 786.685 2387.195 786.975 2387.240 ;
        RECT 288.030 19.280 288.350 19.340 ;
        RECT 541.505 19.280 541.795 19.325 ;
        RECT 288.030 19.140 541.795 19.280 ;
        RECT 288.030 19.080 288.350 19.140 ;
        RECT 541.505 19.095 541.795 19.140 ;
        RECT 541.505 16.220 541.795 16.265 ;
        RECT 569.090 16.220 569.410 16.280 ;
        RECT 541.505 16.080 569.410 16.220 ;
        RECT 541.505 16.035 541.795 16.080 ;
        RECT 569.090 16.020 569.410 16.080 ;
      LAYER via ;
        RECT 569.120 2390.580 569.380 2390.840 ;
        RECT 855.700 2390.580 855.960 2390.840 ;
        RECT 903.540 2390.580 903.800 2390.840 ;
        RECT 1120.660 2390.580 1120.920 2390.840 ;
        RECT 855.700 2387.860 855.960 2388.120 ;
        RECT 903.540 2387.860 903.800 2388.120 ;
        RECT 288.060 19.080 288.320 19.340 ;
        RECT 569.120 16.020 569.380 16.280 ;
      LAYER met2 ;
        RECT 569.120 2390.550 569.380 2390.870 ;
        RECT 855.700 2390.550 855.960 2390.870 ;
        RECT 903.540 2390.550 903.800 2390.870 ;
        RECT 1120.660 2390.550 1120.920 2390.870 ;
        RECT 288.060 19.050 288.320 19.370 ;
        RECT 288.120 2.400 288.260 19.050 ;
        RECT 569.180 16.310 569.320 2390.550 ;
        RECT 855.760 2388.150 855.900 2390.550 ;
        RECT 903.600 2388.150 903.740 2390.550 ;
        RECT 855.700 2387.830 855.960 2388.150 ;
        RECT 903.540 2387.830 903.800 2388.150 ;
        RECT 1120.720 2377.880 1120.860 2390.550 ;
        RECT 1120.700 2373.880 1120.980 2377.880 ;
        RECT 569.120 15.990 569.380 16.310 ;
        RECT 287.910 -4.800 288.470 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 800.010 2389.420 800.330 2389.480 ;
        RECT 1588.910 2389.420 1589.230 2389.480 ;
        RECT 800.010 2389.280 1589.230 2389.420 ;
        RECT 800.010 2389.220 800.330 2389.280 ;
        RECT 1588.910 2389.220 1589.230 2389.280 ;
        RECT 305.970 18.600 306.290 18.660 ;
        RECT 603.590 18.600 603.910 18.660 ;
        RECT 305.970 18.460 603.910 18.600 ;
        RECT 305.970 18.400 306.290 18.460 ;
        RECT 603.590 18.400 603.910 18.460 ;
      LAYER via ;
        RECT 800.040 2389.220 800.300 2389.480 ;
        RECT 1588.940 2389.220 1589.200 2389.480 ;
        RECT 306.000 18.400 306.260 18.660 ;
        RECT 603.620 18.400 603.880 18.660 ;
      LAYER met2 ;
        RECT 603.610 2393.755 603.890 2394.125 ;
        RECT 787.150 2393.755 787.430 2394.125 ;
        RECT 603.680 18.690 603.820 2393.755 ;
        RECT 787.220 2392.085 787.360 2393.755 ;
        RECT 787.150 2391.715 787.430 2392.085 ;
        RECT 800.030 2391.715 800.310 2392.085 ;
        RECT 800.100 2389.510 800.240 2391.715 ;
        RECT 800.040 2389.190 800.300 2389.510 ;
        RECT 1588.940 2389.190 1589.200 2389.510 ;
        RECT 1589.000 2377.880 1589.140 2389.190 ;
        RECT 1588.980 2373.880 1589.260 2377.880 ;
        RECT 306.000 18.370 306.260 18.690 ;
        RECT 603.620 18.370 603.880 18.690 ;
        RECT 306.060 2.400 306.200 18.370 ;
        RECT 305.850 -4.800 306.410 2.400 ;
      LAYER via2 ;
        RECT 603.610 2393.800 603.890 2394.080 ;
        RECT 787.150 2393.800 787.430 2394.080 ;
        RECT 787.150 2391.760 787.430 2392.040 ;
        RECT 800.030 2391.760 800.310 2392.040 ;
      LAYER met3 ;
        RECT 603.585 2394.090 603.915 2394.105 ;
        RECT 787.125 2394.090 787.455 2394.105 ;
        RECT 603.585 2393.790 787.455 2394.090 ;
        RECT 603.585 2393.775 603.915 2393.790 ;
        RECT 787.125 2393.775 787.455 2393.790 ;
        RECT 787.125 2392.050 787.455 2392.065 ;
        RECT 800.005 2392.050 800.335 2392.065 ;
        RECT 787.125 2391.750 800.335 2392.050 ;
        RECT 787.125 2391.735 787.455 2391.750 ;
        RECT 800.005 2391.735 800.335 2391.750 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 323.910 2001.140 324.230 2001.200 ;
        RECT 699.730 2001.140 700.050 2001.200 ;
        RECT 323.910 2001.000 700.050 2001.140 ;
        RECT 323.910 2000.940 324.230 2001.000 ;
        RECT 699.730 2000.940 700.050 2001.000 ;
      LAYER via ;
        RECT 323.940 2000.940 324.200 2001.200 ;
        RECT 699.760 2000.940 700.020 2001.200 ;
      LAYER met2 ;
        RECT 699.750 2002.075 700.030 2002.445 ;
        RECT 699.820 2001.230 699.960 2002.075 ;
        RECT 323.940 2000.910 324.200 2001.230 ;
        RECT 699.760 2000.910 700.020 2001.230 ;
        RECT 324.000 2.400 324.140 2000.910 ;
        RECT 323.790 -4.800 324.350 2.400 ;
      LAYER via2 ;
        RECT 699.750 2002.120 700.030 2002.400 ;
      LAYER met3 ;
        RECT 699.725 2002.410 700.055 2002.425 ;
        RECT 715.810 2002.410 719.810 2002.415 ;
        RECT 699.725 2002.110 719.810 2002.410 ;
        RECT 699.725 2002.095 700.055 2002.110 ;
        RECT 715.810 2001.815 719.810 2002.110 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 348.290 2388.740 348.610 2388.800 ;
        RECT 1166.170 2388.740 1166.490 2388.800 ;
        RECT 348.290 2388.600 1166.490 2388.740 ;
        RECT 348.290 2388.540 348.610 2388.600 ;
        RECT 1166.170 2388.540 1166.490 2388.600 ;
        RECT 341.390 16.560 341.710 16.620 ;
        RECT 348.290 16.560 348.610 16.620 ;
        RECT 341.390 16.420 348.610 16.560 ;
        RECT 341.390 16.360 341.710 16.420 ;
        RECT 348.290 16.360 348.610 16.420 ;
      LAYER via ;
        RECT 348.320 2388.540 348.580 2388.800 ;
        RECT 1166.200 2388.540 1166.460 2388.800 ;
        RECT 341.420 16.360 341.680 16.620 ;
        RECT 348.320 16.360 348.580 16.620 ;
      LAYER met2 ;
        RECT 1166.260 2389.110 1167.320 2389.250 ;
        RECT 1166.260 2388.830 1166.400 2389.110 ;
        RECT 348.320 2388.510 348.580 2388.830 ;
        RECT 1166.200 2388.510 1166.460 2388.830 ;
        RECT 348.380 16.650 348.520 2388.510 ;
        RECT 1167.180 2377.690 1167.320 2389.110 ;
        RECT 1172.220 2377.690 1172.500 2377.880 ;
        RECT 1167.180 2377.550 1172.500 2377.690 ;
        RECT 1172.220 2373.880 1172.500 2377.550 ;
        RECT 341.420 16.330 341.680 16.650 ;
        RECT 348.320 16.330 348.580 16.650 ;
        RECT 341.480 2.400 341.620 16.330 ;
        RECT 341.270 -4.800 341.830 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 359.330 39.340 359.650 39.400 ;
        RECT 1614.670 39.340 1614.990 39.400 ;
        RECT 359.330 39.200 1614.990 39.340 ;
        RECT 359.330 39.140 359.650 39.200 ;
        RECT 1614.670 39.140 1614.990 39.200 ;
      LAYER via ;
        RECT 359.360 39.140 359.620 39.400 ;
        RECT 1614.700 39.140 1614.960 39.400 ;
      LAYER met2 ;
        RECT 1614.740 1323.135 1615.020 1327.135 ;
        RECT 1614.760 39.430 1614.900 1323.135 ;
        RECT 359.360 39.110 359.620 39.430 ;
        RECT 1614.700 39.110 1614.960 39.430 ;
        RECT 359.420 2.400 359.560 39.110 ;
        RECT 359.210 -4.800 359.770 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 379.110 1863.100 379.430 1863.160 ;
        RECT 704.330 1863.100 704.650 1863.160 ;
        RECT 379.110 1862.960 704.650 1863.100 ;
        RECT 379.110 1862.900 379.430 1862.960 ;
        RECT 704.330 1862.900 704.650 1862.960 ;
      LAYER via ;
        RECT 379.140 1862.900 379.400 1863.160 ;
        RECT 704.360 1862.900 704.620 1863.160 ;
      LAYER met2 ;
        RECT 704.350 1866.075 704.630 1866.445 ;
        RECT 704.420 1863.190 704.560 1866.075 ;
        RECT 379.140 1862.870 379.400 1863.190 ;
        RECT 704.360 1862.870 704.620 1863.190 ;
        RECT 379.200 17.410 379.340 1862.870 ;
        RECT 377.360 17.270 379.340 17.410 ;
        RECT 377.360 2.400 377.500 17.270 ;
        RECT 377.150 -4.800 377.710 2.400 ;
      LAYER via2 ;
        RECT 704.350 1866.120 704.630 1866.400 ;
      LAYER met3 ;
        RECT 704.325 1866.410 704.655 1866.425 ;
        RECT 715.810 1866.410 719.810 1866.415 ;
        RECT 704.325 1866.110 719.810 1866.410 ;
        RECT 704.325 1866.095 704.655 1866.110 ;
        RECT 715.810 1865.815 719.810 1866.110 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 395.210 39.000 395.530 39.060 ;
        RECT 1691.030 39.000 1691.350 39.060 ;
        RECT 395.210 38.860 1691.350 39.000 ;
        RECT 395.210 38.800 395.530 38.860 ;
        RECT 1691.030 38.800 1691.350 38.860 ;
      LAYER via ;
        RECT 395.240 38.800 395.500 39.060 ;
        RECT 1691.060 38.800 1691.320 39.060 ;
      LAYER met2 ;
        RECT 1695.700 1323.690 1695.980 1327.135 ;
        RECT 1691.120 1323.550 1695.980 1323.690 ;
        RECT 1691.120 39.090 1691.260 1323.550 ;
        RECT 1695.700 1323.135 1695.980 1323.550 ;
        RECT 395.240 38.770 395.500 39.090 ;
        RECT 1691.060 38.770 1691.320 39.090 ;
        RECT 395.300 2.400 395.440 38.770 ;
        RECT 395.090 -4.800 395.650 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 458.690 1317.060 459.010 1317.120 ;
        RECT 1227.350 1317.060 1227.670 1317.120 ;
        RECT 458.690 1316.920 1227.670 1317.060 ;
        RECT 458.690 1316.860 459.010 1316.920 ;
        RECT 1227.350 1316.860 1227.670 1316.920 ;
        RECT 413.150 18.940 413.470 19.000 ;
        RECT 458.690 18.940 459.010 19.000 ;
        RECT 413.150 18.800 459.010 18.940 ;
        RECT 413.150 18.740 413.470 18.800 ;
        RECT 458.690 18.740 459.010 18.800 ;
      LAYER via ;
        RECT 458.720 1316.860 458.980 1317.120 ;
        RECT 1227.380 1316.860 1227.640 1317.120 ;
        RECT 413.180 18.740 413.440 19.000 ;
        RECT 458.720 18.740 458.980 19.000 ;
      LAYER met2 ;
        RECT 1227.420 1323.135 1227.700 1327.135 ;
        RECT 1227.440 1317.150 1227.580 1323.135 ;
        RECT 458.720 1316.830 458.980 1317.150 ;
        RECT 1227.380 1316.830 1227.640 1317.150 ;
        RECT 458.780 19.030 458.920 1316.830 ;
        RECT 413.180 18.710 413.440 19.030 ;
        RECT 458.720 18.710 458.980 19.030 ;
        RECT 413.240 2.400 413.380 18.710 ;
        RECT 413.030 -4.800 413.590 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 75.510 1642.440 75.830 1642.500 ;
        RECT 699.730 1642.440 700.050 1642.500 ;
        RECT 75.510 1642.300 700.050 1642.440 ;
        RECT 75.510 1642.240 75.830 1642.300 ;
        RECT 699.730 1642.240 700.050 1642.300 ;
      LAYER via ;
        RECT 75.540 1642.240 75.800 1642.500 ;
        RECT 699.760 1642.240 700.020 1642.500 ;
      LAYER met2 ;
        RECT 699.750 1643.035 700.030 1643.405 ;
        RECT 699.820 1642.530 699.960 1643.035 ;
        RECT 75.540 1642.210 75.800 1642.530 ;
        RECT 699.760 1642.210 700.020 1642.530 ;
        RECT 75.600 17.410 75.740 1642.210 ;
        RECT 74.220 17.270 75.740 17.410 ;
        RECT 74.220 2.400 74.360 17.270 ;
        RECT 74.010 -4.800 74.570 2.400 ;
      LAYER via2 ;
        RECT 699.750 1643.080 700.030 1643.360 ;
      LAYER met3 ;
        RECT 699.725 1643.370 700.055 1643.385 ;
        RECT 715.810 1643.370 719.810 1643.375 ;
        RECT 699.725 1643.070 719.810 1643.370 ;
        RECT 699.725 1643.055 700.055 1643.070 ;
        RECT 715.810 1642.775 719.810 1643.070 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 672.590 2388.060 672.910 2388.120 ;
        RECT 825.310 2388.060 825.630 2388.120 ;
        RECT 672.590 2387.920 825.630 2388.060 ;
        RECT 672.590 2387.860 672.910 2387.920 ;
        RECT 825.310 2387.860 825.630 2387.920 ;
        RECT 430.630 19.620 430.950 19.680 ;
        RECT 672.590 19.620 672.910 19.680 ;
        RECT 430.630 19.480 672.910 19.620 ;
        RECT 430.630 19.420 430.950 19.480 ;
        RECT 672.590 19.420 672.910 19.480 ;
      LAYER via ;
        RECT 672.620 2387.860 672.880 2388.120 ;
        RECT 825.340 2387.860 825.600 2388.120 ;
        RECT 430.660 19.420 430.920 19.680 ;
        RECT 672.620 19.420 672.880 19.680 ;
      LAYER met2 ;
        RECT 672.620 2387.830 672.880 2388.150 ;
        RECT 825.340 2387.830 825.600 2388.150 ;
        RECT 672.680 19.710 672.820 2387.830 ;
        RECT 825.400 2377.880 825.540 2387.830 ;
        RECT 825.380 2373.880 825.660 2377.880 ;
        RECT 430.660 19.390 430.920 19.710 ;
        RECT 672.620 19.390 672.880 19.710 ;
        RECT 430.720 2.400 430.860 19.390 ;
        RECT 430.510 -4.800 431.070 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 455.010 2381.600 455.330 2381.660 ;
        RECT 1727.830 2381.600 1728.150 2381.660 ;
        RECT 455.010 2381.460 1728.150 2381.600 ;
        RECT 455.010 2381.400 455.330 2381.460 ;
        RECT 1727.830 2381.400 1728.150 2381.460 ;
        RECT 448.570 15.200 448.890 15.260 ;
        RECT 455.010 15.200 455.330 15.260 ;
        RECT 448.570 15.060 455.330 15.200 ;
        RECT 448.570 15.000 448.890 15.060 ;
        RECT 455.010 15.000 455.330 15.060 ;
      LAYER via ;
        RECT 455.040 2381.400 455.300 2381.660 ;
        RECT 1727.860 2381.400 1728.120 2381.660 ;
        RECT 448.600 15.000 448.860 15.260 ;
        RECT 455.040 15.000 455.300 15.260 ;
      LAYER met2 ;
        RECT 455.040 2381.370 455.300 2381.690 ;
        RECT 1727.860 2381.370 1728.120 2381.690 ;
        RECT 455.100 15.290 455.240 2381.370 ;
        RECT 1727.920 2377.880 1728.060 2381.370 ;
        RECT 1727.900 2373.880 1728.180 2377.880 ;
        RECT 448.600 14.970 448.860 15.290 ;
        RECT 455.040 14.970 455.300 15.290 ;
        RECT 448.660 2.400 448.800 14.970 ;
        RECT 448.450 -4.800 449.010 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1279.790 1311.280 1280.110 1311.340 ;
        RECT 1285.310 1311.280 1285.630 1311.340 ;
        RECT 1279.790 1311.140 1285.630 1311.280 ;
        RECT 1279.790 1311.080 1280.110 1311.140 ;
        RECT 1285.310 1311.080 1285.630 1311.140 ;
        RECT 466.510 18.940 466.830 19.000 ;
        RECT 1279.790 18.940 1280.110 19.000 ;
        RECT 466.510 18.800 1280.110 18.940 ;
        RECT 466.510 18.740 466.830 18.800 ;
        RECT 1279.790 18.740 1280.110 18.800 ;
      LAYER via ;
        RECT 1279.820 1311.080 1280.080 1311.340 ;
        RECT 1285.340 1311.080 1285.600 1311.340 ;
        RECT 466.540 18.740 466.800 19.000 ;
        RECT 1279.820 18.740 1280.080 19.000 ;
      LAYER met2 ;
        RECT 1285.380 1323.135 1285.660 1327.135 ;
        RECT 1285.400 1311.370 1285.540 1323.135 ;
        RECT 1279.820 1311.050 1280.080 1311.370 ;
        RECT 1285.340 1311.050 1285.600 1311.370 ;
        RECT 1279.880 19.030 1280.020 1311.050 ;
        RECT 466.540 18.710 466.800 19.030 ;
        RECT 1279.820 18.710 1280.080 19.030 ;
        RECT 466.600 2.400 466.740 18.710 ;
        RECT 466.390 -4.800 466.950 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 489.510 1312.300 489.830 1312.360 ;
        RECT 822.550 1312.300 822.870 1312.360 ;
        RECT 489.510 1312.160 822.870 1312.300 ;
        RECT 489.510 1312.100 489.830 1312.160 ;
        RECT 822.550 1312.100 822.870 1312.160 ;
        RECT 484.450 16.900 484.770 16.960 ;
        RECT 489.510 16.900 489.830 16.960 ;
        RECT 484.450 16.760 489.830 16.900 ;
        RECT 484.450 16.700 484.770 16.760 ;
        RECT 489.510 16.700 489.830 16.760 ;
      LAYER via ;
        RECT 489.540 1312.100 489.800 1312.360 ;
        RECT 822.580 1312.100 822.840 1312.360 ;
        RECT 484.480 16.700 484.740 16.960 ;
        RECT 489.540 16.700 489.800 16.960 ;
      LAYER met2 ;
        RECT 822.620 1323.135 822.900 1327.135 ;
        RECT 822.640 1312.390 822.780 1323.135 ;
        RECT 489.540 1312.070 489.800 1312.390 ;
        RECT 822.580 1312.070 822.840 1312.390 ;
        RECT 489.600 16.990 489.740 1312.070 ;
        RECT 484.480 16.670 484.740 16.990 ;
        RECT 489.540 16.670 489.800 16.990 ;
        RECT 484.540 2.400 484.680 16.670 ;
        RECT 484.330 -4.800 484.890 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 503.310 2383.300 503.630 2383.360 ;
        RECT 1606.390 2383.300 1606.710 2383.360 ;
        RECT 503.310 2383.160 1606.710 2383.300 ;
        RECT 503.310 2383.100 503.630 2383.160 ;
        RECT 1606.390 2383.100 1606.710 2383.160 ;
      LAYER via ;
        RECT 503.340 2383.100 503.600 2383.360 ;
        RECT 1606.420 2383.100 1606.680 2383.360 ;
      LAYER met2 ;
        RECT 503.340 2383.070 503.600 2383.390 ;
        RECT 1606.420 2383.070 1606.680 2383.390 ;
        RECT 503.400 17.410 503.540 2383.070 ;
        RECT 1606.480 2377.880 1606.620 2383.070 ;
        RECT 1606.460 2373.880 1606.740 2377.880 ;
        RECT 502.480 17.270 503.540 17.410 ;
        RECT 502.480 2.400 502.620 17.270 ;
        RECT 502.270 -4.800 502.830 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 617.390 2392.480 617.710 2392.540 ;
        RECT 952.270 2392.480 952.590 2392.540 ;
        RECT 617.390 2392.340 952.590 2392.480 ;
        RECT 617.390 2392.280 617.710 2392.340 ;
        RECT 952.270 2392.280 952.590 2392.340 ;
        RECT 519.870 16.900 520.190 16.960 ;
        RECT 617.390 16.900 617.710 16.960 ;
        RECT 519.870 16.760 617.710 16.900 ;
        RECT 519.870 16.700 520.190 16.760 ;
        RECT 617.390 16.700 617.710 16.760 ;
      LAYER via ;
        RECT 617.420 2392.280 617.680 2392.540 ;
        RECT 952.300 2392.280 952.560 2392.540 ;
        RECT 519.900 16.700 520.160 16.960 ;
        RECT 617.420 16.700 617.680 16.960 ;
      LAYER met2 ;
        RECT 617.420 2392.250 617.680 2392.570 ;
        RECT 952.300 2392.250 952.560 2392.570 ;
        RECT 617.480 16.990 617.620 2392.250 ;
        RECT 952.360 2377.880 952.500 2392.250 ;
        RECT 952.340 2373.880 952.620 2377.880 ;
        RECT 519.900 16.670 520.160 16.990 ;
        RECT 617.420 16.670 617.680 16.990 ;
        RECT 519.960 2.400 520.100 16.670 ;
        RECT 519.750 -4.800 520.310 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 589.790 2392.140 590.110 2392.200 ;
        RECT 1085.670 2392.140 1085.990 2392.200 ;
        RECT 589.790 2392.000 1085.990 2392.140 ;
        RECT 589.790 2391.940 590.110 2392.000 ;
        RECT 1085.670 2391.940 1085.990 2392.000 ;
        RECT 537.810 16.560 538.130 16.620 ;
        RECT 589.790 16.560 590.110 16.620 ;
        RECT 537.810 16.420 590.110 16.560 ;
        RECT 537.810 16.360 538.130 16.420 ;
        RECT 589.790 16.360 590.110 16.420 ;
      LAYER via ;
        RECT 589.820 2391.940 590.080 2392.200 ;
        RECT 1085.700 2391.940 1085.960 2392.200 ;
        RECT 537.840 16.360 538.100 16.620 ;
        RECT 589.820 16.360 590.080 16.620 ;
      LAYER met2 ;
        RECT 589.820 2391.910 590.080 2392.230 ;
        RECT 1085.700 2391.910 1085.960 2392.230 ;
        RECT 589.880 16.650 590.020 2391.910 ;
        RECT 1085.760 2377.880 1085.900 2391.910 ;
        RECT 1085.740 2373.880 1086.020 2377.880 ;
        RECT 537.840 16.330 538.100 16.650 ;
        RECT 589.820 16.330 590.080 16.650 ;
        RECT 537.900 2.400 538.040 16.330 ;
        RECT 537.690 -4.800 538.250 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 558.510 1311.960 558.830 1312.020 ;
        RECT 851.070 1311.960 851.390 1312.020 ;
        RECT 558.510 1311.820 851.390 1311.960 ;
        RECT 558.510 1311.760 558.830 1311.820 ;
        RECT 851.070 1311.760 851.390 1311.820 ;
        RECT 555.750 17.240 556.070 17.300 ;
        RECT 558.510 17.240 558.830 17.300 ;
        RECT 555.750 17.100 558.830 17.240 ;
        RECT 555.750 17.040 556.070 17.100 ;
        RECT 558.510 17.040 558.830 17.100 ;
      LAYER via ;
        RECT 558.540 1311.760 558.800 1312.020 ;
        RECT 851.100 1311.760 851.360 1312.020 ;
        RECT 555.780 17.040 556.040 17.300 ;
        RECT 558.540 17.040 558.800 17.300 ;
      LAYER met2 ;
        RECT 851.140 1323.135 851.420 1327.135 ;
        RECT 851.160 1312.050 851.300 1323.135 ;
        RECT 558.540 1311.730 558.800 1312.050 ;
        RECT 851.100 1311.730 851.360 1312.050 ;
        RECT 558.600 17.330 558.740 1311.730 ;
        RECT 555.780 17.010 556.040 17.330 ;
        RECT 558.540 17.010 558.800 17.330 ;
        RECT 555.840 2.400 555.980 17.010 ;
        RECT 555.630 -4.800 556.190 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 579.210 886.620 579.530 886.680 ;
        RECT 1762.330 886.620 1762.650 886.680 ;
        RECT 579.210 886.480 1762.650 886.620 ;
        RECT 579.210 886.420 579.530 886.480 ;
        RECT 1762.330 886.420 1762.650 886.480 ;
        RECT 573.690 15.200 574.010 15.260 ;
        RECT 579.210 15.200 579.530 15.260 ;
        RECT 573.690 15.060 579.530 15.200 ;
        RECT 573.690 15.000 574.010 15.060 ;
        RECT 579.210 15.000 579.530 15.060 ;
      LAYER via ;
        RECT 579.240 886.420 579.500 886.680 ;
        RECT 1762.360 886.420 1762.620 886.680 ;
        RECT 573.720 15.000 573.980 15.260 ;
        RECT 579.240 15.000 579.500 15.260 ;
      LAYER met2 ;
        RECT 1762.350 1818.475 1762.630 1818.845 ;
        RECT 1762.420 886.710 1762.560 1818.475 ;
        RECT 579.240 886.390 579.500 886.710 ;
        RECT 1762.360 886.390 1762.620 886.710 ;
        RECT 579.300 15.290 579.440 886.390 ;
        RECT 573.720 14.970 573.980 15.290 ;
        RECT 579.240 14.970 579.500 15.290 ;
        RECT 573.780 2.400 573.920 14.970 ;
        RECT 573.570 -4.800 574.130 2.400 ;
      LAYER via2 ;
        RECT 1762.350 1818.520 1762.630 1818.800 ;
      LAYER met3 ;
        RECT 1755.835 1818.810 1759.835 1818.815 ;
        RECT 1762.325 1818.810 1762.655 1818.825 ;
        RECT 1755.835 1818.510 1762.655 1818.810 ;
        RECT 1755.835 1818.215 1759.835 1818.510 ;
        RECT 1762.325 1818.495 1762.655 1818.510 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 593.010 1312.640 593.330 1312.700 ;
        RECT 995.510 1312.640 995.830 1312.700 ;
        RECT 593.010 1312.500 995.830 1312.640 ;
        RECT 593.010 1312.440 593.330 1312.500 ;
        RECT 995.510 1312.440 995.830 1312.500 ;
      LAYER via ;
        RECT 593.040 1312.440 593.300 1312.700 ;
        RECT 995.540 1312.440 995.800 1312.700 ;
      LAYER met2 ;
        RECT 995.580 1323.135 995.860 1327.135 ;
        RECT 995.600 1312.730 995.740 1323.135 ;
        RECT 593.040 1312.410 593.300 1312.730 ;
        RECT 995.540 1312.410 995.800 1312.730 ;
        RECT 593.100 16.730 593.240 1312.410 ;
        RECT 591.260 16.590 593.240 16.730 ;
        RECT 591.260 2.400 591.400 16.590 ;
        RECT 591.050 -4.800 591.610 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 128.025 16.405 128.195 17.935 ;
      LAYER mcon ;
        RECT 128.025 17.765 128.195 17.935 ;
      LAYER met1 ;
        RECT 1265.990 1317.060 1266.310 1317.120 ;
        RECT 1383.750 1317.060 1384.070 1317.120 ;
        RECT 1265.990 1316.920 1384.070 1317.060 ;
        RECT 1265.990 1316.860 1266.310 1316.920 ;
        RECT 1383.750 1316.860 1384.070 1316.920 ;
        RECT 127.965 17.920 128.255 17.965 ;
        RECT 127.965 17.780 1245.980 17.920 ;
        RECT 127.965 17.735 128.255 17.780 ;
        RECT 1245.840 17.580 1245.980 17.780 ;
        RECT 1265.990 17.580 1266.310 17.640 ;
        RECT 1245.840 17.440 1266.310 17.580 ;
        RECT 1265.990 17.380 1266.310 17.440 ;
        RECT 97.590 16.560 97.910 16.620 ;
        RECT 127.965 16.560 128.255 16.605 ;
        RECT 97.590 16.420 128.255 16.560 ;
        RECT 97.590 16.360 97.910 16.420 ;
        RECT 127.965 16.375 128.255 16.420 ;
      LAYER via ;
        RECT 1266.020 1316.860 1266.280 1317.120 ;
        RECT 1383.780 1316.860 1384.040 1317.120 ;
        RECT 1266.020 17.380 1266.280 17.640 ;
        RECT 97.620 16.360 97.880 16.620 ;
      LAYER met2 ;
        RECT 1383.820 1323.135 1384.100 1327.135 ;
        RECT 1383.840 1317.150 1383.980 1323.135 ;
        RECT 1266.020 1316.830 1266.280 1317.150 ;
        RECT 1383.780 1316.830 1384.040 1317.150 ;
        RECT 1266.080 17.670 1266.220 1316.830 ;
        RECT 1266.020 17.350 1266.280 17.670 ;
        RECT 97.620 16.330 97.880 16.650 ;
        RECT 97.680 2.400 97.820 16.330 ;
        RECT 97.470 -4.800 98.030 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1445.390 1311.280 1445.710 1311.340 ;
        RECT 1475.750 1311.280 1476.070 1311.340 ;
        RECT 1445.390 1311.140 1476.070 1311.280 ;
        RECT 1445.390 1311.080 1445.710 1311.140 ;
        RECT 1475.750 1311.080 1476.070 1311.140 ;
        RECT 609.110 18.600 609.430 18.660 ;
        RECT 1445.390 18.600 1445.710 18.660 ;
        RECT 609.110 18.460 1445.710 18.600 ;
        RECT 609.110 18.400 609.430 18.460 ;
        RECT 1445.390 18.400 1445.710 18.460 ;
      LAYER via ;
        RECT 1445.420 1311.080 1445.680 1311.340 ;
        RECT 1475.780 1311.080 1476.040 1311.340 ;
        RECT 609.140 18.400 609.400 18.660 ;
        RECT 1445.420 18.400 1445.680 18.660 ;
      LAYER met2 ;
        RECT 1475.820 1323.135 1476.100 1327.135 ;
        RECT 1475.840 1311.370 1475.980 1323.135 ;
        RECT 1445.420 1311.050 1445.680 1311.370 ;
        RECT 1475.780 1311.050 1476.040 1311.370 ;
        RECT 1445.480 18.690 1445.620 1311.050 ;
        RECT 609.140 18.370 609.400 18.690 ;
        RECT 1445.420 18.370 1445.680 18.690 ;
        RECT 609.200 2.400 609.340 18.370 ;
        RECT 608.990 -4.800 609.550 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 627.510 2077.300 627.830 2077.360 ;
        RECT 696.970 2077.300 697.290 2077.360 ;
        RECT 627.510 2077.160 697.290 2077.300 ;
        RECT 627.510 2077.100 627.830 2077.160 ;
        RECT 696.970 2077.100 697.290 2077.160 ;
      LAYER via ;
        RECT 627.540 2077.100 627.800 2077.360 ;
        RECT 697.000 2077.100 697.260 2077.360 ;
      LAYER met2 ;
        RECT 696.990 2079.595 697.270 2079.965 ;
        RECT 697.060 2077.390 697.200 2079.595 ;
        RECT 627.540 2077.070 627.800 2077.390 ;
        RECT 697.000 2077.070 697.260 2077.390 ;
        RECT 627.600 17.410 627.740 2077.070 ;
        RECT 627.140 17.270 627.740 17.410 ;
        RECT 627.140 2.400 627.280 17.270 ;
        RECT 626.930 -4.800 627.490 2.400 ;
      LAYER via2 ;
        RECT 696.990 2079.640 697.270 2079.920 ;
      LAYER met3 ;
        RECT 696.965 2079.930 697.295 2079.945 ;
        RECT 715.810 2079.930 719.810 2079.935 ;
        RECT 696.965 2079.630 719.810 2079.930 ;
        RECT 696.965 2079.615 697.295 2079.630 ;
        RECT 715.810 2079.335 719.810 2079.630 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 127.490 2393.160 127.810 2393.220 ;
        RECT 1027.710 2393.160 1028.030 2393.220 ;
        RECT 127.490 2393.020 1028.030 2393.160 ;
        RECT 127.490 2392.960 127.810 2393.020 ;
        RECT 1027.710 2392.960 1028.030 2393.020 ;
        RECT 121.510 17.920 121.830 17.980 ;
        RECT 127.490 17.920 127.810 17.980 ;
        RECT 121.510 17.780 127.810 17.920 ;
        RECT 121.510 17.720 121.830 17.780 ;
        RECT 127.490 17.720 127.810 17.780 ;
      LAYER via ;
        RECT 127.520 2392.960 127.780 2393.220 ;
        RECT 1027.740 2392.960 1028.000 2393.220 ;
        RECT 121.540 17.720 121.800 17.980 ;
        RECT 127.520 17.720 127.780 17.980 ;
      LAYER met2 ;
        RECT 127.520 2392.930 127.780 2393.250 ;
        RECT 1027.740 2392.930 1028.000 2393.250 ;
        RECT 127.580 18.010 127.720 2392.930 ;
        RECT 1027.800 2377.880 1027.940 2392.930 ;
        RECT 1027.780 2373.880 1028.060 2377.880 ;
        RECT 121.540 17.690 121.800 18.010 ;
        RECT 127.520 17.690 127.780 18.010 ;
        RECT 121.600 2.400 121.740 17.690 ;
        RECT 121.390 -4.800 121.950 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 150.950 1315.700 151.270 1315.760 ;
        RECT 897.070 1315.700 897.390 1315.760 ;
        RECT 150.950 1315.560 897.390 1315.700 ;
        RECT 150.950 1315.500 151.270 1315.560 ;
        RECT 897.070 1315.500 897.390 1315.560 ;
        RECT 145.430 17.240 145.750 17.300 ;
        RECT 150.950 17.240 151.270 17.300 ;
        RECT 145.430 17.100 151.270 17.240 ;
        RECT 145.430 17.040 145.750 17.100 ;
        RECT 150.950 17.040 151.270 17.100 ;
      LAYER via ;
        RECT 150.980 1315.500 151.240 1315.760 ;
        RECT 897.100 1315.500 897.360 1315.760 ;
        RECT 145.460 17.040 145.720 17.300 ;
        RECT 150.980 17.040 151.240 17.300 ;
      LAYER met2 ;
        RECT 897.140 1323.135 897.420 1327.135 ;
        RECT 897.160 1315.790 897.300 1323.135 ;
        RECT 150.980 1315.470 151.240 1315.790 ;
        RECT 897.100 1315.470 897.360 1315.790 ;
        RECT 151.040 17.330 151.180 1315.470 ;
        RECT 145.460 17.010 145.720 17.330 ;
        RECT 150.980 17.010 151.240 17.330 ;
        RECT 145.520 2.400 145.660 17.010 ;
        RECT 145.310 -4.800 145.870 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 165.210 2104.840 165.530 2104.900 ;
        RECT 709.390 2104.840 709.710 2104.900 ;
        RECT 165.210 2104.700 709.710 2104.840 ;
        RECT 165.210 2104.640 165.530 2104.700 ;
        RECT 709.390 2104.640 709.710 2104.700 ;
      LAYER via ;
        RECT 165.240 2104.640 165.500 2104.900 ;
        RECT 709.420 2104.640 709.680 2104.900 ;
      LAYER met2 ;
        RECT 709.410 2105.435 709.690 2105.805 ;
        RECT 709.480 2104.930 709.620 2105.435 ;
        RECT 165.240 2104.610 165.500 2104.930 ;
        RECT 709.420 2104.610 709.680 2104.930 ;
        RECT 165.300 16.900 165.440 2104.610 ;
        RECT 163.460 16.760 165.440 16.900 ;
        RECT 163.460 2.400 163.600 16.760 ;
        RECT 163.250 -4.800 163.810 2.400 ;
      LAYER via2 ;
        RECT 709.410 2105.480 709.690 2105.760 ;
      LAYER met3 ;
        RECT 709.385 2105.770 709.715 2105.785 ;
        RECT 715.810 2105.770 719.810 2105.775 ;
        RECT 709.385 2105.470 719.810 2105.770 ;
        RECT 709.385 2105.455 709.715 2105.470 ;
        RECT 715.810 2105.175 719.810 2105.470 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1763.270 2211.515 1763.550 2211.885 ;
        RECT 1763.340 1346.245 1763.480 2211.515 ;
        RECT 1763.270 1345.875 1763.550 1346.245 ;
        RECT 180.870 37.555 181.150 37.925 ;
        RECT 180.940 2.400 181.080 37.555 ;
        RECT 180.730 -4.800 181.290 2.400 ;
      LAYER via2 ;
        RECT 1763.270 2211.560 1763.550 2211.840 ;
        RECT 1763.270 1345.920 1763.550 1346.200 ;
        RECT 180.870 37.600 181.150 37.880 ;
      LAYER met3 ;
        RECT 1755.835 2211.850 1759.835 2211.855 ;
        RECT 1763.245 2211.850 1763.575 2211.865 ;
        RECT 1755.835 2211.550 1763.575 2211.850 ;
        RECT 1755.835 2211.255 1759.835 2211.550 ;
        RECT 1763.245 2211.535 1763.575 2211.550 ;
        RECT 1763.245 1346.210 1763.575 1346.225 ;
        RECT 1763.910 1346.210 1764.290 1346.220 ;
        RECT 1763.245 1345.910 1764.290 1346.210 ;
        RECT 1763.245 1345.895 1763.575 1345.910 ;
        RECT 1763.910 1345.900 1764.290 1345.910 ;
        RECT 180.845 37.890 181.175 37.905 ;
        RECT 1763.910 37.890 1764.290 37.900 ;
        RECT 180.845 37.590 1764.290 37.890 ;
        RECT 180.845 37.575 181.175 37.590 ;
        RECT 1763.910 37.580 1764.290 37.590 ;
      LAYER via3 ;
        RECT 1763.940 1345.900 1764.260 1346.220 ;
        RECT 1763.940 37.580 1764.260 37.900 ;
      LAYER met4 ;
        RECT 1763.935 1345.895 1764.265 1346.225 ;
        RECT 1763.950 37.905 1764.250 1345.895 ;
        RECT 1763.935 37.575 1764.265 37.905 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 224.090 2393.500 224.410 2393.560 ;
        RECT 1108.670 2393.500 1108.990 2393.560 ;
        RECT 224.090 2393.360 1108.990 2393.500 ;
        RECT 224.090 2393.300 224.410 2393.360 ;
        RECT 1108.670 2393.300 1108.990 2393.360 ;
        RECT 198.790 14.520 199.110 14.580 ;
        RECT 224.090 14.520 224.410 14.580 ;
        RECT 198.790 14.380 224.410 14.520 ;
        RECT 198.790 14.320 199.110 14.380 ;
        RECT 224.090 14.320 224.410 14.380 ;
      LAYER via ;
        RECT 224.120 2393.300 224.380 2393.560 ;
        RECT 1108.700 2393.300 1108.960 2393.560 ;
        RECT 198.820 14.320 199.080 14.580 ;
        RECT 224.120 14.320 224.380 14.580 ;
      LAYER met2 ;
        RECT 224.120 2393.270 224.380 2393.590 ;
        RECT 1108.700 2393.270 1108.960 2393.590 ;
        RECT 224.180 14.610 224.320 2393.270 ;
        RECT 1108.760 2377.880 1108.900 2393.270 ;
        RECT 1108.740 2373.880 1109.020 2377.880 ;
        RECT 198.820 14.290 199.080 14.610 ;
        RECT 224.120 14.290 224.380 14.610 ;
        RECT 198.880 2.400 199.020 14.290 ;
        RECT 198.670 -4.800 199.230 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 220.410 1312.980 220.730 1313.040 ;
        RECT 741.590 1312.980 741.910 1313.040 ;
        RECT 220.410 1312.840 741.910 1312.980 ;
        RECT 220.410 1312.780 220.730 1312.840 ;
        RECT 741.590 1312.780 741.910 1312.840 ;
        RECT 216.730 15.200 217.050 15.260 ;
        RECT 220.410 15.200 220.730 15.260 ;
        RECT 216.730 15.060 220.730 15.200 ;
        RECT 216.730 15.000 217.050 15.060 ;
        RECT 220.410 15.000 220.730 15.060 ;
      LAYER via ;
        RECT 220.440 1312.780 220.700 1313.040 ;
        RECT 741.620 1312.780 741.880 1313.040 ;
        RECT 216.760 15.000 217.020 15.260 ;
        RECT 220.440 15.000 220.700 15.260 ;
      LAYER met2 ;
        RECT 741.660 1323.135 741.940 1327.135 ;
        RECT 741.680 1313.070 741.820 1323.135 ;
        RECT 220.440 1312.750 220.700 1313.070 ;
        RECT 741.620 1312.750 741.880 1313.070 ;
        RECT 220.500 15.290 220.640 1312.750 ;
        RECT 216.760 14.970 217.020 15.290 ;
        RECT 220.440 14.970 220.700 15.290 ;
        RECT 216.820 2.400 216.960 14.970 ;
        RECT 216.610 -4.800 217.170 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 241.110 1552.680 241.430 1552.740 ;
        RECT 710.310 1552.680 710.630 1552.740 ;
        RECT 241.110 1552.540 710.630 1552.680 ;
        RECT 241.110 1552.480 241.430 1552.540 ;
        RECT 710.310 1552.480 710.630 1552.540 ;
        RECT 234.670 15.880 234.990 15.940 ;
        RECT 241.110 15.880 241.430 15.940 ;
        RECT 234.670 15.740 241.430 15.880 ;
        RECT 234.670 15.680 234.990 15.740 ;
        RECT 241.110 15.680 241.430 15.740 ;
      LAYER via ;
        RECT 241.140 1552.480 241.400 1552.740 ;
        RECT 710.340 1552.480 710.600 1552.740 ;
        RECT 234.700 15.680 234.960 15.940 ;
        RECT 241.140 15.680 241.400 15.940 ;
      LAYER met2 ;
        RECT 710.330 1557.355 710.610 1557.725 ;
        RECT 710.400 1552.770 710.540 1557.355 ;
        RECT 241.140 1552.450 241.400 1552.770 ;
        RECT 710.340 1552.450 710.600 1552.770 ;
        RECT 241.200 15.970 241.340 1552.450 ;
        RECT 234.700 15.650 234.960 15.970 ;
        RECT 241.140 15.650 241.400 15.970 ;
        RECT 234.760 2.400 234.900 15.650 ;
        RECT 234.550 -4.800 235.110 2.400 ;
      LAYER via2 ;
        RECT 710.330 1557.400 710.610 1557.680 ;
      LAYER met3 ;
        RECT 710.305 1557.690 710.635 1557.705 ;
        RECT 715.810 1557.690 719.810 1557.695 ;
        RECT 710.305 1557.390 719.810 1557.690 ;
        RECT 710.305 1557.375 710.635 1557.390 ;
        RECT 715.810 1557.095 719.810 1557.390 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 793.570 2389.420 793.890 2389.480 ;
        RECT 783.540 2389.280 793.890 2389.420 ;
        RECT 86.090 2389.080 86.410 2389.140 ;
        RECT 783.540 2389.080 783.680 2389.280 ;
        RECT 793.570 2389.220 793.890 2389.280 ;
        RECT 86.090 2388.940 783.680 2389.080 ;
        RECT 86.090 2388.880 86.410 2388.940 ;
        RECT 56.190 15.200 56.510 15.260 ;
        RECT 85.170 15.200 85.490 15.260 ;
        RECT 56.190 15.060 85.490 15.200 ;
        RECT 56.190 15.000 56.510 15.060 ;
        RECT 85.170 15.000 85.490 15.060 ;
      LAYER via ;
        RECT 86.120 2388.880 86.380 2389.140 ;
        RECT 793.600 2389.220 793.860 2389.480 ;
        RECT 56.220 15.000 56.480 15.260 ;
        RECT 85.200 15.000 85.460 15.260 ;
      LAYER met2 ;
        RECT 793.600 2389.190 793.860 2389.510 ;
        RECT 86.120 2388.850 86.380 2389.170 ;
        RECT 86.180 18.770 86.320 2388.850 ;
        RECT 793.660 2377.010 793.800 2389.190 ;
        RECT 796.860 2377.010 797.140 2377.880 ;
        RECT 793.660 2376.870 797.140 2377.010 ;
        RECT 796.860 2373.880 797.140 2376.870 ;
        RECT 85.260 18.630 86.320 18.770 ;
        RECT 85.260 15.290 85.400 18.630 ;
        RECT 56.220 14.970 56.480 15.290 ;
        RECT 85.200 14.970 85.460 15.290 ;
        RECT 56.280 2.400 56.420 14.970 ;
        RECT 56.070 -4.800 56.630 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 80.110 18.260 80.430 18.320 ;
        RECT 99.890 18.260 100.210 18.320 ;
        RECT 80.110 18.120 100.210 18.260 ;
        RECT 80.110 18.060 80.430 18.120 ;
        RECT 99.890 18.060 100.210 18.120 ;
      LAYER via ;
        RECT 80.140 18.060 80.400 18.320 ;
        RECT 99.920 18.060 100.180 18.320 ;
      LAYER met2 ;
        RECT 99.910 2387.635 100.190 2388.005 ;
        RECT 1045.210 2387.635 1045.490 2388.005 ;
        RECT 99.980 18.350 100.120 2387.635 ;
        RECT 1045.280 2377.880 1045.420 2387.635 ;
        RECT 1045.260 2373.880 1045.540 2377.880 ;
        RECT 80.140 18.030 80.400 18.350 ;
        RECT 99.920 18.030 100.180 18.350 ;
        RECT 80.200 2.400 80.340 18.030 ;
        RECT 79.990 -4.800 80.550 2.400 ;
      LAYER via2 ;
        RECT 99.910 2387.680 100.190 2387.960 ;
        RECT 1045.210 2387.680 1045.490 2387.960 ;
      LAYER met3 ;
        RECT 99.885 2387.970 100.215 2387.985 ;
        RECT 1045.185 2387.970 1045.515 2387.985 ;
        RECT 99.885 2387.670 1045.515 2387.970 ;
        RECT 99.885 2387.655 100.215 2387.670 ;
        RECT 1045.185 2387.655 1045.515 2387.670 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 690.145 2380.765 690.315 2384.335 ;
        RECT 727.865 2380.765 728.035 2384.335 ;
      LAYER mcon ;
        RECT 690.145 2384.165 690.315 2384.335 ;
        RECT 727.865 2384.165 728.035 2384.335 ;
      LAYER met1 ;
        RECT 690.085 2384.320 690.375 2384.365 ;
        RECT 727.805 2384.320 728.095 2384.365 ;
        RECT 690.085 2384.180 728.095 2384.320 ;
        RECT 690.085 2384.135 690.375 2384.180 ;
        RECT 727.805 2384.135 728.095 2384.180 ;
        RECT 110.010 2380.920 110.330 2380.980 ;
        RECT 690.085 2380.920 690.375 2380.965 ;
        RECT 110.010 2380.780 690.375 2380.920 ;
        RECT 110.010 2380.720 110.330 2380.780 ;
        RECT 690.085 2380.735 690.375 2380.780 ;
        RECT 727.805 2380.920 728.095 2380.965 ;
        RECT 1519.910 2380.920 1520.230 2380.980 ;
        RECT 727.805 2380.780 1520.230 2380.920 ;
        RECT 727.805 2380.735 728.095 2380.780 ;
        RECT 1519.910 2380.720 1520.230 2380.780 ;
        RECT 103.570 17.920 103.890 17.980 ;
        RECT 110.010 17.920 110.330 17.980 ;
        RECT 103.570 17.780 110.330 17.920 ;
        RECT 103.570 17.720 103.890 17.780 ;
        RECT 110.010 17.720 110.330 17.780 ;
      LAYER via ;
        RECT 110.040 2380.720 110.300 2380.980 ;
        RECT 1519.940 2380.720 1520.200 2380.980 ;
        RECT 103.600 17.720 103.860 17.980 ;
        RECT 110.040 17.720 110.300 17.980 ;
      LAYER met2 ;
        RECT 110.040 2380.690 110.300 2381.010 ;
        RECT 1519.940 2380.690 1520.200 2381.010 ;
        RECT 110.100 18.010 110.240 2380.690 ;
        RECT 1520.000 2377.880 1520.140 2380.690 ;
        RECT 1519.980 2373.880 1520.260 2377.880 ;
        RECT 103.600 17.690 103.860 18.010 ;
        RECT 110.040 17.690 110.300 18.010 ;
        RECT 103.660 2.400 103.800 17.690 ;
        RECT 103.450 -4.800 104.010 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 127.490 16.900 127.810 16.960 ;
        RECT 130.710 16.900 131.030 16.960 ;
        RECT 127.490 16.760 131.030 16.900 ;
        RECT 127.490 16.700 127.810 16.760 ;
        RECT 130.710 16.700 131.030 16.760 ;
      LAYER via ;
        RECT 127.520 16.700 127.780 16.960 ;
        RECT 130.740 16.700 131.000 16.960 ;
      LAYER met2 ;
        RECT 821.260 2376.190 823.240 2376.330 ;
        RECT 821.260 2375.765 821.400 2376.190 ;
        RECT 823.100 2375.765 823.240 2376.190 ;
        RECT 130.730 2375.395 131.010 2375.765 ;
        RECT 821.190 2375.395 821.470 2375.765 ;
        RECT 823.030 2375.395 823.310 2375.765 ;
        RECT 1380.090 2375.650 1380.370 2375.765 ;
        RECT 1381.060 2375.650 1381.340 2377.880 ;
        RECT 1380.090 2375.510 1381.340 2375.650 ;
        RECT 1380.090 2375.395 1380.370 2375.510 ;
        RECT 130.800 16.990 130.940 2375.395 ;
        RECT 1381.060 2373.880 1381.340 2375.510 ;
        RECT 127.520 16.670 127.780 16.990 ;
        RECT 130.740 16.670 131.000 16.990 ;
        RECT 127.580 2.400 127.720 16.670 ;
        RECT 127.370 -4.800 127.930 2.400 ;
      LAYER via2 ;
        RECT 130.730 2375.440 131.010 2375.720 ;
        RECT 821.190 2375.440 821.470 2375.720 ;
        RECT 823.030 2375.440 823.310 2375.720 ;
        RECT 1380.090 2375.440 1380.370 2375.720 ;
      LAYER met3 ;
        RECT 130.705 2375.730 131.035 2375.745 ;
        RECT 821.165 2375.730 821.495 2375.745 ;
        RECT 130.705 2375.430 821.495 2375.730 ;
        RECT 130.705 2375.415 131.035 2375.430 ;
        RECT 821.165 2375.415 821.495 2375.430 ;
        RECT 823.005 2375.730 823.335 2375.745 ;
        RECT 1380.065 2375.730 1380.395 2375.745 ;
        RECT 823.005 2375.430 1380.395 2375.730 ;
        RECT 823.005 2375.415 823.335 2375.430 ;
        RECT 1380.065 2375.415 1380.395 2375.430 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 155.090 2388.400 155.410 2388.460 ;
        RECT 911.790 2388.400 912.110 2388.460 ;
        RECT 155.090 2388.260 912.110 2388.400 ;
        RECT 155.090 2388.200 155.410 2388.260 ;
        RECT 911.790 2388.200 912.110 2388.260 ;
        RECT 26.290 17.240 26.610 17.300 ;
        RECT 26.290 17.100 133.240 17.240 ;
        RECT 26.290 17.040 26.610 17.100 ;
        RECT 133.100 16.900 133.240 17.100 ;
        RECT 155.090 16.900 155.410 16.960 ;
        RECT 133.100 16.760 155.410 16.900 ;
        RECT 155.090 16.700 155.410 16.760 ;
      LAYER via ;
        RECT 155.120 2388.200 155.380 2388.460 ;
        RECT 911.820 2388.200 912.080 2388.460 ;
        RECT 26.320 17.040 26.580 17.300 ;
        RECT 155.120 16.700 155.380 16.960 ;
      LAYER met2 ;
        RECT 155.120 2388.170 155.380 2388.490 ;
        RECT 911.820 2388.170 912.080 2388.490 ;
        RECT 26.320 17.010 26.580 17.330 ;
        RECT 26.380 2.400 26.520 17.010 ;
        RECT 155.180 16.990 155.320 2388.170 ;
        RECT 911.880 2377.880 912.020 2388.170 ;
        RECT 911.860 2373.880 912.140 2377.880 ;
        RECT 155.120 16.670 155.380 16.990 ;
        RECT 26.170 -4.800 26.730 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1245.365 16.065 1245.535 17.595 ;
      LAYER mcon ;
        RECT 1245.365 17.425 1245.535 17.595 ;
      LAYER met1 ;
        RECT 1286.690 1313.660 1287.010 1313.720 ;
        RECT 1325.790 1313.660 1326.110 1313.720 ;
        RECT 1286.690 1313.520 1326.110 1313.660 ;
        RECT 1286.690 1313.460 1287.010 1313.520 ;
        RECT 1325.790 1313.460 1326.110 1313.520 ;
        RECT 32.270 17.580 32.590 17.640 ;
        RECT 1245.305 17.580 1245.595 17.625 ;
        RECT 32.270 17.440 1245.595 17.580 ;
        RECT 32.270 17.380 32.590 17.440 ;
        RECT 1245.305 17.395 1245.595 17.440 ;
        RECT 1245.305 16.220 1245.595 16.265 ;
        RECT 1286.690 16.220 1287.010 16.280 ;
        RECT 1245.305 16.080 1287.010 16.220 ;
        RECT 1245.305 16.035 1245.595 16.080 ;
        RECT 1286.690 16.020 1287.010 16.080 ;
      LAYER via ;
        RECT 1286.720 1313.460 1286.980 1313.720 ;
        RECT 1325.820 1313.460 1326.080 1313.720 ;
        RECT 32.300 17.380 32.560 17.640 ;
        RECT 1286.720 16.020 1286.980 16.280 ;
      LAYER met2 ;
        RECT 1325.860 1323.135 1326.140 1327.135 ;
        RECT 1325.880 1313.750 1326.020 1323.135 ;
        RECT 1286.720 1313.430 1286.980 1313.750 ;
        RECT 1325.820 1313.430 1326.080 1313.750 ;
        RECT 32.300 17.350 32.560 17.670 ;
        RECT 32.360 2.400 32.500 17.350 ;
        RECT 1286.780 16.310 1286.920 1313.430 ;
        RECT 1286.720 15.990 1286.980 16.310 ;
        RECT 32.150 -4.800 32.710 2.400 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INOUT ;
    PORT
      LAYER met4 ;
        RECT 2704.020 3517.600 2707.020 3529.000 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    PORT
      LAYER met4 ;
        RECT 2931.300 -9.320 2934.300 3529.000 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    PORT
      LAYER met4 ;
        RECT 2902.020 3517.600 2905.020 3538.400 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    PORT
      LAYER met4 ;
        RECT 2940.700 -18.720 2943.700 3538.400 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    PORT
      LAYER met4 ;
        RECT 2740.020 3517.600 2743.020 3547.800 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    PORT
      LAYER met4 ;
        RECT 2950.100 -28.120 2953.100 3547.800 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    PORT
      LAYER met4 ;
        RECT 2758.020 3517.600 2761.020 3557.200 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    PORT
      LAYER met4 ;
        RECT 2959.500 -37.520 2962.500 3557.200 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 721.330 1333.930 1754.030 2364.980 ;
      LAYER met1 ;
        RECT 721.330 1333.775 1754.030 2373.695 ;
      LAYER met2 ;
        RECT 721.980 2373.600 726.660 2373.880 ;
        RECT 727.500 2373.600 733.100 2373.880 ;
        RECT 733.940 2373.600 738.620 2373.880 ;
        RECT 739.460 2373.600 744.140 2373.880 ;
        RECT 744.980 2373.600 749.660 2373.880 ;
        RECT 750.500 2373.600 756.100 2373.880 ;
        RECT 756.940 2373.600 761.620 2373.880 ;
        RECT 762.460 2373.600 767.140 2373.880 ;
        RECT 767.980 2373.600 773.580 2373.880 ;
        RECT 774.420 2373.600 779.100 2373.880 ;
        RECT 779.940 2373.600 784.620 2373.880 ;
        RECT 785.460 2373.600 790.140 2373.880 ;
        RECT 790.980 2373.600 796.580 2373.880 ;
        RECT 797.420 2373.600 802.100 2373.880 ;
        RECT 802.940 2373.600 807.620 2373.880 ;
        RECT 808.460 2373.600 814.060 2373.880 ;
        RECT 814.900 2373.600 819.580 2373.880 ;
        RECT 820.420 2373.600 825.100 2373.880 ;
        RECT 825.940 2373.600 830.620 2373.880 ;
        RECT 831.460 2373.600 837.060 2373.880 ;
        RECT 837.900 2373.600 842.580 2373.880 ;
        RECT 843.420 2373.600 848.100 2373.880 ;
        RECT 848.940 2373.600 854.540 2373.880 ;
        RECT 855.380 2373.600 860.060 2373.880 ;
        RECT 860.900 2373.600 865.580 2373.880 ;
        RECT 866.420 2373.600 871.100 2373.880 ;
        RECT 871.940 2373.600 877.540 2373.880 ;
        RECT 878.380 2373.600 883.060 2373.880 ;
        RECT 883.900 2373.600 888.580 2373.880 ;
        RECT 889.420 2373.600 895.020 2373.880 ;
        RECT 895.860 2373.600 900.540 2373.880 ;
        RECT 901.380 2373.600 906.060 2373.880 ;
        RECT 906.900 2373.600 911.580 2373.880 ;
        RECT 912.420 2373.600 918.020 2373.880 ;
        RECT 918.860 2373.600 923.540 2373.880 ;
        RECT 924.380 2373.600 929.060 2373.880 ;
        RECT 929.900 2373.600 935.500 2373.880 ;
        RECT 936.340 2373.600 941.020 2373.880 ;
        RECT 941.860 2373.600 946.540 2373.880 ;
        RECT 947.380 2373.600 952.060 2373.880 ;
        RECT 952.900 2373.600 958.500 2373.880 ;
        RECT 959.340 2373.600 964.020 2373.880 ;
        RECT 964.860 2373.600 969.540 2373.880 ;
        RECT 970.380 2373.600 975.980 2373.880 ;
        RECT 976.820 2373.600 981.500 2373.880 ;
        RECT 982.340 2373.600 987.020 2373.880 ;
        RECT 987.860 2373.600 992.540 2373.880 ;
        RECT 993.380 2373.600 998.980 2373.880 ;
        RECT 999.820 2373.600 1004.500 2373.880 ;
        RECT 1005.340 2373.600 1010.020 2373.880 ;
        RECT 1010.860 2373.600 1016.460 2373.880 ;
        RECT 1017.300 2373.600 1021.980 2373.880 ;
        RECT 1022.820 2373.600 1027.500 2373.880 ;
        RECT 1028.340 2373.600 1033.020 2373.880 ;
        RECT 1033.860 2373.600 1039.460 2373.880 ;
        RECT 1040.300 2373.600 1044.980 2373.880 ;
        RECT 1045.820 2373.600 1050.500 2373.880 ;
        RECT 1051.340 2373.600 1056.940 2373.880 ;
        RECT 1057.780 2373.600 1062.460 2373.880 ;
        RECT 1063.300 2373.600 1067.980 2373.880 ;
        RECT 1068.820 2373.600 1074.420 2373.880 ;
        RECT 1075.260 2373.600 1079.940 2373.880 ;
        RECT 1080.780 2373.600 1085.460 2373.880 ;
        RECT 1086.300 2373.600 1090.980 2373.880 ;
        RECT 1091.820 2373.600 1097.420 2373.880 ;
        RECT 1098.260 2373.600 1102.940 2373.880 ;
        RECT 1103.780 2373.600 1108.460 2373.880 ;
        RECT 1109.300 2373.600 1114.900 2373.880 ;
        RECT 1115.740 2373.600 1120.420 2373.880 ;
        RECT 1121.260 2373.600 1125.940 2373.880 ;
        RECT 1126.780 2373.600 1131.460 2373.880 ;
        RECT 1132.300 2373.600 1137.900 2373.880 ;
        RECT 1138.740 2373.600 1143.420 2373.880 ;
        RECT 1144.260 2373.600 1148.940 2373.880 ;
        RECT 1149.780 2373.600 1155.380 2373.880 ;
        RECT 1156.220 2373.600 1160.900 2373.880 ;
        RECT 1161.740 2373.600 1166.420 2373.880 ;
        RECT 1167.260 2373.600 1171.940 2373.880 ;
        RECT 1172.780 2373.600 1178.380 2373.880 ;
        RECT 1179.220 2373.600 1183.900 2373.880 ;
        RECT 1184.740 2373.600 1189.420 2373.880 ;
        RECT 1190.260 2373.600 1195.860 2373.880 ;
        RECT 1196.700 2373.600 1201.380 2373.880 ;
        RECT 1202.220 2373.600 1206.900 2373.880 ;
        RECT 1207.740 2373.600 1212.420 2373.880 ;
        RECT 1213.260 2373.600 1218.860 2373.880 ;
        RECT 1219.700 2373.600 1224.380 2373.880 ;
        RECT 1225.220 2373.600 1229.900 2373.880 ;
        RECT 1230.740 2373.600 1236.340 2373.880 ;
        RECT 1237.180 2373.600 1241.860 2373.880 ;
        RECT 1242.700 2373.600 1247.380 2373.880 ;
        RECT 1248.220 2373.600 1252.900 2373.880 ;
        RECT 1253.740 2373.600 1259.340 2373.880 ;
        RECT 1260.180 2373.600 1264.860 2373.880 ;
        RECT 1265.700 2373.600 1270.380 2373.880 ;
        RECT 1271.220 2373.600 1276.820 2373.880 ;
        RECT 1277.660 2373.600 1282.340 2373.880 ;
        RECT 1283.180 2373.600 1287.860 2373.880 ;
        RECT 1288.700 2373.600 1293.380 2373.880 ;
        RECT 1294.220 2373.600 1299.820 2373.880 ;
        RECT 1300.660 2373.600 1305.340 2373.880 ;
        RECT 1306.180 2373.600 1310.860 2373.880 ;
        RECT 1311.700 2373.600 1317.300 2373.880 ;
        RECT 1318.140 2373.600 1322.820 2373.880 ;
        RECT 1323.660 2373.600 1328.340 2373.880 ;
        RECT 1329.180 2373.600 1333.860 2373.880 ;
        RECT 1334.700 2373.600 1340.300 2373.880 ;
        RECT 1341.140 2373.600 1345.820 2373.880 ;
        RECT 1346.660 2373.600 1351.340 2373.880 ;
        RECT 1352.180 2373.600 1357.780 2373.880 ;
        RECT 1358.620 2373.600 1363.300 2373.880 ;
        RECT 1364.140 2373.600 1368.820 2373.880 ;
        RECT 1369.660 2373.600 1374.340 2373.880 ;
        RECT 1375.180 2373.600 1380.780 2373.880 ;
        RECT 1381.620 2373.600 1386.300 2373.880 ;
        RECT 1387.140 2373.600 1391.820 2373.880 ;
        RECT 1392.660 2373.600 1398.260 2373.880 ;
        RECT 1399.100 2373.600 1403.780 2373.880 ;
        RECT 1404.620 2373.600 1409.300 2373.880 ;
        RECT 1410.140 2373.600 1415.740 2373.880 ;
        RECT 1416.580 2373.600 1421.260 2373.880 ;
        RECT 1422.100 2373.600 1426.780 2373.880 ;
        RECT 1427.620 2373.600 1432.300 2373.880 ;
        RECT 1433.140 2373.600 1438.740 2373.880 ;
        RECT 1439.580 2373.600 1444.260 2373.880 ;
        RECT 1445.100 2373.600 1449.780 2373.880 ;
        RECT 1450.620 2373.600 1456.220 2373.880 ;
        RECT 1457.060 2373.600 1461.740 2373.880 ;
        RECT 1462.580 2373.600 1467.260 2373.880 ;
        RECT 1468.100 2373.600 1472.780 2373.880 ;
        RECT 1473.620 2373.600 1479.220 2373.880 ;
        RECT 1480.060 2373.600 1484.740 2373.880 ;
        RECT 1485.580 2373.600 1490.260 2373.880 ;
        RECT 1491.100 2373.600 1496.700 2373.880 ;
        RECT 1497.540 2373.600 1502.220 2373.880 ;
        RECT 1503.060 2373.600 1507.740 2373.880 ;
        RECT 1508.580 2373.600 1513.260 2373.880 ;
        RECT 1514.100 2373.600 1519.700 2373.880 ;
        RECT 1520.540 2373.600 1525.220 2373.880 ;
        RECT 1526.060 2373.600 1530.740 2373.880 ;
        RECT 1531.580 2373.600 1537.180 2373.880 ;
        RECT 1538.020 2373.600 1542.700 2373.880 ;
        RECT 1543.540 2373.600 1548.220 2373.880 ;
        RECT 1549.060 2373.600 1553.740 2373.880 ;
        RECT 1554.580 2373.600 1560.180 2373.880 ;
        RECT 1561.020 2373.600 1565.700 2373.880 ;
        RECT 1566.540 2373.600 1571.220 2373.880 ;
        RECT 1572.060 2373.600 1577.660 2373.880 ;
        RECT 1578.500 2373.600 1583.180 2373.880 ;
        RECT 1584.020 2373.600 1588.700 2373.880 ;
        RECT 1589.540 2373.600 1594.220 2373.880 ;
        RECT 1595.060 2373.600 1600.660 2373.880 ;
        RECT 1601.500 2373.600 1606.180 2373.880 ;
        RECT 1607.020 2373.600 1611.700 2373.880 ;
        RECT 1612.540 2373.600 1618.140 2373.880 ;
        RECT 1618.980 2373.600 1623.660 2373.880 ;
        RECT 1624.500 2373.600 1629.180 2373.880 ;
        RECT 1630.020 2373.600 1634.700 2373.880 ;
        RECT 1635.540 2373.600 1641.140 2373.880 ;
        RECT 1641.980 2373.600 1646.660 2373.880 ;
        RECT 1647.500 2373.600 1652.180 2373.880 ;
        RECT 1653.020 2373.600 1658.620 2373.880 ;
        RECT 1659.460 2373.600 1664.140 2373.880 ;
        RECT 1664.980 2373.600 1669.660 2373.880 ;
        RECT 1670.500 2373.600 1675.180 2373.880 ;
        RECT 1676.020 2373.600 1681.620 2373.880 ;
        RECT 1682.460 2373.600 1687.140 2373.880 ;
        RECT 1687.980 2373.600 1692.660 2373.880 ;
        RECT 1693.500 2373.600 1699.100 2373.880 ;
        RECT 1699.940 2373.600 1704.620 2373.880 ;
        RECT 1705.460 2373.600 1710.140 2373.880 ;
        RECT 1710.980 2373.600 1715.660 2373.880 ;
        RECT 1716.500 2373.600 1722.100 2373.880 ;
        RECT 1722.940 2373.600 1727.620 2373.880 ;
        RECT 1728.460 2373.600 1733.140 2373.880 ;
        RECT 1733.980 2373.600 1739.580 2373.880 ;
        RECT 1740.420 2373.600 1745.100 2373.880 ;
        RECT 1745.940 2373.600 1750.620 2373.880 ;
        RECT 721.430 1327.415 1751.170 2373.600 ;
        RECT 721.430 1327.135 723.900 1327.415 ;
        RECT 724.740 1327.135 729.420 1327.415 ;
        RECT 730.260 1327.135 734.940 1327.415 ;
        RECT 735.780 1327.135 741.380 1327.415 ;
        RECT 742.220 1327.135 746.900 1327.415 ;
        RECT 747.740 1327.135 752.420 1327.415 ;
        RECT 753.260 1327.135 758.860 1327.415 ;
        RECT 759.700 1327.135 764.380 1327.415 ;
        RECT 765.220 1327.135 769.900 1327.415 ;
        RECT 770.740 1327.135 775.420 1327.415 ;
        RECT 776.260 1327.135 781.860 1327.415 ;
        RECT 782.700 1327.135 787.380 1327.415 ;
        RECT 788.220 1327.135 792.900 1327.415 ;
        RECT 793.740 1327.135 799.340 1327.415 ;
        RECT 800.180 1327.135 804.860 1327.415 ;
        RECT 805.700 1327.135 810.380 1327.415 ;
        RECT 811.220 1327.135 815.900 1327.415 ;
        RECT 816.740 1327.135 822.340 1327.415 ;
        RECT 823.180 1327.135 827.860 1327.415 ;
        RECT 828.700 1327.135 833.380 1327.415 ;
        RECT 834.220 1327.135 839.820 1327.415 ;
        RECT 840.660 1327.135 845.340 1327.415 ;
        RECT 846.180 1327.135 850.860 1327.415 ;
        RECT 851.700 1327.135 856.380 1327.415 ;
        RECT 857.220 1327.135 862.820 1327.415 ;
        RECT 863.660 1327.135 868.340 1327.415 ;
        RECT 869.180 1327.135 873.860 1327.415 ;
        RECT 874.700 1327.135 880.300 1327.415 ;
        RECT 881.140 1327.135 885.820 1327.415 ;
        RECT 886.660 1327.135 891.340 1327.415 ;
        RECT 892.180 1327.135 896.860 1327.415 ;
        RECT 897.700 1327.135 903.300 1327.415 ;
        RECT 904.140 1327.135 908.820 1327.415 ;
        RECT 909.660 1327.135 914.340 1327.415 ;
        RECT 915.180 1327.135 920.780 1327.415 ;
        RECT 921.620 1327.135 926.300 1327.415 ;
        RECT 927.140 1327.135 931.820 1327.415 ;
        RECT 932.660 1327.135 937.340 1327.415 ;
        RECT 938.180 1327.135 943.780 1327.415 ;
        RECT 944.620 1327.135 949.300 1327.415 ;
        RECT 950.140 1327.135 954.820 1327.415 ;
        RECT 955.660 1327.135 961.260 1327.415 ;
        RECT 962.100 1327.135 966.780 1327.415 ;
        RECT 967.620 1327.135 972.300 1327.415 ;
        RECT 973.140 1327.135 977.820 1327.415 ;
        RECT 978.660 1327.135 984.260 1327.415 ;
        RECT 985.100 1327.135 989.780 1327.415 ;
        RECT 990.620 1327.135 995.300 1327.415 ;
        RECT 996.140 1327.135 1001.740 1327.415 ;
        RECT 1002.580 1327.135 1007.260 1327.415 ;
        RECT 1008.100 1327.135 1012.780 1327.415 ;
        RECT 1013.620 1327.135 1018.300 1327.415 ;
        RECT 1019.140 1327.135 1024.740 1327.415 ;
        RECT 1025.580 1327.135 1030.260 1327.415 ;
        RECT 1031.100 1327.135 1035.780 1327.415 ;
        RECT 1036.620 1327.135 1042.220 1327.415 ;
        RECT 1043.060 1327.135 1047.740 1327.415 ;
        RECT 1048.580 1327.135 1053.260 1327.415 ;
        RECT 1054.100 1327.135 1058.780 1327.415 ;
        RECT 1059.620 1327.135 1065.220 1327.415 ;
        RECT 1066.060 1327.135 1070.740 1327.415 ;
        RECT 1071.580 1327.135 1076.260 1327.415 ;
        RECT 1077.100 1327.135 1082.700 1327.415 ;
        RECT 1083.540 1327.135 1088.220 1327.415 ;
        RECT 1089.060 1327.135 1093.740 1327.415 ;
        RECT 1094.580 1327.135 1100.180 1327.415 ;
        RECT 1101.020 1327.135 1105.700 1327.415 ;
        RECT 1106.540 1327.135 1111.220 1327.415 ;
        RECT 1112.060 1327.135 1116.740 1327.415 ;
        RECT 1117.580 1327.135 1123.180 1327.415 ;
        RECT 1124.020 1327.135 1128.700 1327.415 ;
        RECT 1129.540 1327.135 1134.220 1327.415 ;
        RECT 1135.060 1327.135 1140.660 1327.415 ;
        RECT 1141.500 1327.135 1146.180 1327.415 ;
        RECT 1147.020 1327.135 1151.700 1327.415 ;
        RECT 1152.540 1327.135 1157.220 1327.415 ;
        RECT 1158.060 1327.135 1163.660 1327.415 ;
        RECT 1164.500 1327.135 1169.180 1327.415 ;
        RECT 1170.020 1327.135 1174.700 1327.415 ;
        RECT 1175.540 1327.135 1181.140 1327.415 ;
        RECT 1181.980 1327.135 1186.660 1327.415 ;
        RECT 1187.500 1327.135 1192.180 1327.415 ;
        RECT 1193.020 1327.135 1197.700 1327.415 ;
        RECT 1198.540 1327.135 1204.140 1327.415 ;
        RECT 1204.980 1327.135 1209.660 1327.415 ;
        RECT 1210.500 1327.135 1215.180 1327.415 ;
        RECT 1216.020 1327.135 1221.620 1327.415 ;
        RECT 1222.460 1327.135 1227.140 1327.415 ;
        RECT 1227.980 1327.135 1232.660 1327.415 ;
        RECT 1233.500 1327.135 1238.180 1327.415 ;
        RECT 1239.020 1327.135 1244.620 1327.415 ;
        RECT 1245.460 1327.135 1250.140 1327.415 ;
        RECT 1250.980 1327.135 1255.660 1327.415 ;
        RECT 1256.500 1327.135 1262.100 1327.415 ;
        RECT 1262.940 1327.135 1267.620 1327.415 ;
        RECT 1268.460 1327.135 1273.140 1327.415 ;
        RECT 1273.980 1327.135 1278.660 1327.415 ;
        RECT 1279.500 1327.135 1285.100 1327.415 ;
        RECT 1285.940 1327.135 1290.620 1327.415 ;
        RECT 1291.460 1327.135 1296.140 1327.415 ;
        RECT 1296.980 1327.135 1302.580 1327.415 ;
        RECT 1303.420 1327.135 1308.100 1327.415 ;
        RECT 1308.940 1327.135 1313.620 1327.415 ;
        RECT 1314.460 1327.135 1319.140 1327.415 ;
        RECT 1319.980 1327.135 1325.580 1327.415 ;
        RECT 1326.420 1327.135 1331.100 1327.415 ;
        RECT 1331.940 1327.135 1336.620 1327.415 ;
        RECT 1337.460 1327.135 1343.060 1327.415 ;
        RECT 1343.900 1327.135 1348.580 1327.415 ;
        RECT 1349.420 1327.135 1354.100 1327.415 ;
        RECT 1354.940 1327.135 1359.620 1327.415 ;
        RECT 1360.460 1327.135 1366.060 1327.415 ;
        RECT 1366.900 1327.135 1371.580 1327.415 ;
        RECT 1372.420 1327.135 1377.100 1327.415 ;
        RECT 1377.940 1327.135 1383.540 1327.415 ;
        RECT 1384.380 1327.135 1389.060 1327.415 ;
        RECT 1389.900 1327.135 1394.580 1327.415 ;
        RECT 1395.420 1327.135 1400.100 1327.415 ;
        RECT 1400.940 1327.135 1406.540 1327.415 ;
        RECT 1407.380 1327.135 1412.060 1327.415 ;
        RECT 1412.900 1327.135 1417.580 1327.415 ;
        RECT 1418.420 1327.135 1424.020 1327.415 ;
        RECT 1424.860 1327.135 1429.540 1327.415 ;
        RECT 1430.380 1327.135 1435.060 1327.415 ;
        RECT 1435.900 1327.135 1441.500 1327.415 ;
        RECT 1442.340 1327.135 1447.020 1327.415 ;
        RECT 1447.860 1327.135 1452.540 1327.415 ;
        RECT 1453.380 1327.135 1458.060 1327.415 ;
        RECT 1458.900 1327.135 1464.500 1327.415 ;
        RECT 1465.340 1327.135 1470.020 1327.415 ;
        RECT 1470.860 1327.135 1475.540 1327.415 ;
        RECT 1476.380 1327.135 1481.980 1327.415 ;
        RECT 1482.820 1327.135 1487.500 1327.415 ;
        RECT 1488.340 1327.135 1493.020 1327.415 ;
        RECT 1493.860 1327.135 1498.540 1327.415 ;
        RECT 1499.380 1327.135 1504.980 1327.415 ;
        RECT 1505.820 1327.135 1510.500 1327.415 ;
        RECT 1511.340 1327.135 1516.020 1327.415 ;
        RECT 1516.860 1327.135 1522.460 1327.415 ;
        RECT 1523.300 1327.135 1527.980 1327.415 ;
        RECT 1528.820 1327.135 1533.500 1327.415 ;
        RECT 1534.340 1327.135 1539.020 1327.415 ;
        RECT 1539.860 1327.135 1545.460 1327.415 ;
        RECT 1546.300 1327.135 1550.980 1327.415 ;
        RECT 1551.820 1327.135 1556.500 1327.415 ;
        RECT 1557.340 1327.135 1562.940 1327.415 ;
        RECT 1563.780 1327.135 1568.460 1327.415 ;
        RECT 1569.300 1327.135 1573.980 1327.415 ;
        RECT 1574.820 1327.135 1579.500 1327.415 ;
        RECT 1580.340 1327.135 1585.940 1327.415 ;
        RECT 1586.780 1327.135 1591.460 1327.415 ;
        RECT 1592.300 1327.135 1596.980 1327.415 ;
        RECT 1597.820 1327.135 1603.420 1327.415 ;
        RECT 1604.260 1327.135 1608.940 1327.415 ;
        RECT 1609.780 1327.135 1614.460 1327.415 ;
        RECT 1615.300 1327.135 1619.980 1327.415 ;
        RECT 1620.820 1327.135 1626.420 1327.415 ;
        RECT 1627.260 1327.135 1631.940 1327.415 ;
        RECT 1632.780 1327.135 1637.460 1327.415 ;
        RECT 1638.300 1327.135 1643.900 1327.415 ;
        RECT 1644.740 1327.135 1649.420 1327.415 ;
        RECT 1650.260 1327.135 1654.940 1327.415 ;
        RECT 1655.780 1327.135 1660.460 1327.415 ;
        RECT 1661.300 1327.135 1666.900 1327.415 ;
        RECT 1667.740 1327.135 1672.420 1327.415 ;
        RECT 1673.260 1327.135 1677.940 1327.415 ;
        RECT 1678.780 1327.135 1684.380 1327.415 ;
        RECT 1685.220 1327.135 1689.900 1327.415 ;
        RECT 1690.740 1327.135 1695.420 1327.415 ;
        RECT 1696.260 1327.135 1700.940 1327.415 ;
        RECT 1701.780 1327.135 1707.380 1327.415 ;
        RECT 1708.220 1327.135 1712.900 1327.415 ;
        RECT 1713.740 1327.135 1718.420 1327.415 ;
        RECT 1719.260 1327.135 1724.860 1327.415 ;
        RECT 1725.700 1327.135 1730.380 1327.415 ;
        RECT 1731.220 1327.135 1735.900 1327.415 ;
        RECT 1736.740 1327.135 1741.420 1327.415 ;
        RECT 1742.260 1327.135 1747.860 1327.415 ;
        RECT 1748.700 1327.135 1751.170 1327.415 ;
      LAYER met3 ;
        RECT 719.810 2364.535 1755.435 2365.060 ;
        RECT 719.810 2361.855 1755.835 2364.535 ;
        RECT 720.210 2360.455 1755.835 2361.855 ;
        RECT 719.810 2357.775 1755.835 2360.455 ;
        RECT 719.810 2356.375 1755.435 2357.775 ;
        RECT 719.810 2353.695 1755.835 2356.375 ;
        RECT 720.210 2352.295 1755.835 2353.695 ;
        RECT 719.810 2349.615 1755.835 2352.295 ;
        RECT 719.810 2348.215 1755.435 2349.615 ;
        RECT 719.810 2345.535 1755.835 2348.215 ;
        RECT 720.210 2344.135 1755.835 2345.535 ;
        RECT 719.810 2340.095 1755.835 2344.135 ;
        RECT 719.810 2338.695 1755.435 2340.095 ;
        RECT 719.810 2336.015 1755.835 2338.695 ;
        RECT 720.210 2334.615 1755.835 2336.015 ;
        RECT 719.810 2331.935 1755.835 2334.615 ;
        RECT 719.810 2330.535 1755.435 2331.935 ;
        RECT 719.810 2327.855 1755.835 2330.535 ;
        RECT 720.210 2326.455 1755.835 2327.855 ;
        RECT 719.810 2323.775 1755.835 2326.455 ;
        RECT 719.810 2322.375 1755.435 2323.775 ;
        RECT 719.810 2319.695 1755.835 2322.375 ;
        RECT 720.210 2318.295 1755.835 2319.695 ;
        RECT 719.810 2314.255 1755.835 2318.295 ;
        RECT 719.810 2312.855 1755.435 2314.255 ;
        RECT 719.810 2311.535 1755.835 2312.855 ;
        RECT 720.210 2310.135 1755.835 2311.535 ;
        RECT 719.810 2306.095 1755.835 2310.135 ;
        RECT 719.810 2304.695 1755.435 2306.095 ;
        RECT 719.810 2302.015 1755.835 2304.695 ;
        RECT 720.210 2300.615 1755.835 2302.015 ;
        RECT 719.810 2297.935 1755.835 2300.615 ;
        RECT 719.810 2296.535 1755.435 2297.935 ;
        RECT 719.810 2293.855 1755.835 2296.535 ;
        RECT 720.210 2292.455 1755.835 2293.855 ;
        RECT 719.810 2289.775 1755.835 2292.455 ;
        RECT 719.810 2288.375 1755.435 2289.775 ;
        RECT 719.810 2285.695 1755.835 2288.375 ;
        RECT 720.210 2284.295 1755.835 2285.695 ;
        RECT 719.810 2280.255 1755.835 2284.295 ;
        RECT 719.810 2278.855 1755.435 2280.255 ;
        RECT 719.810 2276.175 1755.835 2278.855 ;
        RECT 720.210 2274.775 1755.835 2276.175 ;
        RECT 719.810 2272.095 1755.835 2274.775 ;
        RECT 719.810 2270.695 1755.435 2272.095 ;
        RECT 719.810 2268.015 1755.835 2270.695 ;
        RECT 720.210 2266.615 1755.835 2268.015 ;
        RECT 719.810 2263.935 1755.835 2266.615 ;
        RECT 719.810 2262.535 1755.435 2263.935 ;
        RECT 719.810 2259.855 1755.835 2262.535 ;
        RECT 720.210 2258.455 1755.835 2259.855 ;
        RECT 719.810 2254.415 1755.835 2258.455 ;
        RECT 719.810 2253.015 1755.435 2254.415 ;
        RECT 719.810 2251.695 1755.835 2253.015 ;
        RECT 720.210 2250.295 1755.835 2251.695 ;
        RECT 719.810 2246.255 1755.835 2250.295 ;
        RECT 719.810 2244.855 1755.435 2246.255 ;
        RECT 719.810 2242.175 1755.835 2244.855 ;
        RECT 720.210 2240.775 1755.835 2242.175 ;
        RECT 719.810 2238.095 1755.835 2240.775 ;
        RECT 719.810 2236.695 1755.435 2238.095 ;
        RECT 719.810 2234.015 1755.835 2236.695 ;
        RECT 720.210 2232.615 1755.835 2234.015 ;
        RECT 719.810 2229.935 1755.835 2232.615 ;
        RECT 719.810 2228.535 1755.435 2229.935 ;
        RECT 719.810 2225.855 1755.835 2228.535 ;
        RECT 720.210 2224.455 1755.835 2225.855 ;
        RECT 719.810 2220.415 1755.835 2224.455 ;
        RECT 719.810 2219.015 1755.435 2220.415 ;
        RECT 719.810 2216.335 1755.835 2219.015 ;
        RECT 720.210 2214.935 1755.835 2216.335 ;
        RECT 719.810 2212.255 1755.835 2214.935 ;
        RECT 719.810 2210.855 1755.435 2212.255 ;
        RECT 719.810 2208.175 1755.835 2210.855 ;
        RECT 720.210 2206.775 1755.835 2208.175 ;
        RECT 719.810 2204.095 1755.835 2206.775 ;
        RECT 719.810 2202.695 1755.435 2204.095 ;
        RECT 719.810 2200.015 1755.835 2202.695 ;
        RECT 720.210 2198.615 1755.835 2200.015 ;
        RECT 719.810 2194.575 1755.835 2198.615 ;
        RECT 719.810 2193.175 1755.435 2194.575 ;
        RECT 719.810 2191.855 1755.835 2193.175 ;
        RECT 720.210 2190.455 1755.835 2191.855 ;
        RECT 719.810 2186.415 1755.835 2190.455 ;
        RECT 719.810 2185.015 1755.435 2186.415 ;
        RECT 719.810 2182.335 1755.835 2185.015 ;
        RECT 720.210 2180.935 1755.835 2182.335 ;
        RECT 719.810 2178.255 1755.835 2180.935 ;
        RECT 719.810 2176.855 1755.435 2178.255 ;
        RECT 719.810 2174.175 1755.835 2176.855 ;
        RECT 720.210 2172.775 1755.835 2174.175 ;
        RECT 719.810 2170.095 1755.835 2172.775 ;
        RECT 719.810 2168.695 1755.435 2170.095 ;
        RECT 719.810 2166.015 1755.835 2168.695 ;
        RECT 720.210 2164.615 1755.835 2166.015 ;
        RECT 719.810 2160.575 1755.835 2164.615 ;
        RECT 719.810 2159.175 1755.435 2160.575 ;
        RECT 719.810 2156.495 1755.835 2159.175 ;
        RECT 720.210 2155.095 1755.835 2156.495 ;
        RECT 719.810 2152.415 1755.835 2155.095 ;
        RECT 719.810 2151.015 1755.435 2152.415 ;
        RECT 719.810 2148.335 1755.835 2151.015 ;
        RECT 720.210 2146.935 1755.835 2148.335 ;
        RECT 719.810 2144.255 1755.835 2146.935 ;
        RECT 719.810 2142.855 1755.435 2144.255 ;
        RECT 719.810 2140.175 1755.835 2142.855 ;
        RECT 720.210 2138.775 1755.835 2140.175 ;
        RECT 719.810 2134.735 1755.835 2138.775 ;
        RECT 719.810 2133.335 1755.435 2134.735 ;
        RECT 719.810 2132.015 1755.835 2133.335 ;
        RECT 720.210 2130.615 1755.835 2132.015 ;
        RECT 719.810 2126.575 1755.835 2130.615 ;
        RECT 719.810 2125.175 1755.435 2126.575 ;
        RECT 719.810 2122.495 1755.835 2125.175 ;
        RECT 720.210 2121.095 1755.835 2122.495 ;
        RECT 719.810 2118.415 1755.835 2121.095 ;
        RECT 719.810 2117.015 1755.435 2118.415 ;
        RECT 719.810 2114.335 1755.835 2117.015 ;
        RECT 720.210 2112.935 1755.835 2114.335 ;
        RECT 719.810 2110.255 1755.835 2112.935 ;
        RECT 719.810 2108.855 1755.435 2110.255 ;
        RECT 719.810 2106.175 1755.835 2108.855 ;
        RECT 720.210 2104.775 1755.835 2106.175 ;
        RECT 719.810 2100.735 1755.835 2104.775 ;
        RECT 719.810 2099.335 1755.435 2100.735 ;
        RECT 719.810 2096.655 1755.835 2099.335 ;
        RECT 720.210 2095.255 1755.835 2096.655 ;
        RECT 719.810 2092.575 1755.835 2095.255 ;
        RECT 719.810 2091.175 1755.435 2092.575 ;
        RECT 719.810 2088.495 1755.835 2091.175 ;
        RECT 720.210 2087.095 1755.835 2088.495 ;
        RECT 719.810 2084.415 1755.835 2087.095 ;
        RECT 719.810 2083.015 1755.435 2084.415 ;
        RECT 719.810 2080.335 1755.835 2083.015 ;
        RECT 720.210 2078.935 1755.835 2080.335 ;
        RECT 719.810 2074.895 1755.835 2078.935 ;
        RECT 719.810 2073.495 1755.435 2074.895 ;
        RECT 719.810 2072.175 1755.835 2073.495 ;
        RECT 720.210 2070.775 1755.835 2072.175 ;
        RECT 719.810 2066.735 1755.835 2070.775 ;
        RECT 719.810 2065.335 1755.435 2066.735 ;
        RECT 719.810 2062.655 1755.835 2065.335 ;
        RECT 720.210 2061.255 1755.835 2062.655 ;
        RECT 719.810 2058.575 1755.835 2061.255 ;
        RECT 719.810 2057.175 1755.435 2058.575 ;
        RECT 719.810 2054.495 1755.835 2057.175 ;
        RECT 720.210 2053.095 1755.835 2054.495 ;
        RECT 719.810 2050.415 1755.835 2053.095 ;
        RECT 719.810 2049.015 1755.435 2050.415 ;
        RECT 719.810 2046.335 1755.835 2049.015 ;
        RECT 720.210 2044.935 1755.835 2046.335 ;
        RECT 719.810 2040.895 1755.835 2044.935 ;
        RECT 719.810 2039.495 1755.435 2040.895 ;
        RECT 719.810 2036.815 1755.835 2039.495 ;
        RECT 720.210 2035.415 1755.835 2036.815 ;
        RECT 719.810 2032.735 1755.835 2035.415 ;
        RECT 719.810 2031.335 1755.435 2032.735 ;
        RECT 719.810 2028.655 1755.835 2031.335 ;
        RECT 720.210 2027.255 1755.835 2028.655 ;
        RECT 719.810 2024.575 1755.835 2027.255 ;
        RECT 719.810 2023.175 1755.435 2024.575 ;
        RECT 719.810 2020.495 1755.835 2023.175 ;
        RECT 720.210 2019.095 1755.835 2020.495 ;
        RECT 719.810 2015.055 1755.835 2019.095 ;
        RECT 719.810 2013.655 1755.435 2015.055 ;
        RECT 719.810 2012.335 1755.835 2013.655 ;
        RECT 720.210 2010.935 1755.835 2012.335 ;
        RECT 719.810 2006.895 1755.835 2010.935 ;
        RECT 719.810 2005.495 1755.435 2006.895 ;
        RECT 719.810 2002.815 1755.835 2005.495 ;
        RECT 720.210 2001.415 1755.835 2002.815 ;
        RECT 719.810 1998.735 1755.835 2001.415 ;
        RECT 719.810 1997.335 1755.435 1998.735 ;
        RECT 719.810 1994.655 1755.835 1997.335 ;
        RECT 720.210 1993.255 1755.835 1994.655 ;
        RECT 719.810 1990.575 1755.835 1993.255 ;
        RECT 719.810 1989.175 1755.435 1990.575 ;
        RECT 719.810 1986.495 1755.835 1989.175 ;
        RECT 720.210 1985.095 1755.835 1986.495 ;
        RECT 719.810 1981.055 1755.835 1985.095 ;
        RECT 719.810 1979.655 1755.435 1981.055 ;
        RECT 719.810 1976.975 1755.835 1979.655 ;
        RECT 720.210 1975.575 1755.835 1976.975 ;
        RECT 719.810 1972.895 1755.835 1975.575 ;
        RECT 719.810 1971.495 1755.435 1972.895 ;
        RECT 719.810 1968.815 1755.835 1971.495 ;
        RECT 720.210 1967.415 1755.835 1968.815 ;
        RECT 719.810 1964.735 1755.835 1967.415 ;
        RECT 719.810 1963.335 1755.435 1964.735 ;
        RECT 719.810 1960.655 1755.835 1963.335 ;
        RECT 720.210 1959.255 1755.835 1960.655 ;
        RECT 719.810 1955.215 1755.835 1959.255 ;
        RECT 719.810 1953.815 1755.435 1955.215 ;
        RECT 719.810 1952.495 1755.835 1953.815 ;
        RECT 720.210 1951.095 1755.835 1952.495 ;
        RECT 719.810 1947.055 1755.835 1951.095 ;
        RECT 719.810 1945.655 1755.435 1947.055 ;
        RECT 719.810 1942.975 1755.835 1945.655 ;
        RECT 720.210 1941.575 1755.835 1942.975 ;
        RECT 719.810 1938.895 1755.835 1941.575 ;
        RECT 719.810 1937.495 1755.435 1938.895 ;
        RECT 719.810 1934.815 1755.835 1937.495 ;
        RECT 720.210 1933.415 1755.835 1934.815 ;
        RECT 719.810 1930.735 1755.835 1933.415 ;
        RECT 719.810 1929.335 1755.435 1930.735 ;
        RECT 719.810 1926.655 1755.835 1929.335 ;
        RECT 720.210 1925.255 1755.835 1926.655 ;
        RECT 719.810 1921.215 1755.835 1925.255 ;
        RECT 719.810 1919.815 1755.435 1921.215 ;
        RECT 719.810 1917.135 1755.835 1919.815 ;
        RECT 720.210 1915.735 1755.835 1917.135 ;
        RECT 719.810 1913.055 1755.835 1915.735 ;
        RECT 719.810 1911.655 1755.435 1913.055 ;
        RECT 719.810 1908.975 1755.835 1911.655 ;
        RECT 720.210 1907.575 1755.835 1908.975 ;
        RECT 719.810 1904.895 1755.835 1907.575 ;
        RECT 719.810 1903.495 1755.435 1904.895 ;
        RECT 719.810 1900.815 1755.835 1903.495 ;
        RECT 720.210 1899.415 1755.835 1900.815 ;
        RECT 719.810 1895.375 1755.835 1899.415 ;
        RECT 719.810 1893.975 1755.435 1895.375 ;
        RECT 719.810 1892.655 1755.835 1893.975 ;
        RECT 720.210 1891.255 1755.835 1892.655 ;
        RECT 719.810 1887.215 1755.835 1891.255 ;
        RECT 719.810 1885.815 1755.435 1887.215 ;
        RECT 719.810 1883.135 1755.835 1885.815 ;
        RECT 720.210 1881.735 1755.835 1883.135 ;
        RECT 719.810 1879.055 1755.835 1881.735 ;
        RECT 719.810 1877.655 1755.435 1879.055 ;
        RECT 719.810 1874.975 1755.835 1877.655 ;
        RECT 720.210 1873.575 1755.835 1874.975 ;
        RECT 719.810 1870.895 1755.835 1873.575 ;
        RECT 719.810 1869.495 1755.435 1870.895 ;
        RECT 719.810 1866.815 1755.835 1869.495 ;
        RECT 720.210 1865.415 1755.835 1866.815 ;
        RECT 719.810 1861.375 1755.835 1865.415 ;
        RECT 719.810 1859.975 1755.435 1861.375 ;
        RECT 719.810 1857.295 1755.835 1859.975 ;
        RECT 720.210 1855.895 1755.835 1857.295 ;
        RECT 719.810 1853.215 1755.835 1855.895 ;
        RECT 719.810 1851.815 1755.435 1853.215 ;
        RECT 719.810 1849.135 1755.835 1851.815 ;
        RECT 720.210 1847.735 1755.835 1849.135 ;
        RECT 719.810 1845.055 1755.835 1847.735 ;
        RECT 719.810 1843.655 1755.435 1845.055 ;
        RECT 719.810 1840.975 1755.835 1843.655 ;
        RECT 720.210 1839.575 1755.835 1840.975 ;
        RECT 719.810 1835.535 1755.835 1839.575 ;
        RECT 719.810 1834.135 1755.435 1835.535 ;
        RECT 719.810 1831.455 1755.835 1834.135 ;
        RECT 720.210 1830.055 1755.835 1831.455 ;
        RECT 719.810 1827.375 1755.835 1830.055 ;
        RECT 719.810 1825.975 1755.435 1827.375 ;
        RECT 719.810 1823.295 1755.835 1825.975 ;
        RECT 720.210 1821.895 1755.835 1823.295 ;
        RECT 719.810 1819.215 1755.835 1821.895 ;
        RECT 719.810 1817.815 1755.435 1819.215 ;
        RECT 719.810 1815.135 1755.835 1817.815 ;
        RECT 720.210 1813.735 1755.835 1815.135 ;
        RECT 719.810 1809.695 1755.835 1813.735 ;
        RECT 719.810 1808.295 1755.435 1809.695 ;
        RECT 719.810 1806.975 1755.835 1808.295 ;
        RECT 720.210 1805.575 1755.835 1806.975 ;
        RECT 719.810 1801.535 1755.835 1805.575 ;
        RECT 719.810 1800.135 1755.435 1801.535 ;
        RECT 719.810 1797.455 1755.835 1800.135 ;
        RECT 720.210 1796.055 1755.835 1797.455 ;
        RECT 719.810 1793.375 1755.835 1796.055 ;
        RECT 719.810 1791.975 1755.435 1793.375 ;
        RECT 719.810 1789.295 1755.835 1791.975 ;
        RECT 720.210 1787.895 1755.835 1789.295 ;
        RECT 719.810 1785.215 1755.835 1787.895 ;
        RECT 719.810 1783.815 1755.435 1785.215 ;
        RECT 719.810 1781.135 1755.835 1783.815 ;
        RECT 720.210 1779.735 1755.835 1781.135 ;
        RECT 719.810 1775.695 1755.835 1779.735 ;
        RECT 719.810 1774.295 1755.435 1775.695 ;
        RECT 719.810 1771.615 1755.835 1774.295 ;
        RECT 720.210 1770.215 1755.835 1771.615 ;
        RECT 719.810 1767.535 1755.835 1770.215 ;
        RECT 719.810 1766.135 1755.435 1767.535 ;
        RECT 719.810 1763.455 1755.835 1766.135 ;
        RECT 720.210 1762.055 1755.835 1763.455 ;
        RECT 719.810 1759.375 1755.835 1762.055 ;
        RECT 719.810 1757.975 1755.435 1759.375 ;
        RECT 719.810 1755.295 1755.835 1757.975 ;
        RECT 720.210 1753.895 1755.835 1755.295 ;
        RECT 719.810 1749.855 1755.835 1753.895 ;
        RECT 719.810 1748.455 1755.435 1749.855 ;
        RECT 719.810 1747.135 1755.835 1748.455 ;
        RECT 720.210 1745.735 1755.835 1747.135 ;
        RECT 719.810 1741.695 1755.835 1745.735 ;
        RECT 719.810 1740.295 1755.435 1741.695 ;
        RECT 719.810 1737.615 1755.835 1740.295 ;
        RECT 720.210 1736.215 1755.835 1737.615 ;
        RECT 719.810 1733.535 1755.835 1736.215 ;
        RECT 719.810 1732.135 1755.435 1733.535 ;
        RECT 719.810 1729.455 1755.835 1732.135 ;
        RECT 720.210 1728.055 1755.835 1729.455 ;
        RECT 719.810 1725.375 1755.835 1728.055 ;
        RECT 719.810 1723.975 1755.435 1725.375 ;
        RECT 719.810 1721.295 1755.835 1723.975 ;
        RECT 720.210 1719.895 1755.835 1721.295 ;
        RECT 719.810 1715.855 1755.835 1719.895 ;
        RECT 719.810 1714.455 1755.435 1715.855 ;
        RECT 719.810 1711.775 1755.835 1714.455 ;
        RECT 720.210 1710.375 1755.835 1711.775 ;
        RECT 719.810 1707.695 1755.835 1710.375 ;
        RECT 719.810 1706.295 1755.435 1707.695 ;
        RECT 719.810 1703.615 1755.835 1706.295 ;
        RECT 720.210 1702.215 1755.835 1703.615 ;
        RECT 719.810 1699.535 1755.835 1702.215 ;
        RECT 719.810 1698.135 1755.435 1699.535 ;
        RECT 719.810 1695.455 1755.835 1698.135 ;
        RECT 720.210 1694.055 1755.835 1695.455 ;
        RECT 719.810 1690.015 1755.835 1694.055 ;
        RECT 719.810 1688.615 1755.435 1690.015 ;
        RECT 719.810 1687.295 1755.835 1688.615 ;
        RECT 720.210 1685.895 1755.835 1687.295 ;
        RECT 719.810 1681.855 1755.835 1685.895 ;
        RECT 719.810 1680.455 1755.435 1681.855 ;
        RECT 719.810 1677.775 1755.835 1680.455 ;
        RECT 720.210 1676.375 1755.835 1677.775 ;
        RECT 719.810 1673.695 1755.835 1676.375 ;
        RECT 719.810 1672.295 1755.435 1673.695 ;
        RECT 719.810 1669.615 1755.835 1672.295 ;
        RECT 720.210 1668.215 1755.835 1669.615 ;
        RECT 719.810 1665.535 1755.835 1668.215 ;
        RECT 719.810 1664.135 1755.435 1665.535 ;
        RECT 719.810 1661.455 1755.835 1664.135 ;
        RECT 720.210 1660.055 1755.835 1661.455 ;
        RECT 719.810 1656.015 1755.835 1660.055 ;
        RECT 719.810 1654.615 1755.435 1656.015 ;
        RECT 719.810 1651.935 1755.835 1654.615 ;
        RECT 720.210 1650.535 1755.835 1651.935 ;
        RECT 719.810 1647.855 1755.835 1650.535 ;
        RECT 719.810 1646.455 1755.435 1647.855 ;
        RECT 719.810 1643.775 1755.835 1646.455 ;
        RECT 720.210 1642.375 1755.835 1643.775 ;
        RECT 719.810 1639.695 1755.835 1642.375 ;
        RECT 719.810 1638.295 1755.435 1639.695 ;
        RECT 719.810 1635.615 1755.835 1638.295 ;
        RECT 720.210 1634.215 1755.835 1635.615 ;
        RECT 719.810 1630.175 1755.835 1634.215 ;
        RECT 719.810 1628.775 1755.435 1630.175 ;
        RECT 719.810 1627.455 1755.835 1628.775 ;
        RECT 720.210 1626.055 1755.835 1627.455 ;
        RECT 719.810 1622.015 1755.835 1626.055 ;
        RECT 719.810 1620.615 1755.435 1622.015 ;
        RECT 719.810 1617.935 1755.835 1620.615 ;
        RECT 720.210 1616.535 1755.835 1617.935 ;
        RECT 719.810 1613.855 1755.835 1616.535 ;
        RECT 719.810 1612.455 1755.435 1613.855 ;
        RECT 719.810 1609.775 1755.835 1612.455 ;
        RECT 720.210 1608.375 1755.835 1609.775 ;
        RECT 719.810 1605.695 1755.835 1608.375 ;
        RECT 719.810 1604.295 1755.435 1605.695 ;
        RECT 719.810 1601.615 1755.835 1604.295 ;
        RECT 720.210 1600.215 1755.835 1601.615 ;
        RECT 719.810 1596.175 1755.835 1600.215 ;
        RECT 719.810 1594.775 1755.435 1596.175 ;
        RECT 719.810 1592.095 1755.835 1594.775 ;
        RECT 720.210 1590.695 1755.835 1592.095 ;
        RECT 719.810 1588.015 1755.835 1590.695 ;
        RECT 719.810 1586.615 1755.435 1588.015 ;
        RECT 719.810 1583.935 1755.835 1586.615 ;
        RECT 720.210 1582.535 1755.835 1583.935 ;
        RECT 719.810 1579.855 1755.835 1582.535 ;
        RECT 719.810 1578.455 1755.435 1579.855 ;
        RECT 719.810 1575.775 1755.835 1578.455 ;
        RECT 720.210 1574.375 1755.835 1575.775 ;
        RECT 719.810 1570.335 1755.835 1574.375 ;
        RECT 719.810 1568.935 1755.435 1570.335 ;
        RECT 719.810 1567.615 1755.835 1568.935 ;
        RECT 720.210 1566.215 1755.835 1567.615 ;
        RECT 719.810 1562.175 1755.835 1566.215 ;
        RECT 719.810 1560.775 1755.435 1562.175 ;
        RECT 719.810 1558.095 1755.835 1560.775 ;
        RECT 720.210 1556.695 1755.835 1558.095 ;
        RECT 719.810 1554.015 1755.835 1556.695 ;
        RECT 719.810 1552.615 1755.435 1554.015 ;
        RECT 719.810 1549.935 1755.835 1552.615 ;
        RECT 720.210 1548.535 1755.835 1549.935 ;
        RECT 719.810 1545.855 1755.835 1548.535 ;
        RECT 719.810 1544.455 1755.435 1545.855 ;
        RECT 719.810 1541.775 1755.835 1544.455 ;
        RECT 720.210 1540.375 1755.835 1541.775 ;
        RECT 719.810 1536.335 1755.835 1540.375 ;
        RECT 719.810 1534.935 1755.435 1536.335 ;
        RECT 719.810 1532.255 1755.835 1534.935 ;
        RECT 720.210 1530.855 1755.835 1532.255 ;
        RECT 719.810 1528.175 1755.835 1530.855 ;
        RECT 719.810 1526.775 1755.435 1528.175 ;
        RECT 719.810 1524.095 1755.835 1526.775 ;
        RECT 720.210 1522.695 1755.835 1524.095 ;
        RECT 719.810 1520.015 1755.835 1522.695 ;
        RECT 719.810 1518.615 1755.435 1520.015 ;
        RECT 719.810 1515.935 1755.835 1518.615 ;
        RECT 720.210 1514.535 1755.835 1515.935 ;
        RECT 719.810 1510.495 1755.835 1514.535 ;
        RECT 719.810 1509.095 1755.435 1510.495 ;
        RECT 719.810 1507.775 1755.835 1509.095 ;
        RECT 720.210 1506.375 1755.835 1507.775 ;
        RECT 719.810 1502.335 1755.835 1506.375 ;
        RECT 719.810 1500.935 1755.435 1502.335 ;
        RECT 719.810 1498.255 1755.835 1500.935 ;
        RECT 720.210 1496.855 1755.835 1498.255 ;
        RECT 719.810 1494.175 1755.835 1496.855 ;
        RECT 719.810 1492.775 1755.435 1494.175 ;
        RECT 719.810 1490.095 1755.835 1492.775 ;
        RECT 720.210 1488.695 1755.835 1490.095 ;
        RECT 719.810 1486.015 1755.835 1488.695 ;
        RECT 719.810 1484.615 1755.435 1486.015 ;
        RECT 719.810 1481.935 1755.835 1484.615 ;
        RECT 720.210 1480.535 1755.835 1481.935 ;
        RECT 719.810 1476.495 1755.835 1480.535 ;
        RECT 719.810 1475.095 1755.435 1476.495 ;
        RECT 719.810 1472.415 1755.835 1475.095 ;
        RECT 720.210 1471.015 1755.835 1472.415 ;
        RECT 719.810 1468.335 1755.835 1471.015 ;
        RECT 719.810 1466.935 1755.435 1468.335 ;
        RECT 719.810 1464.255 1755.835 1466.935 ;
        RECT 720.210 1462.855 1755.835 1464.255 ;
        RECT 719.810 1460.175 1755.835 1462.855 ;
        RECT 719.810 1458.775 1755.435 1460.175 ;
        RECT 719.810 1456.095 1755.835 1458.775 ;
        RECT 720.210 1454.695 1755.835 1456.095 ;
        RECT 719.810 1450.655 1755.835 1454.695 ;
        RECT 719.810 1449.255 1755.435 1450.655 ;
        RECT 719.810 1447.935 1755.835 1449.255 ;
        RECT 720.210 1446.535 1755.835 1447.935 ;
        RECT 719.810 1442.495 1755.835 1446.535 ;
        RECT 719.810 1441.095 1755.435 1442.495 ;
        RECT 719.810 1438.415 1755.835 1441.095 ;
        RECT 720.210 1437.015 1755.835 1438.415 ;
        RECT 719.810 1434.335 1755.835 1437.015 ;
        RECT 719.810 1432.935 1755.435 1434.335 ;
        RECT 719.810 1430.255 1755.835 1432.935 ;
        RECT 720.210 1428.855 1755.835 1430.255 ;
        RECT 719.810 1426.175 1755.835 1428.855 ;
        RECT 719.810 1424.775 1755.435 1426.175 ;
        RECT 719.810 1422.095 1755.835 1424.775 ;
        RECT 720.210 1420.695 1755.835 1422.095 ;
        RECT 719.810 1416.655 1755.835 1420.695 ;
        RECT 719.810 1415.255 1755.435 1416.655 ;
        RECT 719.810 1412.575 1755.835 1415.255 ;
        RECT 720.210 1411.175 1755.835 1412.575 ;
        RECT 719.810 1408.495 1755.835 1411.175 ;
        RECT 719.810 1407.095 1755.435 1408.495 ;
        RECT 719.810 1404.415 1755.835 1407.095 ;
        RECT 720.210 1403.015 1755.835 1404.415 ;
        RECT 719.810 1400.335 1755.835 1403.015 ;
        RECT 719.810 1398.935 1755.435 1400.335 ;
        RECT 719.810 1396.255 1755.835 1398.935 ;
        RECT 720.210 1394.855 1755.835 1396.255 ;
        RECT 719.810 1390.815 1755.835 1394.855 ;
        RECT 719.810 1389.415 1755.435 1390.815 ;
        RECT 719.810 1388.095 1755.835 1389.415 ;
        RECT 720.210 1386.695 1755.835 1388.095 ;
        RECT 719.810 1382.655 1755.835 1386.695 ;
        RECT 719.810 1381.255 1755.435 1382.655 ;
        RECT 719.810 1378.575 1755.835 1381.255 ;
        RECT 720.210 1377.175 1755.835 1378.575 ;
        RECT 719.810 1374.495 1755.835 1377.175 ;
        RECT 719.810 1373.095 1755.435 1374.495 ;
        RECT 719.810 1370.415 1755.835 1373.095 ;
        RECT 720.210 1369.015 1755.835 1370.415 ;
        RECT 719.810 1366.335 1755.835 1369.015 ;
        RECT 719.810 1364.935 1755.435 1366.335 ;
        RECT 719.810 1362.255 1755.835 1364.935 ;
        RECT 720.210 1360.855 1755.835 1362.255 ;
        RECT 719.810 1356.815 1755.835 1360.855 ;
        RECT 719.810 1355.415 1755.435 1356.815 ;
        RECT 719.810 1352.735 1755.835 1355.415 ;
        RECT 720.210 1351.335 1755.835 1352.735 ;
        RECT 719.810 1348.655 1755.835 1351.335 ;
        RECT 719.810 1347.255 1755.435 1348.655 ;
        RECT 719.810 1344.575 1755.835 1347.255 ;
        RECT 720.210 1343.175 1755.835 1344.575 ;
        RECT 719.810 1340.495 1755.835 1343.175 ;
        RECT 719.810 1339.095 1755.435 1340.495 ;
        RECT 719.810 1336.415 1755.835 1339.095 ;
        RECT 720.210 1335.015 1755.835 1336.415 ;
        RECT 719.810 1330.975 1755.835 1335.015 ;
        RECT 719.810 1329.575 1755.435 1330.975 ;
        RECT 719.810 1327.390 1755.835 1329.575 ;
      LAYER met4 ;
        RECT 732.665 1333.775 1742.235 2365.135 ;
      LAYER met5 ;
        RECT 721.330 1502.805 1754.030 2346.895 ;
      LAYER met5 ;
        RECT 721.330 1426.215 1754.030 1427.815 ;
        RECT 721.330 1349.625 1754.030 1351.225 ;
  END
END user_project_wrapper
END LIBRARY

