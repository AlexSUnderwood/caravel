magic
tech sky130A
magscale 1 2
timestamp 1608153117
<< checkpaint >>
rect -1260 -1260 718860 1038860
<< metal1 >>
rect 93904 1010925 93910 1010977
rect 93962 1010965 93968 1010977
rect 97072 1010965 97078 1010977
rect 93962 1010937 97078 1010965
rect 93962 1010925 93968 1010937
rect 97072 1010925 97078 1010937
rect 97130 1010925 97136 1010977
rect 440656 1005671 440662 1005723
rect 440714 1005711 440720 1005723
rect 446608 1005711 446614 1005723
rect 440714 1005683 446614 1005711
rect 440714 1005671 440720 1005683
rect 446608 1005671 446614 1005683
rect 446666 1005671 446672 1005723
rect 115696 1005637 115702 1005649
rect 113602 1005609 115702 1005637
rect 93712 1005523 93718 1005575
rect 93770 1005563 93776 1005575
rect 113602 1005563 113630 1005609
rect 115696 1005597 115702 1005609
rect 115754 1005597 115760 1005649
rect 93770 1005535 113630 1005563
rect 93770 1005523 93776 1005535
rect 439216 1005523 439222 1005575
rect 439274 1005563 439280 1005575
rect 446416 1005563 446422 1005575
rect 439274 1005535 446422 1005563
rect 439274 1005523 439280 1005535
rect 446416 1005523 446422 1005535
rect 446474 1005523 446480 1005575
rect 97072 1005449 97078 1005501
rect 97130 1005489 97136 1005501
rect 118192 1005489 118198 1005501
rect 97130 1005461 118198 1005489
rect 97130 1005449 97136 1005461
rect 118192 1005449 118198 1005461
rect 118250 1005449 118256 1005501
rect 298480 1005449 298486 1005501
rect 298538 1005489 298544 1005501
rect 312784 1005489 312790 1005501
rect 298538 1005461 312790 1005489
rect 298538 1005449 298544 1005461
rect 312784 1005449 312790 1005461
rect 312842 1005449 312848 1005501
rect 365104 1005449 365110 1005501
rect 365162 1005489 365168 1005501
rect 383632 1005489 383638 1005501
rect 365162 1005461 383638 1005489
rect 365162 1005449 365168 1005461
rect 383632 1005449 383638 1005461
rect 383690 1005449 383696 1005501
rect 433168 1005449 433174 1005501
rect 433226 1005489 433232 1005501
rect 460816 1005489 460822 1005501
rect 433226 1005461 460822 1005489
rect 433226 1005449 433232 1005461
rect 460816 1005449 460822 1005461
rect 460874 1005449 460880 1005501
rect 558736 1005449 558742 1005501
rect 558794 1005489 558800 1005501
rect 572848 1005489 572854 1005501
rect 558794 1005461 572854 1005489
rect 558794 1005449 558800 1005461
rect 572848 1005449 572854 1005461
rect 572906 1005449 572912 1005501
rect 92560 1005375 92566 1005427
rect 92618 1005415 92624 1005427
rect 102160 1005415 102166 1005427
rect 92618 1005387 102166 1005415
rect 92618 1005375 92624 1005387
rect 102160 1005375 102166 1005387
rect 102218 1005375 102224 1005427
rect 298384 1005375 298390 1005427
rect 298442 1005415 298448 1005427
rect 313840 1005415 313846 1005427
rect 298442 1005387 313846 1005415
rect 298442 1005375 298448 1005387
rect 313840 1005375 313846 1005387
rect 313898 1005375 313904 1005427
rect 430864 1005375 430870 1005427
rect 430922 1005415 430928 1005427
rect 446032 1005415 446038 1005427
rect 430922 1005387 446038 1005415
rect 430922 1005375 430928 1005387
rect 446032 1005375 446038 1005387
rect 446090 1005375 446096 1005427
rect 446608 1005375 446614 1005427
rect 446666 1005415 446672 1005427
rect 469840 1005415 469846 1005427
rect 446666 1005387 469846 1005415
rect 446666 1005375 446672 1005387
rect 469840 1005375 469846 1005387
rect 469898 1005375 469904 1005427
rect 554512 1005375 554518 1005427
rect 554570 1005415 554576 1005427
rect 570448 1005415 570454 1005427
rect 554570 1005387 570454 1005415
rect 554570 1005375 554576 1005387
rect 570448 1005375 570454 1005387
rect 570506 1005375 570512 1005427
rect 92656 1005301 92662 1005353
rect 92714 1005341 92720 1005353
rect 101488 1005341 101494 1005353
rect 92714 1005313 101494 1005341
rect 92714 1005301 92720 1005313
rect 101488 1005301 101494 1005313
rect 101546 1005301 101552 1005353
rect 298672 1005301 298678 1005353
rect 298730 1005341 298736 1005353
rect 309616 1005341 309622 1005353
rect 298730 1005313 309622 1005341
rect 298730 1005301 298736 1005313
rect 309616 1005301 309622 1005313
rect 309674 1005301 309680 1005353
rect 358672 1005301 358678 1005353
rect 358730 1005341 358736 1005353
rect 366256 1005341 366262 1005353
rect 358730 1005313 366262 1005341
rect 358730 1005301 358736 1005313
rect 366256 1005301 366262 1005313
rect 366314 1005301 366320 1005353
rect 431536 1005301 431542 1005353
rect 431594 1005341 431600 1005353
rect 446320 1005341 446326 1005353
rect 431594 1005313 446326 1005341
rect 431594 1005301 431600 1005313
rect 446320 1005301 446326 1005313
rect 446378 1005301 446384 1005353
rect 446416 1005301 446422 1005353
rect 446474 1005341 446480 1005353
rect 470032 1005341 470038 1005353
rect 446474 1005313 470038 1005341
rect 446474 1005301 446480 1005313
rect 470032 1005301 470038 1005313
rect 470090 1005301 470096 1005353
rect 556912 1005301 556918 1005353
rect 556970 1005341 556976 1005353
rect 574480 1005341 574486 1005353
rect 556970 1005313 574486 1005341
rect 556970 1005301 556976 1005313
rect 574480 1005301 574486 1005313
rect 574538 1005301 574544 1005353
rect 92944 1005227 92950 1005279
rect 93002 1005267 93008 1005279
rect 114160 1005267 114166 1005279
rect 93002 1005239 114166 1005267
rect 93002 1005227 93008 1005239
rect 114160 1005227 114166 1005239
rect 114218 1005227 114224 1005279
rect 298768 1005227 298774 1005279
rect 298826 1005267 298832 1005279
rect 308752 1005267 308758 1005279
rect 298826 1005239 308758 1005267
rect 298826 1005227 298832 1005239
rect 308752 1005227 308758 1005239
rect 308810 1005227 308816 1005279
rect 318640 1005227 318646 1005279
rect 318698 1005267 318704 1005279
rect 328720 1005267 328726 1005279
rect 318698 1005239 328726 1005267
rect 318698 1005227 318704 1005239
rect 328720 1005227 328726 1005239
rect 328778 1005227 328784 1005279
rect 359920 1005227 359926 1005279
rect 359978 1005267 359984 1005279
rect 381712 1005267 381718 1005279
rect 359978 1005239 368702 1005267
rect 359978 1005227 359984 1005239
rect 92464 1005153 92470 1005205
rect 92522 1005193 92528 1005205
rect 105424 1005193 105430 1005205
rect 92522 1005165 105430 1005193
rect 92522 1005153 92528 1005165
rect 105424 1005153 105430 1005165
rect 105482 1005153 105488 1005205
rect 195472 1005153 195478 1005205
rect 195530 1005193 195536 1005205
rect 209008 1005193 209014 1005205
rect 195530 1005165 209014 1005193
rect 195530 1005153 195536 1005165
rect 209008 1005153 209014 1005165
rect 209066 1005153 209072 1005205
rect 299536 1005153 299542 1005205
rect 299594 1005193 299600 1005205
rect 310288 1005193 310294 1005205
rect 299594 1005165 310294 1005193
rect 299594 1005153 299600 1005165
rect 310288 1005153 310294 1005165
rect 310346 1005153 310352 1005205
rect 325456 1005153 325462 1005205
rect 325514 1005193 325520 1005205
rect 331216 1005193 331222 1005205
rect 325514 1005165 331222 1005193
rect 325514 1005153 325520 1005165
rect 331216 1005153 331222 1005165
rect 331274 1005153 331280 1005205
rect 357040 1005153 357046 1005205
rect 357098 1005193 357104 1005205
rect 368560 1005193 368566 1005205
rect 357098 1005165 368566 1005193
rect 357098 1005153 357104 1005165
rect 368560 1005153 368566 1005165
rect 368618 1005153 368624 1005205
rect 368674 1005193 368702 1005239
rect 368866 1005239 381718 1005267
rect 368866 1005193 368894 1005239
rect 381712 1005227 381718 1005239
rect 381770 1005227 381776 1005279
rect 425296 1005227 425302 1005279
rect 425354 1005267 425360 1005279
rect 463600 1005267 463606 1005279
rect 425354 1005239 463606 1005267
rect 425354 1005227 425360 1005239
rect 463600 1005227 463606 1005239
rect 463658 1005227 463664 1005279
rect 500656 1005227 500662 1005279
rect 500714 1005267 500720 1005279
rect 512560 1005267 512566 1005279
rect 500714 1005239 512566 1005267
rect 500714 1005227 500720 1005239
rect 512560 1005227 512566 1005239
rect 512618 1005227 512624 1005279
rect 368674 1005165 368894 1005193
rect 368962 1005165 380126 1005193
rect 364240 1005079 364246 1005131
rect 364298 1005119 364304 1005131
rect 368962 1005119 368990 1005165
rect 364298 1005091 368990 1005119
rect 380098 1005119 380126 1005165
rect 427600 1005153 427606 1005205
rect 427658 1005193 427664 1005205
rect 466576 1005193 466582 1005205
rect 427658 1005165 466582 1005193
rect 427658 1005153 427664 1005165
rect 466576 1005153 466582 1005165
rect 466634 1005153 466640 1005205
rect 501136 1005153 501142 1005205
rect 501194 1005193 501200 1005205
rect 512464 1005193 512470 1005205
rect 501194 1005165 512470 1005193
rect 501194 1005153 501200 1005165
rect 512464 1005153 512470 1005165
rect 512522 1005153 512528 1005205
rect 553744 1005153 553750 1005205
rect 553802 1005193 553808 1005205
rect 558736 1005193 558742 1005205
rect 553802 1005165 558742 1005193
rect 553802 1005153 553808 1005165
rect 558736 1005153 558742 1005165
rect 558794 1005153 558800 1005205
rect 562480 1005153 562486 1005205
rect 562538 1005193 562544 1005205
rect 570544 1005193 570550 1005205
rect 562538 1005165 570550 1005193
rect 562538 1005153 562544 1005165
rect 570544 1005153 570550 1005165
rect 570602 1005153 570608 1005205
rect 382960 1005119 382966 1005131
rect 380098 1005091 382966 1005119
rect 364298 1005079 364304 1005091
rect 382960 1005079 382966 1005091
rect 383018 1005079 383024 1005131
rect 435568 1005079 435574 1005131
rect 435626 1005119 435632 1005131
rect 440656 1005119 440662 1005131
rect 435626 1005091 440662 1005119
rect 435626 1005079 435632 1005091
rect 440656 1005079 440662 1005091
rect 440714 1005079 440720 1005131
rect 428080 1003895 428086 1003947
rect 428138 1003935 428144 1003947
rect 457840 1003935 457846 1003947
rect 428138 1003907 457846 1003935
rect 428138 1003895 428144 1003907
rect 457840 1003895 457846 1003907
rect 457898 1003895 457904 1003947
rect 357616 1003821 357622 1003873
rect 357674 1003861 357680 1003873
rect 380080 1003861 380086 1003873
rect 357674 1003833 380086 1003861
rect 357674 1003821 357680 1003833
rect 380080 1003821 380086 1003833
rect 380138 1003821 380144 1003873
rect 426448 1003821 426454 1003873
rect 426506 1003861 426512 1003873
rect 456304 1003861 456310 1003873
rect 426506 1003833 456310 1003861
rect 426506 1003821 426512 1003833
rect 456304 1003821 456310 1003833
rect 456362 1003821 456368 1003873
rect 554896 1003821 554902 1003873
rect 554954 1003861 554960 1003873
rect 567184 1003861 567190 1003873
rect 554954 1003833 567190 1003861
rect 554954 1003821 554960 1003833
rect 567184 1003821 567190 1003833
rect 567242 1003821 567248 1003873
rect 359056 1003747 359062 1003799
rect 359114 1003787 359120 1003799
rect 378256 1003787 378262 1003799
rect 359114 1003759 378262 1003787
rect 359114 1003747 359120 1003759
rect 378256 1003747 378262 1003759
rect 378314 1003747 378320 1003799
rect 423376 1003747 423382 1003799
rect 423434 1003787 423440 1003799
rect 466480 1003787 466486 1003799
rect 423434 1003759 466486 1003787
rect 423434 1003747 423440 1003759
rect 466480 1003747 466486 1003759
rect 466538 1003747 466544 1003799
rect 498160 1003747 498166 1003799
rect 498218 1003787 498224 1003799
rect 515728 1003787 515734 1003799
rect 498218 1003759 515734 1003787
rect 498218 1003747 498224 1003759
rect 515728 1003747 515734 1003759
rect 515786 1003747 515792 1003799
rect 92368 1003673 92374 1003725
rect 92426 1003713 92432 1003725
rect 108880 1003713 108886 1003725
rect 92426 1003685 108886 1003713
rect 92426 1003673 92432 1003685
rect 108880 1003673 108886 1003685
rect 108938 1003673 108944 1003725
rect 355984 1003673 355990 1003725
rect 356042 1003713 356048 1003725
rect 379312 1003713 379318 1003725
rect 356042 1003685 379318 1003713
rect 356042 1003673 356048 1003685
rect 379312 1003673 379318 1003685
rect 379370 1003673 379376 1003725
rect 425776 1003673 425782 1003725
rect 425834 1003713 425840 1003725
rect 471760 1003713 471766 1003725
rect 425834 1003685 471766 1003713
rect 425834 1003673 425840 1003685
rect 471760 1003673 471766 1003685
rect 471818 1003673 471824 1003725
rect 555664 1003673 555670 1003725
rect 555722 1003713 555728 1003725
rect 567280 1003713 567286 1003725
rect 555722 1003685 567286 1003713
rect 555722 1003673 555728 1003685
rect 567280 1003673 567286 1003685
rect 567338 1003673 567344 1003725
rect 501040 1002563 501046 1002615
rect 501098 1002603 501104 1002615
rect 519280 1002603 519286 1002615
rect 501098 1002575 519286 1002603
rect 501098 1002563 501104 1002575
rect 519280 1002563 519286 1002575
rect 519338 1002563 519344 1002615
rect 143728 1002489 143734 1002541
rect 143786 1002529 143792 1002541
rect 157936 1002529 157942 1002541
rect 143786 1002501 157942 1002529
rect 143786 1002489 143792 1002501
rect 157936 1002489 157942 1002501
rect 157994 1002489 158000 1002541
rect 503440 1002489 503446 1002541
rect 503498 1002529 503504 1002541
rect 503498 1002501 509726 1002529
rect 503498 1002489 503504 1002501
rect 97840 1002415 97846 1002467
rect 97898 1002455 97904 1002467
rect 102832 1002455 102838 1002467
rect 97898 1002427 102838 1002455
rect 97898 1002415 97904 1002427
rect 102832 1002415 102838 1002427
rect 102890 1002415 102896 1002467
rect 144016 1002415 144022 1002467
rect 144074 1002455 144080 1002467
rect 151216 1002455 151222 1002467
rect 144074 1002427 151222 1002455
rect 144074 1002415 144080 1002427
rect 151216 1002415 151222 1002427
rect 151274 1002415 151280 1002467
rect 99760 1002341 99766 1002393
rect 99818 1002381 99824 1002393
rect 103792 1002381 103798 1002393
rect 99818 1002353 103798 1002381
rect 99818 1002341 99824 1002353
rect 103792 1002341 103798 1002353
rect 103850 1002341 103856 1002393
rect 143920 1002341 143926 1002393
rect 143978 1002381 143984 1002393
rect 150352 1002381 150358 1002393
rect 143978 1002353 150358 1002381
rect 143978 1002341 143984 1002353
rect 150352 1002341 150358 1002353
rect 150410 1002341 150416 1002393
rect 509698 1002381 509726 1002501
rect 559120 1002489 559126 1002541
rect 559178 1002529 559184 1002541
rect 566128 1002529 566134 1002541
rect 559178 1002501 566134 1002529
rect 559178 1002489 559184 1002501
rect 566128 1002489 566134 1002501
rect 566186 1002489 566192 1002541
rect 560560 1002415 560566 1002467
rect 560618 1002455 560624 1002467
rect 566416 1002455 566422 1002467
rect 560618 1002427 566422 1002455
rect 560618 1002415 560624 1002427
rect 566416 1002415 566422 1002427
rect 566474 1002415 566480 1002467
rect 517168 1002381 517174 1002393
rect 509698 1002353 517174 1002381
rect 517168 1002341 517174 1002353
rect 517226 1002341 517232 1002393
rect 560080 1002341 560086 1002393
rect 560138 1002381 560144 1002393
rect 564688 1002381 564694 1002393
rect 560138 1002353 564694 1002381
rect 560138 1002341 560144 1002353
rect 564688 1002341 564694 1002353
rect 564746 1002341 564752 1002393
rect 564784 1002341 564790 1002393
rect 564842 1002381 564848 1002393
rect 567664 1002381 567670 1002393
rect 564842 1002353 567670 1002381
rect 564842 1002341 564848 1002353
rect 567664 1002341 567670 1002353
rect 567722 1002341 567728 1002393
rect 97744 1002267 97750 1002319
rect 97802 1002307 97808 1002319
rect 100528 1002307 100534 1002319
rect 97802 1002279 100534 1002307
rect 97802 1002267 97808 1002279
rect 100528 1002267 100534 1002279
rect 100586 1002267 100592 1002319
rect 100720 1002267 100726 1002319
rect 100778 1002307 100784 1002319
rect 104464 1002307 104470 1002319
rect 100778 1002279 104470 1002307
rect 100778 1002267 100784 1002279
rect 104464 1002267 104470 1002279
rect 104522 1002267 104528 1002319
rect 144112 1002267 144118 1002319
rect 144170 1002307 144176 1002319
rect 178480 1002307 178486 1002319
rect 144170 1002279 178486 1002307
rect 144170 1002267 144176 1002279
rect 178480 1002267 178486 1002279
rect 178538 1002267 178544 1002319
rect 446032 1002267 446038 1002319
rect 446090 1002307 446096 1002319
rect 446512 1002307 446518 1002319
rect 446090 1002279 446518 1002307
rect 446090 1002267 446096 1002279
rect 446512 1002267 446518 1002279
rect 446570 1002267 446576 1002319
rect 505072 1002267 505078 1002319
rect 505130 1002307 505136 1002319
rect 523600 1002307 523606 1002319
rect 505130 1002279 523606 1002307
rect 505130 1002267 505136 1002279
rect 523600 1002267 523606 1002279
rect 523658 1002267 523664 1002319
rect 561520 1002267 561526 1002319
rect 561578 1002307 561584 1002319
rect 565168 1002307 565174 1002319
rect 561578 1002279 565174 1002307
rect 561578 1002267 561584 1002279
rect 565168 1002267 565174 1002279
rect 565226 1002267 565232 1002319
rect 378256 1001897 378262 1001949
rect 378314 1001937 378320 1001949
rect 380464 1001937 380470 1001949
rect 378314 1001909 380470 1001937
rect 378314 1001897 378320 1001909
rect 380464 1001897 380470 1001909
rect 380522 1001897 380528 1001949
rect 446512 1001157 446518 1001209
rect 446570 1001197 446576 1001209
rect 467056 1001197 467062 1001209
rect 446570 1001169 467062 1001197
rect 446570 1001157 446576 1001169
rect 467056 1001157 467062 1001169
rect 467114 1001157 467120 1001209
rect 434032 1001083 434038 1001135
rect 434090 1001123 434096 1001135
rect 472624 1001123 472630 1001135
rect 434090 1001095 472630 1001123
rect 434090 1001083 434096 1001095
rect 472624 1001083 472630 1001095
rect 472682 1001083 472688 1001135
rect 195280 1001009 195286 1001061
rect 195338 1001049 195344 1001061
rect 208336 1001049 208342 1001061
rect 195338 1001021 208342 1001049
rect 195338 1001009 195344 1001021
rect 208336 1001009 208342 1001021
rect 208394 1001009 208400 1001061
rect 446416 1001009 446422 1001061
rect 446474 1001049 446480 1001061
rect 472336 1001049 472342 1001061
rect 446474 1001021 472342 1001049
rect 446474 1001009 446480 1001021
rect 472336 1001009 472342 1001021
rect 472394 1001009 472400 1001061
rect 564688 1001009 564694 1001061
rect 564746 1001049 564752 1001061
rect 570160 1001049 570166 1001061
rect 564746 1001021 570166 1001049
rect 564746 1001009 564752 1001021
rect 570160 1001009 570166 1001021
rect 570218 1001009 570224 1001061
rect 432496 1000935 432502 1000987
rect 432554 1000975 432560 1000987
rect 472624 1000975 472630 1000987
rect 432554 1000947 472630 1000975
rect 432554 1000935 432560 1000947
rect 472624 1000935 472630 1000947
rect 472682 1000935 472688 1000987
rect 361552 1000861 361558 1000913
rect 361610 1000901 361616 1000913
rect 383632 1000901 383638 1000913
rect 361610 1000873 383638 1000901
rect 361610 1000861 361616 1000873
rect 383632 1000861 383638 1000873
rect 383690 1000861 383696 1000913
rect 428944 1000861 428950 1000913
rect 429002 1000901 429008 1000913
rect 472528 1000901 472534 1000913
rect 429002 1000873 472534 1000901
rect 429002 1000861 429008 1000873
rect 472528 1000861 472534 1000873
rect 472586 1000861 472592 1000913
rect 565168 1000861 565174 1000913
rect 565226 1000901 565232 1000913
rect 568336 1000901 568342 1000913
rect 565226 1000873 568342 1000901
rect 565226 1000861 565232 1000873
rect 568336 1000861 568342 1000873
rect 568394 1000861 568400 1000913
rect 143824 1000787 143830 1000839
rect 143882 1000827 143888 1000839
rect 160240 1000827 160246 1000839
rect 143882 1000799 160246 1000827
rect 143882 1000787 143888 1000799
rect 160240 1000787 160246 1000799
rect 160298 1000787 160304 1000839
rect 195376 1000787 195382 1000839
rect 195434 1000827 195440 1000839
rect 211696 1000827 211702 1000839
rect 195434 1000799 211702 1000827
rect 195434 1000787 195440 1000799
rect 211696 1000787 211702 1000799
rect 211754 1000787 211760 1000839
rect 360688 1000787 360694 1000839
rect 360746 1000827 360752 1000839
rect 383536 1000827 383542 1000839
rect 360746 1000799 383542 1000827
rect 360746 1000787 360752 1000799
rect 383536 1000787 383542 1000799
rect 383594 1000787 383600 1000839
rect 424144 1000787 424150 1000839
rect 424202 1000827 424208 1000839
rect 471952 1000827 471958 1000839
rect 424202 1000799 471958 1000827
rect 424202 1000787 424208 1000799
rect 471952 1000787 471958 1000799
rect 472010 1000787 472016 1000839
rect 463696 1000713 463702 1000765
rect 463754 1000753 463760 1000765
rect 472144 1000753 472150 1000765
rect 463754 1000725 472150 1000753
rect 463754 1000713 463760 1000725
rect 472144 1000713 472150 1000725
rect 472202 1000713 472208 1000765
rect 509392 1000639 509398 1000691
rect 509450 1000679 509456 1000691
rect 516688 1000679 516694 1000691
rect 509450 1000651 516694 1000679
rect 509450 1000639 509456 1000651
rect 516688 1000639 516694 1000651
rect 516746 1000639 516752 1000691
rect 456304 1000269 456310 1000321
rect 456362 1000309 456368 1000321
rect 458800 1000309 458806 1000321
rect 456362 1000281 458806 1000309
rect 456362 1000269 456368 1000281
rect 458800 1000269 458806 1000281
rect 458858 1000269 458864 1000321
rect 298096 999973 298102 1000025
rect 298154 1000013 298160 1000025
rect 308080 1000013 308086 1000025
rect 298154 999985 308086 1000013
rect 298154 999973 298160 999985
rect 308080 999973 308086 999985
rect 308138 999973 308144 1000025
rect 503056 999899 503062 999951
rect 503114 999939 503120 999951
rect 516688 999939 516694 999951
rect 503114 999911 516694 999939
rect 503114 999899 503120 999911
rect 516688 999899 516694 999911
rect 516746 999899 516752 999951
rect 509872 999751 509878 999803
rect 509930 999791 509936 999803
rect 521680 999791 521686 999803
rect 509930 999763 521686 999791
rect 509930 999751 509936 999763
rect 521680 999751 521686 999763
rect 521738 999751 521744 999803
rect 298288 999677 298294 999729
rect 298346 999717 298352 999729
rect 298346 999689 318302 999717
rect 298346 999677 298352 999689
rect 298576 999529 298582 999581
rect 298634 999569 298640 999581
rect 315472 999569 315478 999581
rect 298634 999541 315478 999569
rect 298634 999529 298640 999541
rect 315472 999529 315478 999541
rect 315530 999529 315536 999581
rect 92752 999455 92758 999507
rect 92810 999495 92816 999507
rect 97744 999495 97750 999507
rect 92810 999467 97750 999495
rect 92810 999455 92816 999467
rect 97744 999455 97750 999467
rect 97802 999455 97808 999507
rect 246928 999455 246934 999507
rect 246986 999495 246992 999507
rect 256432 999495 256438 999507
rect 246986 999467 256438 999495
rect 246986 999455 246992 999467
rect 256432 999455 256438 999467
rect 256490 999455 256496 999507
rect 298192 999455 298198 999507
rect 298250 999495 298256 999507
rect 314704 999495 314710 999507
rect 298250 999467 314710 999495
rect 298250 999455 298256 999467
rect 314704 999455 314710 999467
rect 314762 999455 314768 999507
rect 92848 999381 92854 999433
rect 92906 999421 92912 999433
rect 126640 999421 126646 999433
rect 92906 999393 126646 999421
rect 92906 999381 92912 999393
rect 126640 999381 126646 999393
rect 126698 999381 126704 999433
rect 143728 999381 143734 999433
rect 143786 999421 143792 999433
rect 156880 999421 156886 999433
rect 143786 999393 156886 999421
rect 143786 999381 143792 999393
rect 156880 999381 156886 999393
rect 156938 999381 156944 999433
rect 195760 999381 195766 999433
rect 195818 999421 195824 999433
rect 224656 999421 224662 999433
rect 195818 999393 224662 999421
rect 195818 999381 195824 999393
rect 224656 999381 224662 999393
rect 224714 999381 224720 999433
rect 246544 999381 246550 999433
rect 246602 999421 246608 999433
rect 259504 999421 259510 999433
rect 246602 999393 259510 999421
rect 246602 999381 246608 999393
rect 259504 999381 259510 999393
rect 259562 999381 259568 999433
rect 298096 999381 298102 999433
rect 298154 999421 298160 999433
rect 311440 999421 311446 999433
rect 298154 999393 311446 999421
rect 298154 999381 298160 999393
rect 311440 999381 311446 999393
rect 311498 999381 311504 999433
rect 318274 999421 318302 999689
rect 506224 999677 506230 999729
rect 506282 999717 506288 999729
rect 516784 999717 516790 999729
rect 506282 999689 516790 999717
rect 506282 999677 506288 999689
rect 516784 999677 516790 999689
rect 516842 999677 516848 999729
rect 616048 999677 616054 999729
rect 616106 999717 616112 999729
rect 625744 999717 625750 999729
rect 616106 999689 625750 999717
rect 616106 999677 616112 999689
rect 625744 999677 625750 999689
rect 625802 999677 625808 999729
rect 507760 999603 507766 999655
rect 507818 999643 507824 999655
rect 521584 999643 521590 999655
rect 507818 999615 521590 999643
rect 507818 999603 507824 999615
rect 521584 999603 521590 999615
rect 521642 999603 521648 999655
rect 540304 999603 540310 999655
rect 540362 999643 540368 999655
rect 540362 999615 555998 999643
rect 540362 999603 540368 999615
rect 502384 999529 502390 999581
rect 502442 999569 502448 999581
rect 516784 999569 516790 999581
rect 502442 999541 516790 999569
rect 502442 999529 502448 999541
rect 516784 999529 516790 999541
rect 516842 999529 516848 999581
rect 466576 999455 466582 999507
rect 466634 999495 466640 999507
rect 472432 999495 472438 999507
rect 466634 999467 472438 999495
rect 466634 999455 466640 999467
rect 472432 999455 472438 999467
rect 472490 999455 472496 999507
rect 508624 999455 508630 999507
rect 508682 999495 508688 999507
rect 523984 999495 523990 999507
rect 508682 999467 523990 999495
rect 508682 999455 508688 999467
rect 523984 999455 523990 999467
rect 524042 999455 524048 999507
rect 331792 999421 331798 999433
rect 318274 999393 331798 999421
rect 331792 999381 331798 999393
rect 331850 999381 331856 999433
rect 399952 999381 399958 999433
rect 400010 999421 400016 999433
rect 471664 999421 471670 999433
rect 400010 999393 471670 999421
rect 400010 999381 400016 999393
rect 471664 999381 471670 999393
rect 471722 999381 471728 999433
rect 488944 999381 488950 999433
rect 489002 999421 489008 999433
rect 489002 999393 519806 999421
rect 489002 999381 489008 999393
rect 368560 999307 368566 999359
rect 368618 999347 368624 999359
rect 383056 999347 383062 999359
rect 368618 999319 383062 999347
rect 368618 999307 368624 999319
rect 383056 999307 383062 999319
rect 383114 999307 383120 999359
rect 422512 999307 422518 999359
rect 422570 999347 422576 999359
rect 429136 999347 429142 999359
rect 422570 999319 429142 999347
rect 422570 999307 422576 999319
rect 429136 999307 429142 999319
rect 429194 999307 429200 999359
rect 497584 999307 497590 999359
rect 497642 999347 497648 999359
rect 516880 999347 516886 999359
rect 497642 999319 516886 999347
rect 497642 999307 497648 999319
rect 516880 999307 516886 999319
rect 516938 999307 516944 999359
rect 519778 999347 519806 999393
rect 552976 999381 552982 999433
rect 553034 999421 553040 999433
rect 555856 999421 555862 999433
rect 553034 999393 555862 999421
rect 553034 999381 553040 999393
rect 555856 999381 555862 999393
rect 555914 999381 555920 999433
rect 555970 999421 555998 999615
rect 616144 999603 616150 999655
rect 616202 999643 616208 999655
rect 625840 999643 625846 999655
rect 616202 999615 625846 999643
rect 616202 999603 616208 999615
rect 625840 999603 625846 999615
rect 625898 999603 625904 999655
rect 600400 999529 600406 999581
rect 600458 999569 600464 999581
rect 600458 999541 616286 999569
rect 600458 999529 600464 999541
rect 598768 999455 598774 999507
rect 598826 999495 598832 999507
rect 616048 999495 616054 999507
rect 598826 999467 616054 999495
rect 598826 999455 598832 999467
rect 616048 999455 616054 999467
rect 616106 999455 616112 999507
rect 616258 999495 616286 999541
rect 625648 999495 625654 999507
rect 616258 999467 625654 999495
rect 625648 999455 625654 999467
rect 625706 999455 625712 999507
rect 572464 999421 572470 999433
rect 555970 999393 572470 999421
rect 572464 999381 572470 999393
rect 572522 999381 572528 999433
rect 596080 999381 596086 999433
rect 596138 999421 596144 999433
rect 616144 999421 616150 999433
rect 596138 999393 616150 999421
rect 596138 999381 596144 999393
rect 616144 999381 616150 999393
rect 616202 999381 616208 999433
rect 616240 999381 616246 999433
rect 616298 999421 616304 999433
rect 625840 999421 625846 999433
rect 616298 999393 625846 999421
rect 616298 999381 616304 999393
rect 625840 999381 625846 999393
rect 625898 999381 625904 999433
rect 521296 999347 521302 999359
rect 519778 999319 521302 999347
rect 521296 999307 521302 999319
rect 521354 999307 521360 999359
rect 366256 999233 366262 999285
rect 366314 999273 366320 999285
rect 383248 999273 383254 999285
rect 366314 999245 383254 999273
rect 366314 999233 366320 999245
rect 383248 999233 383254 999245
rect 383306 999233 383312 999285
rect 512464 999233 512470 999285
rect 512522 999273 512528 999285
rect 521776 999273 521782 999285
rect 512522 999245 521782 999273
rect 512522 999233 512528 999245
rect 521776 999233 521782 999245
rect 521834 999233 521840 999285
rect 566128 999233 566134 999285
rect 566186 999273 566192 999285
rect 573040 999273 573046 999285
rect 566186 999245 573046 999273
rect 566186 999233 566192 999245
rect 573040 999233 573046 999245
rect 573098 999233 573104 999285
rect 567184 999159 567190 999211
rect 567242 999199 567248 999211
rect 575344 999199 575350 999211
rect 567242 999171 575350 999199
rect 567242 999159 567248 999171
rect 575344 999159 575350 999171
rect 575402 999159 575408 999211
rect 460816 999085 460822 999137
rect 460874 999125 460880 999137
rect 471856 999125 471862 999137
rect 460874 999097 471862 999125
rect 460874 999085 460880 999097
rect 471856 999085 471862 999097
rect 471914 999085 471920 999137
rect 567376 998567 567382 998619
rect 567434 998607 567440 998619
rect 575440 998607 575446 998619
rect 567434 998579 575446 998607
rect 567434 998567 567440 998579
rect 575440 998567 575446 998579
rect 575498 998567 575504 998619
rect 568336 998271 568342 998323
rect 568394 998311 568400 998323
rect 572944 998311 572950 998323
rect 568394 998283 572950 998311
rect 568394 998271 568400 998283
rect 572944 998271 572950 998283
rect 573002 998271 573008 998323
rect 320944 997901 320950 997953
rect 321002 997941 321008 997953
rect 367888 997941 367894 997953
rect 321002 997913 367894 997941
rect 321002 997901 321008 997913
rect 367888 997901 367894 997913
rect 367946 997941 367952 997953
rect 380176 997941 380182 997953
rect 367946 997913 380182 997941
rect 367946 997901 367952 997913
rect 380176 997901 380182 997913
rect 380234 997901 380240 997953
rect 572464 997901 572470 997953
rect 572522 997941 572528 997953
rect 617776 997941 617782 997953
rect 572522 997913 617782 997941
rect 572522 997901 572528 997913
rect 617776 997901 617782 997913
rect 617834 997901 617840 997953
rect 331792 997827 331798 997879
rect 331850 997867 331856 997879
rect 383152 997867 383158 997879
rect 331850 997839 383158 997867
rect 331850 997827 331856 997839
rect 383152 997827 383158 997839
rect 383210 997827 383216 997879
rect 557296 997827 557302 997879
rect 557354 997867 557360 997879
rect 596080 997867 596086 997879
rect 557354 997839 596086 997867
rect 557354 997827 557360 997839
rect 596080 997827 596086 997839
rect 596138 997827 596144 997879
rect 302416 997753 302422 997805
rect 302474 997793 302480 997805
rect 348688 997793 348694 997805
rect 302474 997765 348694 997793
rect 302474 997753 302480 997765
rect 348688 997753 348694 997765
rect 348746 997753 348752 997805
rect 566416 997753 566422 997805
rect 566474 997793 566480 997805
rect 598768 997793 598774 997805
rect 566474 997765 598774 997793
rect 566474 997753 566480 997765
rect 598768 997753 598774 997765
rect 598826 997753 598832 997805
rect 328720 997679 328726 997731
rect 328778 997719 328784 997731
rect 369040 997719 369046 997731
rect 328778 997691 369046 997719
rect 328778 997679 328784 997691
rect 369040 997679 369046 997691
rect 369098 997679 369104 997731
rect 457936 997679 457942 997731
rect 457994 997719 458000 997731
rect 472240 997719 472246 997731
rect 457994 997691 472246 997719
rect 457994 997679 458000 997691
rect 472240 997679 472246 997691
rect 472298 997679 472304 997731
rect 574480 997679 574486 997731
rect 574538 997719 574544 997731
rect 619120 997719 619126 997731
rect 574538 997691 619126 997719
rect 574538 997679 574544 997691
rect 619120 997679 619126 997691
rect 619178 997679 619184 997731
rect 570544 997605 570550 997657
rect 570602 997645 570608 997657
rect 600400 997645 600406 997657
rect 570602 997617 600406 997645
rect 570602 997605 570608 997617
rect 600400 997605 600406 997617
rect 600458 997605 600464 997657
rect 570448 997531 570454 997583
rect 570506 997571 570512 997583
rect 616240 997571 616246 997583
rect 570506 997543 616246 997571
rect 570506 997531 570512 997543
rect 616240 997531 616246 997543
rect 616298 997531 616304 997583
rect 458800 996791 458806 996843
rect 458858 996831 458864 996843
rect 472048 996831 472054 996843
rect 458858 996803 472054 996831
rect 458858 996791 458864 996803
rect 472048 996791 472054 996803
rect 472106 996791 472112 996843
rect 195184 996495 195190 996547
rect 195242 996535 195248 996547
rect 204208 996535 204214 996547
rect 195242 996507 204214 996535
rect 195242 996495 195248 996507
rect 204208 996495 204214 996507
rect 204266 996495 204272 996547
rect 251248 996495 251254 996547
rect 251306 996535 251312 996547
rect 263056 996535 263062 996547
rect 251306 996507 263062 996535
rect 251306 996495 251312 996507
rect 263056 996495 263062 996507
rect 263114 996495 263120 996547
rect 512656 996495 512662 996547
rect 512714 996535 512720 996547
rect 521488 996535 521494 996547
rect 512714 996507 521494 996535
rect 512714 996495 512720 996507
rect 521488 996495 521494 996507
rect 521546 996495 521552 996547
rect 555856 996495 555862 996547
rect 555914 996535 555920 996547
rect 561424 996535 561430 996547
rect 555914 996507 561430 996535
rect 555914 996495 555920 996507
rect 561424 996495 561430 996507
rect 561482 996495 561488 996547
rect 319792 996421 319798 996473
rect 319850 996461 319856 996473
rect 367120 996461 367126 996473
rect 319850 996433 367126 996461
rect 319850 996421 319856 996433
rect 367120 996421 367126 996433
rect 367178 996421 367184 996473
rect 604816 996347 604822 996399
rect 604874 996387 604880 996399
rect 624880 996387 624886 996399
rect 604874 996359 624886 996387
rect 604874 996347 604880 996359
rect 624880 996347 624886 996359
rect 624938 996347 624944 996399
rect 511888 996199 511894 996251
rect 511946 996239 511952 996251
rect 511946 996211 517310 996239
rect 511946 996199 511952 996211
rect 163120 996165 163126 996177
rect 136930 996137 163126 996165
rect 115312 996051 115318 996103
rect 115370 996091 115376 996103
rect 127504 996091 127510 996103
rect 115370 996063 127510 996091
rect 115370 996051 115376 996063
rect 127504 996051 127510 996063
rect 127562 996051 127568 996103
rect 136930 996091 136958 996137
rect 163120 996125 163126 996137
rect 163178 996165 163184 996177
rect 214096 996165 214102 996177
rect 163178 996137 214102 996165
rect 163178 996125 163184 996137
rect 214096 996125 214102 996137
rect 214154 996165 214160 996177
rect 265936 996165 265942 996177
rect 214154 996137 265942 996165
rect 214154 996125 214160 996137
rect 265936 996125 265942 996137
rect 265994 996165 266000 996177
rect 265994 996137 267134 996165
rect 265994 996125 266000 996137
rect 162256 996091 162262 996103
rect 127618 996063 136958 996091
rect 137218 996063 162262 996091
rect 127408 995977 127414 996029
rect 127466 996017 127472 996029
rect 127618 996017 127646 996063
rect 127466 995989 127646 996017
rect 127466 995977 127472 995989
rect 81634 995915 94046 995943
rect 81634 995807 81662 995915
rect 93904 995869 93910 995881
rect 89026 995841 93910 995869
rect 89026 995807 89054 995841
rect 93904 995829 93910 995841
rect 93962 995829 93968 995881
rect 94018 995869 94046 995915
rect 97840 995869 97846 995881
rect 94018 995841 97846 995869
rect 97840 995829 97846 995841
rect 97898 995829 97904 995881
rect 115216 995829 115222 995881
rect 115274 995869 115280 995881
rect 127408 995869 127414 995881
rect 115274 995841 127414 995869
rect 115274 995829 115280 995841
rect 127408 995829 127414 995841
rect 127466 995829 127472 995881
rect 127504 995829 127510 995881
rect 127562 995869 127568 995881
rect 137218 995869 137246 996063
rect 162256 996051 162262 996063
rect 162314 996091 162320 996103
rect 213328 996091 213334 996103
rect 162314 996063 213334 996091
rect 162314 996051 162320 996063
rect 213328 996051 213334 996063
rect 213386 996051 213392 996103
rect 215632 996051 215638 996103
rect 215690 996091 215696 996103
rect 266992 996091 266998 996103
rect 215690 996063 266998 996091
rect 215690 996051 215696 996063
rect 266992 996051 266998 996063
rect 267050 996051 267056 996103
rect 267106 996091 267134 996137
rect 270736 996125 270742 996177
rect 270794 996165 270800 996177
rect 318640 996165 318646 996177
rect 270794 996137 318646 996165
rect 270794 996125 270800 996137
rect 318640 996125 318646 996137
rect 318698 996125 318704 996177
rect 368656 996125 368662 996177
rect 368714 996165 368720 996177
rect 436336 996165 436342 996177
rect 368714 996137 436342 996165
rect 368714 996125 368720 996137
rect 436336 996125 436342 996137
rect 436394 996125 436400 996177
rect 436432 996125 436438 996177
rect 436490 996165 436496 996177
rect 513424 996165 513430 996177
rect 436490 996137 513430 996165
rect 436490 996125 436496 996137
rect 513424 996125 513430 996137
rect 513482 996125 513488 996177
rect 517282 996165 517310 996211
rect 563728 996165 563734 996177
rect 517282 996137 563734 996165
rect 563728 996125 563734 996137
rect 563786 996125 563792 996177
rect 317104 996091 317110 996103
rect 267106 996063 317110 996091
rect 317104 996051 317110 996063
rect 317162 996091 317168 996103
rect 320944 996091 320950 996103
rect 317162 996063 320950 996091
rect 317162 996051 317168 996063
rect 320944 996051 320950 996063
rect 321002 996051 321008 996103
rect 380176 996051 380182 996103
rect 380234 996091 380240 996103
rect 440656 996091 440662 996103
rect 380234 996063 440662 996091
rect 380234 996051 380240 996063
rect 440656 996051 440662 996063
rect 440714 996051 440720 996103
rect 470032 996051 470038 996103
rect 470090 996091 470096 996103
rect 511120 996091 511126 996103
rect 470090 996063 511126 996091
rect 470090 996051 470096 996063
rect 511120 996051 511126 996063
rect 511178 996091 511184 996103
rect 562864 996091 562870 996103
rect 511178 996063 562870 996091
rect 511178 996051 511184 996063
rect 562864 996051 562870 996063
rect 562922 996051 562928 996103
rect 164080 996017 164086 996029
rect 127562 995841 137246 995869
rect 137602 995989 164086 996017
rect 127562 995829 127568 995841
rect 137602 995807 137630 995989
rect 164080 995977 164086 995989
rect 164138 995977 164144 996029
rect 164176 995977 164182 996029
rect 164234 996017 164240 996029
rect 215440 996017 215446 996029
rect 164234 995989 215446 996017
rect 164234 995977 164240 995989
rect 215440 995977 215446 995989
rect 215498 995977 215504 996029
rect 264688 996017 264694 996029
rect 250402 995989 264694 996017
rect 151984 995943 151990 995955
rect 140146 995915 151990 995943
rect 81616 995755 81622 995807
rect 81674 995755 81680 995807
rect 89008 995755 89014 995807
rect 89066 995755 89072 995807
rect 91504 995755 91510 995807
rect 91562 995795 91568 995807
rect 92464 995795 92470 995807
rect 91562 995767 92470 995795
rect 91562 995755 91568 995767
rect 92464 995755 92470 995767
rect 92522 995755 92528 995807
rect 106096 995755 106102 995807
rect 106154 995795 106160 995807
rect 113296 995795 113302 995807
rect 106154 995767 113302 995795
rect 106154 995755 106160 995767
rect 113296 995755 113302 995767
rect 113354 995755 113360 995807
rect 113392 995755 113398 995807
rect 113450 995795 113456 995807
rect 118096 995795 118102 995807
rect 113450 995767 118102 995795
rect 113450 995755 113456 995767
rect 118096 995755 118102 995767
rect 118154 995755 118160 995807
rect 137584 995755 137590 995807
rect 137642 995755 137648 995807
rect 89776 995681 89782 995733
rect 89834 995721 89840 995733
rect 92368 995721 92374 995733
rect 89834 995693 92374 995721
rect 89834 995681 89840 995693
rect 92368 995681 92374 995693
rect 92426 995681 92432 995733
rect 133648 995681 133654 995733
rect 133706 995721 133712 995733
rect 140146 995721 140174 995915
rect 151984 995903 151990 995915
rect 152042 995903 152048 995955
rect 198640 995903 198646 995955
rect 198698 995943 198704 995955
rect 203440 995943 203446 995955
rect 198698 995915 203446 995943
rect 198698 995903 198704 995915
rect 203440 995903 203446 995915
rect 203498 995903 203504 995955
rect 213040 995903 213046 995955
rect 213098 995943 213104 995955
rect 217072 995943 217078 995955
rect 213098 995915 217078 995943
rect 213098 995903 213104 995915
rect 217072 995903 217078 995915
rect 217130 995903 217136 995955
rect 250402 995943 250430 995989
rect 264688 995977 264694 995989
rect 264746 996017 264752 996029
rect 267760 996017 267766 996029
rect 264746 995989 267766 996017
rect 264746 995977 264752 995989
rect 267760 995977 267766 995989
rect 267818 995977 267824 996029
rect 267856 995977 267862 996029
rect 267914 996017 267920 996029
rect 316336 996017 316342 996029
rect 267914 995989 316342 996017
rect 267914 995977 267920 995989
rect 316336 995977 316342 995989
rect 316394 996017 316400 996029
rect 319696 996017 319702 996029
rect 316394 995989 319702 996017
rect 316394 995977 316400 995989
rect 319696 995977 319702 995989
rect 319754 995977 319760 996029
rect 367120 995977 367126 996029
rect 367178 996017 367184 996029
rect 434128 996017 434134 996029
rect 367178 995989 434134 996017
rect 367178 995977 367184 995989
rect 434128 995977 434134 995989
rect 434186 996017 434192 996029
rect 439216 996017 439222 996029
rect 434186 995989 439222 996017
rect 434186 995977 434192 995989
rect 439216 995977 439222 995989
rect 439274 995977 439280 996029
rect 469840 995977 469846 996029
rect 469898 996017 469904 996029
rect 511888 996017 511894 996029
rect 469898 995989 511894 996017
rect 469898 995977 469904 995989
rect 511888 995977 511894 995989
rect 511946 995977 511952 996029
rect 513328 995977 513334 996029
rect 513386 996017 513392 996029
rect 564784 996017 564790 996029
rect 513386 995989 564790 996017
rect 513386 995977 513392 995989
rect 564784 995977 564790 995989
rect 564842 995977 564848 996029
rect 227458 995915 250430 995943
rect 144016 995829 144022 995881
rect 144074 995869 144080 995881
rect 155344 995869 155350 995881
rect 144074 995841 155350 995869
rect 144074 995829 144080 995841
rect 155344 995829 155350 995841
rect 155402 995829 155408 995881
rect 195472 995869 195478 995881
rect 187714 995841 195478 995869
rect 187714 995807 187742 995841
rect 195472 995829 195478 995841
rect 195530 995829 195536 995881
rect 213328 995829 213334 995881
rect 213386 995869 213392 995881
rect 227458 995869 227486 995915
rect 250480 995903 250486 995955
rect 250538 995943 250544 995955
rect 258832 995943 258838 995955
rect 250538 995915 258838 995943
rect 250538 995903 250544 995915
rect 258832 995903 258838 995915
rect 258890 995903 258896 995955
rect 299440 995943 299446 995955
rect 283810 995915 299446 995943
rect 213386 995841 227486 995869
rect 213386 995829 213392 995841
rect 250096 995829 250102 995881
rect 250154 995869 250160 995881
rect 255568 995869 255574 995881
rect 250154 995841 255574 995869
rect 250154 995829 250160 995841
rect 255568 995829 255574 995841
rect 255626 995829 255632 995881
rect 283810 995807 283838 995915
rect 299440 995903 299446 995915
rect 299498 995903 299504 995955
rect 472048 995903 472054 995955
rect 472106 995943 472112 995955
rect 472106 995915 483902 995943
rect 472106 995903 472112 995915
rect 298768 995869 298774 995881
rect 289474 995841 298774 995869
rect 289474 995807 289502 995841
rect 298768 995829 298774 995841
rect 298826 995829 298832 995881
rect 382960 995829 382966 995881
rect 383018 995869 383024 995881
rect 383018 995841 387518 995869
rect 383018 995829 383024 995841
rect 387490 995807 387518 995841
rect 472432 995829 472438 995881
rect 472490 995869 472496 995881
rect 472490 995841 477758 995869
rect 472490 995829 472496 995841
rect 477730 995807 477758 995841
rect 483874 995807 483902 995915
rect 524080 995903 524086 995955
rect 524138 995943 524144 995955
rect 524138 995915 533342 995943
rect 524138 995903 524144 995915
rect 523696 995829 523702 995881
rect 523754 995869 523760 995881
rect 523754 995841 529694 995869
rect 523754 995829 523760 995841
rect 142960 995755 142966 995807
rect 143018 995795 143024 995807
rect 143728 995795 143734 995807
rect 143018 995767 143734 995795
rect 143018 995755 143024 995767
rect 143728 995755 143734 995767
rect 143786 995755 143792 995807
rect 146800 995755 146806 995807
rect 146858 995795 146864 995807
rect 154288 995795 154294 995807
rect 146858 995767 154294 995795
rect 146858 995755 146864 995767
rect 154288 995755 154294 995767
rect 154346 995755 154352 995807
rect 164080 995755 164086 995807
rect 164138 995795 164144 995807
rect 165616 995795 165622 995807
rect 164138 995767 165622 995795
rect 164138 995755 164144 995767
rect 165616 995755 165622 995767
rect 165674 995755 165680 995807
rect 187696 995755 187702 995807
rect 187754 995755 187760 995807
rect 190576 995755 190582 995807
rect 190634 995795 190640 995807
rect 204976 995795 204982 995807
rect 190634 995767 204982 995795
rect 190634 995755 190640 995767
rect 204976 995755 204982 995767
rect 205034 995755 205040 995807
rect 224656 995755 224662 995807
rect 224714 995795 224720 995807
rect 224714 995767 236414 995795
rect 224714 995755 224720 995767
rect 133706 995693 140174 995721
rect 133706 995681 133712 995693
rect 141040 995681 141046 995733
rect 141098 995721 141104 995733
rect 143824 995721 143830 995733
rect 141098 995693 143830 995721
rect 141098 995681 141104 995693
rect 143824 995681 143830 995693
rect 143882 995681 143888 995733
rect 151696 995681 151702 995733
rect 151754 995721 151760 995733
rect 156304 995721 156310 995733
rect 151754 995693 156310 995721
rect 151754 995681 151760 995693
rect 156304 995681 156310 995693
rect 156362 995681 156368 995733
rect 163984 995681 163990 995733
rect 164042 995721 164048 995733
rect 166192 995721 166198 995733
rect 164042 995693 166198 995721
rect 164042 995681 164048 995693
rect 166192 995681 166198 995693
rect 166250 995681 166256 995733
rect 188080 995681 188086 995733
rect 188138 995721 188144 995733
rect 202864 995721 202870 995733
rect 188138 995693 202870 995721
rect 188138 995681 188144 995693
rect 202864 995681 202870 995693
rect 202922 995681 202928 995733
rect 194416 995607 194422 995659
rect 194474 995647 194480 995659
rect 195280 995647 195286 995659
rect 194474 995619 195286 995647
rect 194474 995607 194480 995619
rect 195280 995607 195286 995619
rect 195338 995607 195344 995659
rect 201616 995607 201622 995659
rect 201674 995647 201680 995659
rect 206992 995647 206998 995659
rect 201674 995619 206998 995647
rect 201674 995607 201680 995619
rect 206992 995607 206998 995619
rect 207050 995607 207056 995659
rect 236386 995647 236414 995767
rect 236464 995755 236470 995807
rect 236522 995795 236528 995807
rect 254800 995795 254806 995807
rect 236522 995767 254806 995795
rect 236522 995755 236528 995767
rect 254800 995755 254806 995767
rect 254858 995755 254864 995807
rect 268240 995755 268246 995807
rect 268298 995795 268304 995807
rect 273712 995795 273718 995807
rect 268298 995767 273718 995795
rect 268298 995755 268304 995767
rect 273712 995755 273718 995767
rect 273770 995755 273776 995807
rect 283792 995755 283798 995807
rect 283850 995755 283856 995807
rect 289456 995755 289462 995807
rect 289514 995755 289520 995807
rect 291184 995755 291190 995807
rect 291242 995795 291248 995807
rect 305584 995795 305590 995807
rect 291242 995767 305590 995795
rect 291242 995755 291248 995767
rect 305584 995755 305590 995767
rect 305642 995755 305648 995807
rect 366640 995755 366646 995807
rect 366698 995795 366704 995807
rect 371824 995795 371830 995807
rect 366698 995767 371830 995795
rect 366698 995755 366704 995767
rect 371824 995755 371830 995767
rect 371882 995755 371888 995807
rect 383632 995755 383638 995807
rect 383690 995795 383696 995807
rect 384976 995795 384982 995807
rect 383690 995767 384982 995795
rect 383690 995755 383696 995767
rect 384976 995755 384982 995767
rect 385034 995755 385040 995807
rect 387472 995755 387478 995807
rect 387530 995755 387536 995807
rect 396592 995755 396598 995807
rect 396650 995795 396656 995807
rect 399952 995795 399958 995807
rect 396650 995767 399958 995795
rect 396650 995755 396656 995767
rect 399952 995755 399958 995767
rect 400010 995755 400016 995807
rect 438736 995755 438742 995807
rect 438794 995795 438800 995807
rect 444496 995795 444502 995807
rect 438794 995767 444502 995795
rect 438794 995755 438800 995767
rect 444496 995755 444502 995767
rect 444554 995755 444560 995807
rect 472624 995755 472630 995807
rect 472682 995795 472688 995807
rect 473296 995795 473302 995807
rect 472682 995767 473302 995795
rect 472682 995755 472688 995767
rect 473296 995755 473302 995767
rect 473354 995755 473360 995807
rect 477712 995755 477718 995807
rect 477770 995755 477776 995807
rect 483856 995755 483862 995807
rect 483914 995755 483920 995807
rect 485680 995755 485686 995807
rect 485738 995795 485744 995807
rect 488944 995795 488950 995807
rect 485738 995767 488950 995795
rect 485738 995755 485744 995767
rect 488944 995755 488950 995767
rect 489002 995755 489008 995807
rect 504688 995755 504694 995807
rect 504746 995795 504752 995807
rect 518704 995795 518710 995807
rect 504746 995767 518710 995795
rect 504746 995755 504752 995767
rect 518704 995755 518710 995767
rect 518762 995755 518768 995807
rect 523888 995755 523894 995807
rect 523946 995795 523952 995807
rect 525328 995795 525334 995807
rect 523946 995767 525334 995795
rect 523946 995755 523952 995767
rect 525328 995755 525334 995767
rect 525386 995755 525392 995807
rect 529666 995795 529694 995841
rect 529840 995795 529846 995807
rect 529666 995767 529846 995795
rect 529840 995755 529846 995767
rect 529898 995755 529904 995807
rect 533314 995795 533342 995915
rect 567088 995903 567094 995955
rect 567146 995943 567152 995955
rect 570256 995943 570262 995955
rect 567146 995915 570262 995943
rect 567146 995903 567152 995915
rect 570256 995903 570262 995915
rect 570314 995903 570320 995955
rect 625840 995903 625846 995955
rect 625898 995943 625904 995955
rect 625898 995915 635102 995943
rect 625898 995903 625904 995915
rect 562864 995829 562870 995881
rect 562922 995869 562928 995881
rect 567376 995869 567382 995881
rect 562922 995841 567382 995869
rect 562922 995829 562928 995841
rect 567376 995829 567382 995841
rect 567434 995829 567440 995881
rect 619120 995829 619126 995881
rect 619178 995869 619184 995881
rect 635074 995869 635102 995915
rect 619178 995841 630206 995869
rect 635074 995841 635294 995869
rect 619178 995829 619184 995841
rect 630178 995807 630206 995841
rect 635266 995807 635294 995841
rect 533392 995795 533398 995807
rect 533314 995767 533398 995795
rect 533392 995755 533398 995767
rect 533450 995755 533456 995807
rect 537136 995755 537142 995807
rect 537194 995795 537200 995807
rect 540304 995795 540310 995807
rect 537194 995767 540310 995795
rect 537194 995755 537200 995767
rect 540304 995755 540310 995767
rect 540362 995755 540368 995807
rect 566320 995755 566326 995807
rect 566378 995795 566384 995807
rect 570352 995795 570358 995807
rect 566378 995767 570358 995795
rect 566378 995755 566384 995767
rect 570352 995755 570358 995767
rect 570410 995755 570416 995807
rect 625744 995755 625750 995807
rect 625802 995795 625808 995807
rect 626512 995795 626518 995807
rect 625802 995767 626518 995795
rect 625802 995755 625808 995767
rect 626512 995755 626518 995767
rect 626570 995755 626576 995807
rect 630160 995755 630166 995807
rect 630218 995755 630224 995807
rect 635248 995755 635254 995807
rect 635306 995755 635312 995807
rect 245680 995681 245686 995733
rect 245738 995721 245744 995733
rect 246544 995721 246550 995733
rect 245738 995693 246550 995721
rect 245738 995681 245744 995693
rect 246544 995681 246550 995693
rect 246602 995681 246608 995733
rect 247600 995681 247606 995733
rect 247658 995721 247664 995733
rect 257488 995721 257494 995733
rect 247658 995693 257494 995721
rect 247658 995681 247664 995693
rect 257488 995681 257494 995693
rect 257546 995681 257552 995733
rect 291760 995681 291766 995733
rect 291818 995721 291824 995733
rect 307408 995721 307414 995733
rect 291818 995693 307414 995721
rect 291818 995681 291824 995693
rect 307408 995681 307414 995693
rect 307466 995681 307472 995733
rect 365872 995681 365878 995733
rect 365930 995721 365936 995733
rect 377392 995721 377398 995733
rect 365930 995693 377398 995721
rect 365930 995681 365936 995693
rect 377392 995681 377398 995693
rect 377450 995681 377456 995733
rect 383536 995681 383542 995733
rect 383594 995721 383600 995733
rect 388048 995721 388054 995733
rect 383594 995693 388054 995721
rect 383594 995681 383600 995693
rect 388048 995681 388054 995693
rect 388106 995681 388112 995733
rect 472528 995681 472534 995733
rect 472586 995721 472592 995733
rect 474064 995721 474070 995733
rect 472586 995693 474070 995721
rect 472586 995681 472592 995693
rect 474064 995681 474070 995693
rect 474122 995681 474128 995733
rect 523792 995681 523798 995733
rect 523850 995721 523856 995733
rect 524752 995721 524758 995733
rect 523850 995693 524758 995721
rect 523850 995681 523856 995693
rect 524752 995681 524758 995693
rect 524810 995681 524816 995733
rect 563728 995681 563734 995733
rect 563786 995721 563792 995733
rect 567472 995721 567478 995733
rect 563786 995693 567478 995721
rect 563786 995681 563792 995693
rect 567472 995681 567478 995693
rect 567530 995681 567536 995733
rect 625936 995681 625942 995733
rect 625994 995721 626000 995733
rect 627088 995721 627094 995733
rect 625994 995693 627094 995721
rect 625994 995681 626000 995693
rect 627088 995681 627094 995693
rect 627146 995681 627152 995733
rect 237232 995647 237238 995659
rect 236386 995619 237238 995647
rect 237232 995607 237238 995619
rect 237290 995607 237296 995659
rect 253072 995607 253078 995659
rect 253130 995647 253136 995659
rect 258256 995647 258262 995659
rect 253130 995619 258262 995647
rect 253130 995607 253136 995619
rect 258256 995607 258262 995619
rect 258314 995607 258320 995659
rect 297328 995607 297334 995659
rect 297386 995647 297392 995659
rect 298096 995647 298102 995659
rect 297386 995619 298102 995647
rect 297386 995607 297392 995619
rect 298096 995607 298102 995619
rect 298154 995607 298160 995659
rect 383728 995607 383734 995659
rect 383786 995647 383792 995659
rect 384400 995647 384406 995659
rect 383786 995619 384406 995647
rect 383786 995607 383792 995619
rect 384400 995607 384406 995619
rect 384458 995607 384464 995659
rect 472720 995607 472726 995659
rect 472778 995647 472784 995659
rect 474640 995647 474646 995659
rect 472778 995619 474646 995647
rect 472778 995607 472784 995619
rect 474640 995607 474646 995619
rect 474698 995607 474704 995659
rect 523600 995607 523606 995659
rect 523658 995647 523664 995659
rect 528400 995647 528406 995659
rect 523658 995619 528406 995647
rect 523658 995607 523664 995619
rect 528400 995607 528406 995619
rect 528458 995607 528464 995659
rect 625648 995607 625654 995659
rect 625706 995647 625712 995659
rect 627856 995647 627862 995659
rect 625706 995619 627862 995647
rect 625706 995607 625712 995619
rect 627856 995607 627862 995619
rect 627914 995607 627920 995659
rect 132400 995533 132406 995585
rect 132458 995573 132464 995585
rect 144016 995573 144022 995585
rect 132458 995545 144022 995573
rect 132458 995533 132464 995545
rect 144016 995533 144022 995545
rect 144074 995533 144080 995585
rect 192496 995533 192502 995585
rect 192554 995573 192560 995585
rect 195376 995573 195382 995585
rect 192554 995545 195382 995573
rect 192554 995533 192560 995545
rect 195376 995533 195382 995545
rect 195434 995533 195440 995585
rect 295408 995533 295414 995585
rect 295466 995573 295472 995585
rect 298192 995573 298198 995585
rect 295466 995545 298198 995573
rect 295466 995533 295472 995545
rect 298192 995533 298198 995545
rect 298250 995533 298256 995585
rect 383056 995533 383062 995585
rect 383114 995573 383120 995585
rect 392368 995573 392374 995585
rect 383114 995545 392374 995573
rect 383114 995533 383120 995545
rect 392368 995533 392374 995545
rect 392426 995533 392432 995585
rect 472336 995533 472342 995585
rect 472394 995573 472400 995585
rect 476368 995573 476374 995585
rect 472394 995545 476374 995573
rect 472394 995533 472400 995545
rect 476368 995533 476374 995545
rect 476426 995533 476432 995585
rect 617776 995533 617782 995585
rect 617834 995573 617840 995585
rect 629200 995573 629206 995585
rect 617834 995545 629206 995573
rect 617834 995533 617840 995545
rect 629200 995533 629206 995545
rect 629258 995533 629264 995585
rect 82288 995459 82294 995511
rect 82346 995499 82352 995511
rect 92752 995499 92758 995511
rect 82346 995471 92758 995499
rect 82346 995459 82352 995471
rect 92752 995459 92758 995471
rect 92810 995459 92816 995511
rect 284368 995459 284374 995511
rect 284426 995499 284432 995511
rect 284426 995471 293630 995499
rect 284426 995459 284432 995471
rect 133072 995385 133078 995437
rect 133130 995425 133136 995437
rect 133130 995397 136190 995425
rect 133130 995385 133136 995397
rect 136162 995351 136190 995397
rect 136240 995385 136246 995437
rect 136298 995425 136304 995437
rect 143632 995425 143638 995437
rect 136298 995397 143638 995425
rect 136298 995385 136304 995397
rect 143632 995385 143638 995397
rect 143690 995385 143696 995437
rect 286768 995385 286774 995437
rect 286826 995425 286832 995437
rect 293602 995425 293630 995471
rect 293680 995459 293686 995511
rect 293738 995499 293744 995511
rect 298000 995499 298006 995511
rect 293738 995471 298006 995499
rect 293738 995459 293744 995471
rect 298000 995459 298006 995471
rect 298058 995459 298064 995511
rect 380464 995459 380470 995511
rect 380522 995499 380528 995511
rect 394864 995499 394870 995511
rect 380522 995471 394870 995499
rect 380522 995459 380528 995471
rect 394864 995459 394870 995471
rect 394922 995459 394928 995511
rect 466576 995459 466582 995511
rect 466634 995499 466640 995511
rect 482704 995499 482710 995511
rect 466634 995471 482710 995499
rect 466634 995459 466640 995471
rect 482704 995459 482710 995471
rect 482762 995459 482768 995511
rect 521776 995459 521782 995511
rect 521834 995499 521840 995511
rect 532816 995499 532822 995511
rect 521834 995471 532822 995499
rect 521834 995459 521840 995471
rect 532816 995459 532822 995471
rect 532874 995459 532880 995511
rect 298576 995425 298582 995437
rect 286826 995397 289598 995425
rect 293602 995397 298582 995425
rect 286826 995385 286832 995397
rect 146800 995351 146806 995363
rect 136162 995323 146806 995351
rect 146800 995311 146806 995323
rect 146858 995311 146864 995363
rect 133984 995237 133990 995289
rect 134042 995277 134048 995289
rect 143920 995277 143926 995289
rect 134042 995249 143926 995277
rect 134042 995237 134048 995249
rect 143920 995237 143926 995249
rect 143978 995237 143984 995289
rect 201712 995237 201718 995289
rect 201770 995277 201776 995289
rect 206512 995277 206518 995289
rect 201770 995249 206518 995277
rect 201770 995237 201776 995249
rect 206512 995237 206518 995249
rect 206570 995237 206576 995289
rect 82576 995163 82582 995215
rect 82634 995203 82640 995215
rect 134002 995203 134030 995237
rect 82634 995175 134030 995203
rect 82634 995163 82640 995175
rect 141232 995163 141238 995215
rect 141290 995203 141296 995215
rect 161200 995203 161206 995215
rect 141290 995175 161206 995203
rect 141290 995163 141296 995175
rect 161200 995163 161206 995175
rect 161258 995163 161264 995215
rect 181456 995163 181462 995215
rect 181514 995203 181520 995215
rect 201520 995203 201526 995215
rect 181514 995175 201526 995203
rect 181514 995163 181520 995175
rect 201520 995163 201526 995175
rect 201578 995163 201584 995215
rect 287152 995163 287158 995215
rect 287210 995203 287216 995215
rect 289456 995203 289462 995215
rect 287210 995175 289462 995203
rect 287210 995163 287216 995175
rect 289456 995163 289462 995175
rect 289514 995163 289520 995215
rect 289570 995203 289598 995397
rect 298576 995385 298582 995397
rect 298634 995385 298640 995437
rect 471952 995385 471958 995437
rect 472010 995425 472016 995437
rect 481360 995425 481366 995437
rect 472010 995397 481366 995425
rect 472010 995385 472016 995397
rect 481360 995385 481366 995397
rect 481418 995385 481424 995437
rect 523504 995385 523510 995437
rect 523562 995425 523568 995437
rect 531088 995425 531094 995437
rect 523562 995397 531094 995425
rect 523562 995385 523568 995397
rect 531088 995385 531094 995397
rect 531146 995385 531152 995437
rect 561712 995385 561718 995437
rect 561770 995425 561776 995437
rect 581680 995425 581686 995437
rect 561770 995397 581686 995425
rect 561770 995385 561776 995397
rect 581680 995385 581686 995397
rect 581738 995385 581744 995437
rect 521296 995311 521302 995363
rect 521354 995351 521360 995363
rect 640720 995351 640726 995363
rect 521354 995323 640726 995351
rect 521354 995311 521360 995323
rect 640720 995311 640726 995323
rect 640778 995311 640784 995363
rect 443536 995237 443542 995289
rect 443594 995277 443600 995289
rect 463600 995277 463606 995289
rect 443594 995249 463606 995277
rect 443594 995237 443600 995249
rect 463600 995237 463606 995249
rect 463658 995237 463664 995289
rect 515728 995237 515734 995289
rect 515786 995277 515792 995289
rect 642640 995277 642646 995289
rect 515786 995249 642646 995277
rect 515786 995237 515792 995249
rect 642640 995237 642646 995249
rect 642698 995237 642704 995289
rect 298672 995203 298678 995215
rect 289570 995175 298678 995203
rect 298672 995163 298678 995175
rect 298730 995163 298736 995215
rect 471664 995163 471670 995215
rect 471722 995203 471728 995215
rect 643408 995203 643414 995215
rect 471722 995175 643414 995203
rect 471722 995163 471728 995175
rect 643408 995163 643414 995175
rect 643466 995163 643472 995215
rect 69136 995089 69142 995141
rect 69194 995129 69200 995141
rect 302416 995129 302422 995141
rect 69194 995101 302422 995129
rect 69194 995089 69200 995101
rect 302416 995089 302422 995101
rect 302474 995089 302480 995141
rect 383152 995089 383158 995141
rect 383210 995129 383216 995141
rect 636496 995129 636502 995141
rect 383210 995101 636502 995129
rect 383210 995089 383216 995101
rect 636496 995089 636502 995101
rect 636554 995089 636560 995141
rect 118192 995015 118198 995067
rect 118250 995055 118256 995067
rect 561520 995055 561526 995067
rect 118250 995027 561526 995055
rect 118250 995015 118256 995027
rect 561520 995015 561526 995027
rect 561578 995015 561584 995067
rect 584752 995015 584758 995067
rect 584810 995055 584816 995067
rect 604720 995055 604726 995067
rect 584810 995027 604726 995055
rect 584810 995015 584816 995027
rect 604720 995015 604726 995027
rect 604778 995015 604784 995067
rect 247408 994941 247414 994993
rect 247466 994981 247472 994993
rect 259120 994981 259126 994993
rect 247466 994953 259126 994981
rect 247466 994941 247472 994953
rect 259120 994941 259126 994953
rect 259178 994941 259184 994993
rect 287824 994941 287830 994993
rect 287882 994981 287888 994993
rect 306448 994981 306454 994993
rect 287882 994953 306454 994981
rect 287882 994941 287888 994953
rect 306448 994941 306454 994953
rect 306506 994941 306512 994993
rect 290320 994793 290326 994845
rect 290378 994833 290384 994845
rect 311920 994833 311926 994845
rect 290378 994805 311926 994833
rect 290378 994793 290384 994805
rect 311920 994793 311926 994805
rect 311978 994793 311984 994845
rect 289264 994497 289270 994549
rect 289322 994537 289328 994549
rect 296656 994537 296662 994549
rect 289322 994509 296662 994537
rect 289322 994497 289328 994509
rect 296656 994497 296662 994509
rect 296714 994497 296720 994549
rect 131824 994127 131830 994179
rect 131882 994167 131888 994179
rect 158800 994167 158806 994179
rect 131882 994139 158806 994167
rect 131882 994127 131888 994139
rect 158800 994127 158806 994139
rect 158858 994127 158864 994179
rect 244816 994053 244822 994105
rect 244874 994093 244880 994105
rect 279280 994093 279286 994105
rect 244874 994065 279286 994093
rect 244874 994053 244880 994065
rect 279280 994053 279286 994065
rect 279338 994053 279344 994105
rect 234928 993905 234934 993957
rect 234986 993945 234992 993957
rect 253072 993945 253078 993957
rect 234986 993917 253078 993945
rect 234986 993905 234992 993917
rect 253072 993905 253078 993917
rect 253130 993905 253136 993957
rect 61840 993831 61846 993883
rect 61898 993871 61904 993883
rect 82576 993871 82582 993883
rect 61898 993843 82582 993871
rect 61898 993831 61904 993843
rect 82576 993831 82582 993843
rect 82634 993831 82640 993883
rect 238672 993831 238678 993883
rect 238730 993871 238736 993883
rect 260752 993871 260758 993883
rect 238730 993843 260758 993871
rect 238730 993831 238736 993843
rect 260752 993831 260758 993843
rect 260810 993831 260816 993883
rect 558160 993831 558166 993883
rect 558218 993871 558224 993883
rect 641008 993871 641014 993883
rect 558218 993843 641014 993871
rect 558218 993831 558224 993843
rect 641008 993831 641014 993843
rect 641066 993831 641072 993883
rect 77680 993757 77686 993809
rect 77738 993797 77744 993809
rect 100720 993797 100726 993809
rect 77738 993769 100726 993797
rect 77738 993757 77744 993769
rect 100720 993757 100726 993769
rect 100778 993757 100784 993809
rect 129328 993757 129334 993809
rect 129386 993797 129392 993809
rect 151696 993797 151702 993809
rect 129386 993769 151702 993797
rect 129386 993757 129392 993769
rect 151696 993757 151702 993769
rect 151754 993757 151760 993809
rect 180496 993757 180502 993809
rect 180554 993797 180560 993809
rect 201616 993797 201622 993809
rect 180554 993769 201622 993797
rect 180554 993757 180560 993769
rect 201616 993757 201622 993769
rect 201674 993757 201680 993809
rect 231472 993757 231478 993809
rect 231530 993797 231536 993809
rect 262384 993797 262390 993809
rect 231530 993769 262390 993797
rect 231530 993757 231536 993769
rect 262384 993757 262390 993769
rect 262442 993757 262448 993809
rect 78352 993683 78358 993735
rect 78410 993723 78416 993735
rect 109840 993723 109846 993735
rect 78410 993695 109846 993723
rect 78410 993683 78416 993695
rect 109840 993683 109846 993695
rect 109898 993683 109904 993735
rect 181360 993683 181366 993735
rect 181418 993723 181424 993735
rect 212656 993723 212662 993735
rect 181418 993695 212662 993723
rect 181418 993683 181424 993695
rect 212656 993683 212662 993695
rect 212714 993683 212720 993735
rect 232528 993683 232534 993735
rect 232586 993723 232592 993735
rect 264016 993723 264022 993735
rect 232586 993695 264022 993723
rect 232586 993683 232592 993695
rect 264016 993683 264022 993695
rect 264074 993683 264080 993735
rect 506608 993683 506614 993735
rect 506666 993723 506672 993735
rect 538960 993723 538966 993735
rect 506666 993695 538966 993723
rect 506666 993683 506672 993695
rect 538960 993683 538966 993695
rect 539018 993683 539024 993735
rect 77296 993609 77302 993661
rect 77354 993649 77360 993661
rect 108208 993649 108214 993661
rect 77354 993621 108214 993649
rect 77354 993609 77360 993621
rect 108208 993609 108214 993621
rect 108266 993609 108272 993661
rect 128464 993609 128470 993661
rect 128522 993649 128528 993661
rect 159568 993649 159574 993661
rect 128522 993621 159574 993649
rect 128522 993609 128528 993621
rect 159568 993609 159574 993621
rect 159626 993609 159632 993661
rect 179824 993609 179830 993661
rect 179882 993649 179888 993661
rect 211024 993649 211030 993661
rect 179882 993621 211030 993649
rect 179882 993609 179888 993621
rect 211024 993609 211030 993621
rect 211082 993609 211088 993661
rect 237424 993609 237430 993661
rect 237482 993649 237488 993661
rect 289264 993649 289270 993661
rect 237482 993621 289270 993649
rect 237482 993609 237488 993621
rect 289264 993609 289270 993621
rect 289322 993609 289328 993661
rect 362320 993609 362326 993661
rect 362378 993649 362384 993661
rect 398800 993649 398806 993661
rect 362378 993621 398806 993649
rect 362378 993609 362384 993621
rect 398800 993609 398806 993621
rect 398858 993609 398864 993661
rect 429712 993609 429718 993661
rect 429770 993649 429776 993661
rect 487792 993649 487798 993661
rect 429770 993621 487798 993649
rect 429770 993609 429776 993621
rect 487792 993609 487798 993621
rect 487850 993609 487856 993661
rect 531184 993609 531190 993661
rect 531242 993649 531248 993661
rect 633040 993649 633046 993661
rect 531242 993621 633046 993649
rect 531242 993609 531248 993621
rect 633040 993609 633046 993621
rect 633098 993609 633104 993661
rect 126640 993535 126646 993587
rect 126698 993575 126704 993587
rect 134608 993575 134614 993587
rect 126698 993547 134614 993575
rect 126698 993535 126704 993547
rect 134608 993535 134614 993547
rect 134666 993575 134672 993587
rect 186160 993575 186166 993587
rect 134666 993547 186166 993575
rect 134666 993535 134672 993547
rect 186160 993535 186166 993547
rect 186218 993575 186224 993587
rect 195760 993575 195766 993587
rect 186218 993547 195766 993575
rect 186218 993535 186224 993547
rect 195760 993535 195766 993547
rect 195818 993535 195824 993587
rect 279280 993535 279286 993587
rect 279338 993575 279344 993587
rect 288112 993575 288118 993587
rect 279338 993547 288118 993575
rect 279338 993535 279344 993547
rect 288112 993535 288118 993547
rect 288170 993575 288176 993587
rect 390160 993575 390166 993587
rect 288170 993547 390166 993575
rect 288170 993535 288176 993547
rect 390160 993535 390166 993547
rect 390218 993575 390224 993587
rect 479152 993575 479158 993587
rect 390218 993547 479158 993575
rect 390218 993535 390224 993547
rect 479152 993535 479158 993547
rect 479210 993575 479216 993587
rect 501040 993575 501046 993587
rect 479210 993547 501046 993575
rect 479210 993535 479216 993547
rect 501040 993535 501046 993547
rect 501098 993535 501104 993587
rect 636496 993535 636502 993587
rect 636554 993575 636560 993587
rect 643600 993575 643606 993587
rect 636554 993547 643606 993575
rect 636554 993535 636560 993547
rect 643600 993535 643606 993547
rect 643658 993535 643664 993587
rect 642640 993461 642646 993513
rect 642698 993501 642704 993513
rect 649456 993501 649462 993513
rect 642698 993473 649462 993501
rect 642698 993461 642704 993473
rect 649456 993461 649462 993473
rect 649514 993461 649520 993513
rect 331216 992573 331222 992625
rect 331274 992613 331280 992625
rect 332560 992613 332566 992625
rect 331274 992585 332566 992613
rect 331274 992573 331280 992585
rect 332560 992573 332566 992585
rect 332618 992573 332624 992625
rect 640720 990723 640726 990775
rect 640778 990763 640784 990775
rect 640778 990735 642302 990763
rect 640778 990723 640784 990735
rect 642274 990689 642302 990735
rect 645136 990689 645142 990701
rect 642274 990661 645142 990689
rect 645136 990649 645142 990661
rect 645194 990649 645200 990701
rect 89584 990501 89590 990553
rect 89642 990541 89648 990553
rect 93712 990541 93718 990553
rect 89642 990513 93718 990541
rect 89642 990501 89648 990513
rect 93712 990501 93718 990513
rect 93770 990501 93776 990553
rect 219472 990501 219478 990553
rect 219530 990541 219536 990553
rect 221776 990541 221782 990553
rect 219530 990513 221782 990541
rect 219530 990501 219536 990513
rect 221776 990501 221782 990513
rect 221834 990501 221840 990553
rect 444496 990501 444502 990553
rect 444554 990541 444560 990553
rect 462736 990541 462742 990553
rect 444554 990513 462742 990541
rect 444554 990501 444560 990513
rect 462736 990501 462742 990513
rect 462794 990501 462800 990553
rect 521392 989465 521398 989517
rect 521450 989505 521456 989517
rect 521450 989477 538526 989505
rect 521450 989465 521456 989477
rect 374416 989391 374422 989443
rect 374474 989431 374480 989443
rect 397840 989431 397846 989443
rect 374474 989403 397846 989431
rect 374474 989391 374480 989403
rect 397840 989391 397846 989403
rect 397898 989391 397904 989443
rect 154480 989317 154486 989369
rect 154538 989357 154544 989369
rect 163984 989357 163990 989369
rect 154538 989329 163990 989357
rect 154538 989317 154544 989329
rect 163984 989317 163990 989329
rect 164042 989317 164048 989369
rect 222928 989317 222934 989369
rect 222986 989357 222992 989369
rect 235600 989357 235606 989369
rect 222986 989329 235606 989357
rect 222986 989317 222992 989329
rect 235600 989317 235606 989329
rect 235658 989317 235664 989369
rect 273616 989317 273622 989369
rect 273674 989357 273680 989369
rect 284272 989357 284278 989369
rect 273674 989329 284278 989357
rect 273674 989317 273680 989329
rect 284272 989317 284278 989329
rect 284330 989317 284336 989369
rect 328240 989317 328246 989369
rect 328298 989357 328304 989369
rect 349168 989357 349174 989369
rect 328298 989329 349174 989357
rect 328298 989317 328304 989329
rect 349168 989317 349174 989329
rect 349226 989317 349232 989369
rect 377296 989317 377302 989369
rect 377354 989357 377360 989369
rect 414064 989357 414070 989369
rect 377354 989329 414070 989357
rect 377354 989317 377360 989329
rect 414064 989317 414070 989329
rect 414122 989317 414128 989369
rect 446224 989317 446230 989369
rect 446282 989357 446288 989369
rect 478960 989357 478966 989369
rect 446282 989329 478966 989357
rect 446282 989317 446288 989329
rect 478960 989317 478966 989329
rect 479018 989317 479024 989369
rect 518512 989317 518518 989369
rect 518570 989357 518576 989369
rect 527632 989357 527638 989369
rect 518570 989329 527638 989357
rect 518570 989317 518576 989329
rect 527632 989317 527638 989329
rect 527690 989317 527696 989369
rect 538498 989357 538526 989477
rect 570256 989465 570262 989517
rect 570314 989505 570320 989517
rect 592432 989505 592438 989517
rect 570314 989477 592438 989505
rect 570314 989465 570320 989477
rect 592432 989465 592438 989477
rect 592490 989465 592496 989517
rect 573136 989391 573142 989443
rect 573194 989431 573200 989443
rect 608752 989431 608758 989443
rect 573194 989403 608758 989431
rect 573194 989391 573200 989403
rect 608752 989391 608758 989403
rect 608810 989391 608816 989443
rect 543760 989357 543766 989369
rect 538498 989329 543766 989357
rect 543760 989317 543766 989329
rect 543818 989317 543824 989369
rect 570352 989317 570358 989369
rect 570410 989357 570416 989369
rect 624976 989357 624982 989369
rect 570410 989329 624982 989357
rect 570410 989317 570416 989329
rect 624976 989317 624982 989329
rect 625034 989317 625040 989369
rect 73456 989243 73462 989295
rect 73514 989283 73520 989295
rect 92944 989283 92950 989295
rect 73514 989255 92950 989283
rect 73514 989243 73520 989255
rect 92944 989243 92950 989255
rect 93002 989243 93008 989295
rect 138256 989243 138262 989295
rect 138314 989283 138320 989295
rect 164080 989283 164086 989295
rect 138314 989255 164086 989283
rect 138314 989243 138320 989255
rect 164080 989243 164086 989255
rect 164138 989243 164144 989295
rect 273712 989243 273718 989295
rect 273770 989283 273776 989295
rect 300496 989283 300502 989295
rect 273770 989255 300502 989283
rect 273770 989243 273776 989255
rect 300496 989243 300502 989255
rect 300554 989243 300560 989295
rect 325264 989243 325270 989295
rect 325322 989283 325328 989295
rect 365392 989283 365398 989295
rect 325322 989255 365398 989283
rect 325322 989243 325328 989255
rect 365392 989243 365398 989255
rect 365450 989243 365456 989295
rect 374512 989243 374518 989295
rect 374570 989283 374576 989295
rect 430288 989283 430294 989295
rect 374570 989255 430294 989283
rect 374570 989243 374576 989255
rect 430288 989243 430294 989255
rect 430346 989243 430352 989295
rect 440752 989243 440758 989295
rect 440810 989283 440816 989295
rect 495184 989283 495190 989295
rect 440810 989255 495190 989283
rect 440810 989243 440816 989255
rect 495184 989243 495190 989255
rect 495242 989243 495248 989295
rect 518704 989243 518710 989295
rect 518762 989283 518768 989295
rect 560080 989283 560086 989295
rect 518762 989255 560086 989283
rect 518762 989243 518768 989255
rect 560080 989243 560086 989255
rect 560138 989243 560144 989295
rect 567664 989243 567670 989295
rect 567722 989283 567728 989295
rect 658000 989283 658006 989295
rect 567722 989255 658006 989283
rect 567722 989243 567728 989255
rect 658000 989243 658006 989255
rect 658058 989243 658064 989295
rect 203152 988799 203158 988851
rect 203210 988839 203216 988851
rect 213040 988839 213046 988851
rect 203210 988811 213046 988839
rect 203210 988799 203216 988811
rect 213040 988799 213046 988811
rect 213098 988799 213104 988851
rect 288016 988651 288022 988703
rect 288074 988691 288080 988703
rect 299152 988691 299158 988703
rect 288074 988663 299158 988691
rect 288074 988651 288080 988663
rect 299152 988651 299158 988663
rect 299210 988651 299216 988703
rect 47632 988281 47638 988333
rect 47690 988321 47696 988333
rect 122032 988321 122038 988333
rect 47690 988293 122038 988321
rect 47690 988281 47696 988293
rect 122032 988281 122038 988293
rect 122090 988281 122096 988333
rect 44752 988207 44758 988259
rect 44810 988247 44816 988259
rect 186928 988247 186934 988259
rect 44810 988219 186934 988247
rect 44810 988207 44816 988219
rect 186928 988207 186934 988219
rect 186986 988207 186992 988259
rect 561520 988207 561526 988259
rect 561578 988247 561584 988259
rect 576304 988247 576310 988259
rect 561578 988219 576310 988247
rect 561578 988207 561584 988219
rect 576304 988207 576310 988219
rect 576362 988207 576368 988259
rect 44848 988133 44854 988185
rect 44906 988173 44912 988185
rect 251824 988173 251830 988185
rect 44906 988145 251830 988173
rect 44906 988133 44912 988145
rect 251824 988133 251830 988145
rect 251882 988133 251888 988185
rect 44944 988059 44950 988111
rect 45002 988099 45008 988111
rect 316720 988099 316726 988111
rect 45002 988071 316726 988099
rect 45002 988059 45008 988071
rect 316720 988059 316726 988071
rect 316778 988059 316784 988111
rect 45040 987985 45046 988037
rect 45098 988025 45104 988037
rect 381616 988025 381622 988037
rect 45098 987997 381622 988025
rect 45098 987985 45104 987997
rect 381616 987985 381622 987997
rect 381674 987985 381680 988037
rect 45136 987911 45142 987963
rect 45194 987951 45200 987963
rect 446512 987951 446518 987963
rect 45194 987923 446518 987951
rect 45194 987911 45200 987923
rect 446512 987911 446518 987923
rect 446570 987911 446576 987963
rect 43120 987837 43126 987889
rect 43178 987877 43184 987889
rect 511408 987877 511414 987889
rect 43178 987849 511414 987877
rect 43178 987837 43184 987849
rect 511408 987837 511414 987849
rect 511466 987837 511472 987889
rect 244720 987763 244726 987815
rect 244778 987803 244784 987815
rect 247504 987803 247510 987815
rect 244778 987775 247510 987803
rect 244778 987763 244784 987775
rect 247504 987763 247510 987775
rect 247562 987763 247568 987815
rect 640528 987763 640534 987815
rect 640586 987803 640592 987815
rect 649552 987803 649558 987815
rect 640586 987775 649558 987803
rect 640586 987763 640592 987775
rect 649552 987763 649558 987775
rect 649610 987763 649616 987815
rect 643600 987689 643606 987741
rect 643658 987729 643664 987741
rect 650128 987729 650134 987741
rect 643658 987701 650134 987729
rect 643658 987689 643664 987701
rect 650128 987689 650134 987701
rect 650186 987689 650192 987741
rect 643408 987615 643414 987667
rect 643466 987655 643472 987667
rect 649648 987655 649654 987667
rect 643466 987627 649654 987655
rect 643466 987615 643472 987627
rect 649648 987615 649654 987627
rect 649706 987615 649712 987667
rect 640912 987541 640918 987593
rect 640970 987581 640976 987593
rect 650032 987581 650038 987593
rect 640970 987553 650038 987581
rect 640970 987541 640976 987553
rect 650032 987541 650038 987553
rect 650090 987541 650096 987593
rect 47920 986653 47926 986705
rect 47978 986693 47984 986705
rect 115312 986693 115318 986705
rect 47978 986665 115318 986693
rect 47978 986653 47984 986665
rect 115312 986653 115318 986665
rect 115370 986653 115376 986705
rect 47728 986579 47734 986631
rect 47786 986619 47792 986631
rect 115216 986619 115222 986631
rect 47786 986591 115222 986619
rect 47786 986579 47792 986591
rect 115216 986579 115222 986591
rect 115274 986579 115280 986631
rect 629200 986579 629206 986631
rect 629258 986619 629264 986631
rect 649744 986619 649750 986631
rect 629258 986591 649750 986619
rect 629258 986579 629264 986591
rect 649744 986579 649750 986591
rect 649802 986579 649808 986631
rect 47440 986505 47446 986557
rect 47498 986545 47504 986557
rect 118096 986545 118102 986557
rect 47498 986517 118102 986545
rect 47498 986505 47504 986517
rect 118096 986505 118102 986517
rect 118154 986505 118160 986557
rect 567376 986505 567382 986557
rect 567434 986545 567440 986557
rect 660880 986545 660886 986557
rect 567434 986517 660886 986545
rect 567434 986505 567440 986517
rect 660880 986505 660886 986517
rect 660938 986505 660944 986557
rect 63280 986431 63286 986483
rect 63338 986471 63344 986483
rect 145264 986471 145270 986483
rect 63338 986443 145270 986471
rect 63338 986431 63344 986443
rect 145264 986431 145270 986443
rect 145322 986431 145328 986483
rect 567472 986431 567478 986483
rect 567530 986471 567536 986483
rect 660976 986471 660982 986483
rect 567530 986443 660982 986471
rect 567530 986431 567536 986443
rect 660976 986431 660982 986443
rect 661034 986431 661040 986483
rect 65200 986357 65206 986409
rect 65258 986397 65264 986409
rect 195088 986397 195094 986409
rect 65258 986369 195094 986397
rect 65258 986357 65264 986369
rect 195088 986357 195094 986369
rect 195146 986357 195152 986409
rect 544240 986357 544246 986409
rect 544298 986397 544304 986409
rect 650992 986397 650998 986409
rect 544298 986369 650998 986397
rect 544298 986357 544304 986369
rect 650992 986357 650998 986369
rect 651050 986357 651056 986409
rect 277936 985099 277942 985151
rect 277994 985139 278000 985151
rect 288016 985139 288022 985151
rect 277994 985111 288022 985139
rect 277994 985099 278000 985111
rect 288016 985099 288022 985111
rect 288074 985099 288080 985151
rect 65104 984951 65110 985003
rect 65162 984991 65168 985003
rect 94960 984991 94966 985003
rect 65162 984963 94966 984991
rect 65162 984951 65168 984963
rect 94960 984951 94966 984963
rect 95018 984951 95024 985003
rect 645136 984877 645142 984929
rect 645194 984917 645200 984929
rect 649936 984917 649942 984929
rect 645194 984889 649942 984917
rect 645194 984877 645200 984889
rect 649936 984877 649942 984889
rect 649994 984877 650000 984929
rect 64816 984137 64822 984189
rect 64874 984177 64880 984189
rect 69040 984177 69046 984189
rect 64874 984149 69046 984177
rect 64874 984137 64880 984149
rect 69040 984137 69046 984149
rect 69098 984137 69104 984189
rect 632368 983619 632374 983671
rect 632426 983659 632432 983671
rect 674512 983659 674518 983671
rect 632426 983631 674518 983659
rect 632426 983619 632432 983631
rect 674512 983619 674518 983631
rect 674570 983619 674576 983671
rect 64912 983545 64918 983597
rect 64970 983585 64976 983597
rect 244720 983585 244726 983597
rect 64970 983557 244726 983585
rect 64970 983545 64976 983557
rect 244720 983545 244726 983557
rect 244778 983545 244784 983597
rect 633040 983545 633046 983597
rect 633098 983585 633104 983597
rect 674320 983585 674326 983597
rect 633098 983557 674326 983585
rect 633098 983545 633104 983557
rect 674320 983545 674326 983557
rect 674378 983545 674384 983597
rect 65008 983471 65014 983523
rect 65066 983511 65072 983523
rect 277936 983511 277942 983523
rect 65066 983483 277942 983511
rect 65066 983471 65072 983483
rect 277936 983471 277942 983483
rect 277994 983471 278000 983523
rect 429136 983471 429142 983523
rect 429194 983511 429200 983523
rect 649360 983511 649366 983523
rect 429194 983483 649366 983511
rect 429194 983471 429200 983483
rect 649360 983471 649366 983483
rect 649418 983471 649424 983523
rect 50512 973481 50518 973533
rect 50570 973521 50576 973533
rect 59440 973521 59446 973533
rect 50570 973493 59446 973521
rect 50570 973481 50576 973493
rect 59440 973481 59446 973493
rect 59498 973481 59504 973533
rect 42160 967265 42166 967317
rect 42218 967305 42224 967317
rect 43120 967305 43126 967317
rect 42218 967277 43126 967305
rect 42218 967265 42224 967277
rect 43120 967265 43126 967277
rect 43178 967265 43184 967317
rect 42160 960975 42166 961027
rect 42218 961015 42224 961027
rect 42448 961015 42454 961027
rect 42218 960987 42454 961015
rect 42218 960975 42224 960987
rect 42448 960975 42454 960987
rect 42506 960975 42512 961027
rect 46096 959051 46102 959103
rect 46154 959091 46160 959103
rect 59536 959091 59542 959103
rect 46154 959063 59542 959091
rect 46154 959051 46160 959063
rect 59536 959051 59542 959063
rect 59594 959051 59600 959103
rect 675088 958163 675094 958215
rect 675146 958203 675152 958215
rect 675376 958203 675382 958215
rect 675146 958175 675382 958203
rect 675146 958163 675152 958175
rect 675376 958163 675382 958175
rect 675434 958163 675440 958215
rect 675184 956979 675190 957031
rect 675242 957019 675248 957031
rect 675472 957019 675478 957031
rect 675242 956991 675478 957019
rect 675242 956979 675248 956991
rect 675472 956979 675478 956991
rect 675530 956979 675536 957031
rect 42064 955203 42070 955255
rect 42122 955243 42128 955255
rect 42832 955243 42838 955255
rect 42122 955215 42838 955243
rect 42122 955203 42128 955215
rect 42832 955203 42838 955215
rect 42890 955203 42896 955255
rect 669520 954685 669526 954737
rect 669578 954725 669584 954737
rect 675376 954725 675382 954737
rect 669578 954697 675382 954725
rect 669578 954685 669584 954697
rect 675376 954685 675382 954697
rect 675434 954685 675440 954737
rect 41776 954611 41782 954663
rect 41834 954611 41840 954663
rect 41794 954441 41822 954611
rect 41776 954389 41782 954441
rect 41834 954389 41840 954441
rect 673936 953945 673942 953997
rect 673994 953985 674000 953997
rect 675472 953985 675478 953997
rect 673994 953957 675478 953985
rect 673994 953945 674000 953957
rect 675472 953945 675478 953957
rect 675530 953945 675536 953997
rect 37360 952169 37366 952221
rect 37418 952209 37424 952221
rect 41776 952209 41782 952221
rect 37418 952181 41782 952209
rect 37418 952169 37424 952181
rect 41776 952169 41782 952181
rect 41834 952169 41840 952221
rect 674032 952021 674038 952073
rect 674090 952061 674096 952073
rect 675472 952061 675478 952073
rect 674090 952033 675478 952061
rect 674090 952021 674096 952033
rect 675472 952021 675478 952033
rect 675530 952021 675536 952073
rect 42352 948395 42358 948447
rect 42410 948435 42416 948447
rect 53200 948435 53206 948447
rect 42410 948407 53206 948435
rect 42410 948395 42416 948407
rect 53200 948395 53206 948407
rect 53258 948395 53264 948447
rect 42640 947877 42646 947929
rect 42698 947917 42704 947929
rect 46096 947917 46102 947929
rect 42698 947889 46102 947917
rect 42698 947877 42704 947889
rect 46096 947877 46102 947889
rect 46154 947877 46160 947929
rect 42448 947433 42454 947485
rect 42506 947473 42512 947485
rect 57808 947473 57814 947485
rect 42506 947445 57814 947473
rect 42506 947433 42512 947445
rect 57808 947433 57814 947445
rect 57866 947433 57872 947485
rect 655216 944843 655222 944895
rect 655274 944883 655280 944895
rect 674512 944883 674518 944895
rect 655274 944855 674518 944883
rect 655274 944843 655280 944855
rect 674512 944843 674518 944855
rect 674570 944843 674576 944895
rect 655120 944621 655126 944673
rect 655178 944661 655184 944673
rect 674512 944661 674518 944673
rect 655178 944633 674518 944661
rect 655178 944621 655184 944633
rect 674512 944621 674518 944633
rect 674570 944621 674576 944673
rect 658000 942031 658006 942083
rect 658058 942071 658064 942083
rect 674512 942071 674518 942083
rect 658058 942043 674518 942071
rect 658058 942031 658064 942043
rect 674512 942031 674518 942043
rect 674570 942031 674576 942083
rect 660976 941957 660982 942009
rect 661034 941997 661040 942009
rect 674416 941997 674422 942009
rect 661034 941969 674422 941997
rect 661034 941957 661040 941969
rect 674416 941957 674422 941969
rect 674474 941957 674480 942009
rect 654448 941883 654454 941935
rect 654506 941923 654512 941935
rect 674896 941923 674902 941935
rect 654506 941895 674902 941923
rect 654506 941883 654512 941895
rect 674896 941883 674902 941895
rect 674954 941883 674960 941935
rect 660880 941143 660886 941195
rect 660938 941183 660944 941195
rect 674416 941183 674422 941195
rect 660938 941155 674422 941183
rect 660938 941143 660944 941155
rect 674416 941143 674422 941155
rect 674474 941143 674480 941195
rect 674032 938997 674038 939049
rect 674090 939037 674096 939049
rect 676816 939037 676822 939049
rect 674090 939009 676822 939037
rect 674090 938997 674096 939009
rect 676816 938997 676822 939009
rect 676874 938997 676880 939049
rect 53200 933077 53206 933129
rect 53258 933117 53264 933129
rect 59536 933117 59542 933129
rect 53258 933089 59542 933117
rect 53258 933077 53264 933089
rect 59536 933077 59542 933089
rect 59594 933077 59600 933129
rect 42352 930931 42358 930983
rect 42410 930971 42416 930983
rect 44656 930971 44662 930983
rect 42410 930943 44662 930971
rect 42410 930931 42416 930943
rect 44656 930931 44662 930943
rect 44714 930931 44720 930983
rect 654448 927453 654454 927505
rect 654506 927493 654512 927505
rect 666736 927493 666742 927505
rect 654506 927465 666742 927493
rect 654506 927453 654512 927465
rect 666736 927453 666742 927465
rect 666794 927453 666800 927505
rect 40048 927379 40054 927431
rect 40106 927419 40112 927431
rect 40240 927419 40246 927431
rect 40106 927391 40246 927419
rect 40106 927379 40112 927391
rect 40240 927379 40246 927391
rect 40298 927379 40304 927431
rect 649552 927379 649558 927431
rect 649610 927419 649616 927431
rect 679792 927419 679798 927431
rect 649610 927391 679798 927419
rect 649610 927379 649616 927391
rect 679792 927379 679798 927391
rect 679850 927379 679856 927431
rect 53392 915835 53398 915887
rect 53450 915875 53456 915887
rect 59536 915875 59542 915887
rect 53450 915847 59542 915875
rect 53450 915835 53456 915847
rect 59536 915835 59542 915847
rect 59594 915835 59600 915887
rect 653968 915835 653974 915887
rect 654026 915875 654032 915887
rect 660976 915875 660982 915887
rect 654026 915847 660982 915875
rect 654026 915835 654032 915847
rect 660976 915835 660982 915847
rect 661034 915835 661040 915887
rect 654448 904365 654454 904417
rect 654506 904405 654512 904417
rect 663952 904405 663958 904417
rect 654506 904377 663958 904405
rect 654506 904365 654512 904377
rect 663952 904365 663958 904377
rect 664010 904365 664016 904417
rect 50320 901479 50326 901531
rect 50378 901519 50384 901531
rect 59536 901519 59542 901531
rect 50378 901491 59542 901519
rect 50378 901479 50384 901491
rect 59536 901479 59542 901491
rect 59594 901479 59600 901531
rect 39952 892821 39958 892873
rect 40010 892861 40016 892873
rect 40144 892861 40150 892873
rect 40010 892833 40150 892861
rect 40010 892821 40016 892833
rect 40144 892821 40150 892833
rect 40202 892821 40208 892873
rect 53200 887123 53206 887175
rect 53258 887163 53264 887175
rect 59536 887163 59542 887175
rect 53258 887135 59542 887163
rect 53258 887123 53264 887135
rect 59536 887123 59542 887135
rect 59594 887123 59600 887175
rect 653968 881277 653974 881329
rect 654026 881317 654032 881329
rect 660880 881317 660886 881329
rect 654026 881289 660886 881317
rect 654026 881277 654032 881289
rect 660880 881277 660886 881289
rect 660938 881277 660944 881329
rect 673168 872841 673174 872893
rect 673226 872881 673232 872893
rect 675376 872881 675382 872893
rect 673226 872853 675382 872881
rect 673226 872841 673232 872853
rect 675376 872841 675382 872853
rect 675434 872841 675440 872893
rect 47536 872619 47542 872671
rect 47594 872659 47600 872671
rect 59536 872659 59542 872671
rect 47594 872631 59542 872659
rect 47594 872619 47600 872631
rect 59536 872619 59542 872631
rect 59594 872619 59600 872671
rect 673360 872101 673366 872153
rect 673418 872141 673424 872153
rect 675472 872141 675478 872153
rect 673418 872113 675478 872141
rect 673418 872101 673424 872113
rect 675472 872101 675478 872113
rect 675530 872101 675536 872153
rect 674032 871657 674038 871709
rect 674090 871697 674096 871709
rect 675088 871697 675094 871709
rect 674090 871669 675094 871697
rect 674090 871657 674096 871669
rect 675088 871657 675094 871669
rect 675146 871697 675152 871709
rect 675376 871697 675382 871709
rect 675146 871669 675382 871697
rect 675146 871657 675152 871669
rect 675376 871657 675382 871669
rect 675434 871657 675440 871709
rect 674224 871435 674230 871487
rect 674282 871475 674288 871487
rect 675184 871475 675190 871487
rect 674282 871447 675190 871475
rect 674282 871435 674288 871447
rect 675184 871435 675190 871447
rect 675242 871475 675248 871487
rect 675376 871475 675382 871487
rect 675242 871447 675382 871475
rect 675242 871435 675248 871447
rect 675376 871435 675382 871447
rect 675434 871435 675440 871487
rect 654448 869807 654454 869859
rect 654506 869847 654512 869859
rect 663760 869847 663766 869859
rect 654506 869819 663766 869847
rect 654506 869807 654512 869819
rect 663760 869807 663766 869819
rect 663818 869807 663824 869859
rect 673072 869141 673078 869193
rect 673130 869181 673136 869193
rect 675472 869181 675478 869193
rect 673130 869153 675478 869181
rect 673130 869141 673136 869153
rect 675472 869141 675478 869153
rect 675530 869141 675536 869193
rect 674512 868327 674518 868379
rect 674570 868367 674576 868379
rect 675376 868367 675382 868379
rect 674570 868339 675382 868367
rect 674570 868327 674576 868339
rect 675376 868327 675382 868339
rect 675434 868327 675440 868379
rect 673264 867809 673270 867861
rect 673322 867849 673328 867861
rect 675376 867849 675382 867861
rect 673322 867821 675382 867849
rect 673322 867809 673328 867821
rect 675376 867809 675382 867821
rect 675434 867809 675440 867861
rect 674128 866477 674134 866529
rect 674186 866517 674192 866529
rect 675376 866517 675382 866529
rect 674186 866489 675382 866517
rect 674186 866477 674192 866489
rect 675376 866477 675382 866489
rect 675434 866477 675440 866529
rect 666640 865293 666646 865345
rect 666698 865333 666704 865345
rect 675376 865333 675382 865345
rect 666698 865305 675382 865333
rect 666698 865293 666704 865305
rect 675376 865293 675382 865305
rect 675434 865293 675440 865345
rect 40048 863961 40054 864013
rect 40106 864001 40112 864013
rect 40240 864001 40246 864013
rect 40106 863973 40246 864001
rect 40106 863961 40112 863973
rect 40240 863961 40246 863973
rect 40298 863961 40304 864013
rect 47440 858263 47446 858315
rect 47498 858303 47504 858315
rect 58576 858303 58582 858315
rect 47498 858275 58582 858303
rect 47498 858263 47504 858275
rect 58576 858263 58582 858275
rect 58634 858263 58640 858315
rect 654160 858263 654166 858315
rect 654218 858303 654224 858315
rect 661072 858303 661078 858315
rect 654218 858275 661078 858303
rect 654218 858263 654224 858275
rect 661072 858263 661078 858275
rect 661130 858263 661136 858315
rect 53296 843833 53302 843885
rect 53354 843873 53360 843885
rect 59536 843873 59542 843885
rect 53354 843845 59542 843873
rect 53354 843833 53360 843845
rect 59536 843833 59542 843845
rect 59594 843833 59600 843885
rect 653968 835175 653974 835227
rect 654026 835215 654032 835227
rect 669712 835215 669718 835227
rect 654026 835187 669718 835215
rect 654026 835175 654032 835187
rect 669712 835175 669718 835187
rect 669770 835175 669776 835227
rect 40240 832363 40246 832415
rect 40298 832363 40304 832415
rect 40048 832289 40054 832341
rect 40106 832329 40112 832341
rect 40258 832329 40286 832363
rect 40106 832301 40286 832329
rect 40106 832289 40112 832301
rect 47728 829477 47734 829529
rect 47786 829517 47792 829529
rect 59536 829517 59542 829529
rect 47786 829489 59542 829517
rect 47786 829477 47792 829489
rect 59536 829477 59542 829489
rect 59594 829477 59600 829529
rect 40048 826591 40054 826643
rect 40106 826631 40112 826643
rect 40240 826631 40246 826643
rect 40106 826603 40246 826631
rect 40106 826591 40112 826603
rect 40240 826591 40246 826603
rect 40298 826591 40304 826643
rect 42160 823853 42166 823905
rect 42218 823893 42224 823905
rect 53200 823893 53206 823905
rect 42218 823865 53206 823893
rect 42218 823853 42224 823865
rect 53200 823853 53206 823865
rect 53258 823853 53264 823905
rect 653968 823705 653974 823757
rect 654026 823745 654032 823757
rect 672496 823745 672502 823757
rect 654026 823717 672502 823745
rect 654026 823705 654032 823717
rect 672496 823705 672502 823717
rect 672554 823705 672560 823757
rect 42160 823113 42166 823165
rect 42218 823153 42224 823165
rect 47536 823153 47542 823165
rect 42218 823125 47542 823153
rect 42218 823113 42224 823125
rect 47536 823113 47542 823125
rect 47594 823113 47600 823165
rect 42160 822225 42166 822277
rect 42218 822265 42224 822277
rect 50320 822265 50326 822277
rect 42218 822237 50326 822265
rect 42218 822225 42224 822237
rect 50320 822225 50326 822237
rect 50378 822225 50384 822277
rect 50416 815047 50422 815099
rect 50474 815087 50480 815099
rect 59536 815087 59542 815099
rect 50474 815059 59542 815087
rect 50474 815047 50480 815059
rect 59536 815047 59542 815059
rect 59594 815047 59600 815099
rect 654448 812161 654454 812213
rect 654506 812201 654512 812213
rect 664048 812201 664054 812213
rect 654506 812173 664054 812201
rect 654506 812161 654512 812173
rect 664048 812161 664054 812173
rect 664106 812161 664112 812213
rect 42160 810459 42166 810511
rect 42218 810499 42224 810511
rect 43024 810499 43030 810511
rect 42218 810471 43030 810499
rect 42218 810459 42224 810471
rect 43024 810459 43030 810471
rect 43082 810459 43088 810511
rect 42448 807055 42454 807107
rect 42506 807095 42512 807107
rect 42832 807095 42838 807107
rect 42506 807067 42838 807095
rect 42506 807055 42512 807067
rect 42832 807055 42838 807067
rect 42890 807055 42896 807107
rect 42832 805427 42838 805479
rect 42890 805467 42896 805479
rect 53200 805467 53206 805479
rect 42890 805439 53206 805467
rect 42890 805427 42896 805439
rect 53200 805427 53206 805439
rect 53258 805427 53264 805479
rect 40144 803429 40150 803481
rect 40202 803469 40208 803481
rect 42832 803469 42838 803481
rect 40202 803441 42838 803469
rect 40202 803429 40208 803441
rect 42832 803429 42838 803441
rect 42890 803429 42896 803481
rect 41968 802023 41974 802075
rect 42026 802063 42032 802075
rect 42448 802063 42454 802075
rect 42026 802035 42454 802063
rect 42026 802023 42032 802035
rect 42448 802023 42454 802035
rect 42506 802023 42512 802075
rect 43408 800617 43414 800669
rect 43466 800657 43472 800669
rect 45136 800657 45142 800669
rect 43466 800629 45142 800657
rect 43466 800617 43472 800629
rect 45136 800617 45142 800629
rect 45194 800617 45200 800669
rect 50320 800617 50326 800669
rect 50378 800657 50384 800669
rect 59536 800657 59542 800669
rect 50378 800629 59542 800657
rect 50378 800617 50384 800629
rect 59536 800617 59542 800629
rect 59594 800617 59600 800669
rect 41488 800543 41494 800595
rect 41546 800583 41552 800595
rect 43600 800583 43606 800595
rect 41546 800555 43606 800583
rect 41546 800543 41552 800555
rect 43600 800543 43606 800555
rect 43658 800543 43664 800595
rect 41584 800469 41590 800521
rect 41642 800509 41648 800521
rect 43504 800509 43510 800521
rect 41642 800481 43510 800509
rect 41642 800469 41648 800481
rect 43504 800469 43510 800481
rect 43562 800469 43568 800521
rect 41872 800173 41878 800225
rect 41930 800173 41936 800225
rect 42160 800173 42166 800225
rect 42218 800213 42224 800225
rect 43312 800213 43318 800225
rect 42218 800185 43318 800213
rect 42218 800173 42224 800185
rect 43312 800173 43318 800185
rect 43370 800173 43376 800225
rect 41890 800003 41918 800173
rect 41872 799951 41878 800003
rect 41930 799951 41936 800003
rect 43024 798471 43030 798523
rect 43082 798471 43088 798523
rect 42832 798323 42838 798375
rect 42890 798323 42896 798375
rect 42160 798101 42166 798153
rect 42218 798141 42224 798153
rect 42850 798141 42878 798323
rect 42218 798113 42878 798141
rect 42218 798101 42224 798113
rect 42736 798027 42742 798079
rect 42794 798067 42800 798079
rect 43042 798067 43070 798471
rect 42794 798039 43070 798067
rect 42794 798027 42800 798039
rect 42064 797287 42070 797339
rect 42122 797327 42128 797339
rect 43408 797327 43414 797339
rect 42122 797299 43414 797327
rect 42122 797287 42128 797299
rect 43408 797287 43414 797299
rect 43466 797287 43472 797339
rect 42160 796251 42166 796303
rect 42218 796291 42224 796303
rect 42736 796291 42742 796303
rect 42218 796263 42742 796291
rect 42218 796251 42224 796263
rect 42736 796251 42742 796263
rect 42794 796251 42800 796303
rect 42736 796103 42742 796155
rect 42794 796143 42800 796155
rect 43312 796143 43318 796155
rect 42794 796115 43318 796143
rect 42794 796103 42800 796115
rect 43312 796103 43318 796115
rect 43370 796103 43376 796155
rect 42160 794993 42166 795045
rect 42218 795033 42224 795045
rect 43120 795033 43126 795045
rect 42218 795005 43126 795033
rect 42218 794993 42224 795005
rect 43120 794993 43126 795005
rect 43178 794993 43184 795045
rect 43120 794845 43126 794897
rect 43178 794885 43184 794897
rect 43504 794885 43510 794897
rect 43178 794857 43510 794885
rect 43178 794845 43184 794857
rect 43504 794845 43510 794857
rect 43562 794845 43568 794897
rect 42160 792995 42166 793047
rect 42218 793035 42224 793047
rect 42736 793035 42742 793047
rect 42218 793007 42742 793035
rect 42218 792995 42224 793007
rect 42736 792995 42742 793007
rect 42794 792995 42800 793047
rect 42736 792847 42742 792899
rect 42794 792887 42800 792899
rect 43120 792887 43126 792899
rect 42794 792859 43126 792887
rect 42794 792847 42800 792859
rect 43120 792847 43126 792859
rect 43178 792847 43184 792899
rect 42160 790627 42166 790679
rect 42218 790667 42224 790679
rect 42736 790667 42742 790679
rect 42218 790639 42742 790667
rect 42218 790627 42224 790639
rect 42736 790627 42742 790639
rect 42794 790627 42800 790679
rect 42160 789887 42166 789939
rect 42218 789927 42224 789939
rect 43600 789927 43606 789939
rect 42218 789899 43606 789927
rect 42218 789887 42224 789899
rect 43600 789887 43606 789899
rect 43658 789887 43664 789939
rect 42160 789443 42166 789495
rect 42218 789483 42224 789495
rect 42448 789483 42454 789495
rect 42218 789455 42454 789483
rect 42218 789443 42224 789455
rect 42448 789443 42454 789455
rect 42506 789443 42512 789495
rect 674032 789147 674038 789199
rect 674090 789187 674096 789199
rect 675088 789187 675094 789199
rect 674090 789159 675094 789187
rect 674090 789147 674096 789159
rect 675088 789147 675094 789159
rect 675146 789147 675152 789199
rect 42160 787001 42166 787053
rect 42218 787041 42224 787053
rect 42928 787041 42934 787053
rect 42218 787013 42934 787041
rect 42218 787001 42224 787013
rect 42928 787001 42934 787013
rect 42986 787001 42992 787053
rect 42160 786409 42166 786461
rect 42218 786449 42224 786461
rect 42832 786449 42838 786461
rect 42218 786421 42838 786449
rect 42218 786409 42224 786421
rect 42832 786409 42838 786421
rect 42890 786409 42896 786461
rect 47536 786261 47542 786313
rect 47594 786301 47600 786313
rect 59536 786301 59542 786313
rect 47594 786273 59542 786301
rect 47594 786261 47600 786273
rect 59536 786261 59542 786273
rect 59594 786261 59600 786313
rect 654064 786261 654070 786313
rect 654122 786301 654128 786313
rect 666832 786301 666838 786313
rect 654122 786273 666838 786301
rect 654122 786261 654128 786273
rect 666832 786261 666838 786273
rect 666890 786261 666896 786313
rect 42064 785743 42070 785795
rect 42122 785783 42128 785795
rect 42736 785783 42742 785795
rect 42122 785755 42742 785783
rect 42122 785743 42128 785755
rect 42736 785743 42742 785755
rect 42794 785743 42800 785795
rect 672304 784263 672310 784315
rect 672362 784303 672368 784315
rect 675472 784303 675478 784315
rect 672362 784275 675478 784303
rect 672362 784263 672368 784275
rect 675472 784263 675478 784275
rect 675530 784263 675536 784315
rect 671920 783449 671926 783501
rect 671978 783489 671984 783501
rect 675376 783489 675382 783501
rect 671978 783461 675382 783489
rect 671978 783449 671984 783461
rect 675376 783449 675382 783461
rect 675434 783449 675440 783501
rect 672784 783079 672790 783131
rect 672842 783119 672848 783131
rect 675088 783119 675094 783131
rect 672842 783091 675094 783119
rect 672842 783079 672848 783091
rect 675088 783079 675094 783091
rect 675146 783119 675152 783131
rect 675472 783119 675478 783131
rect 675146 783091 675478 783119
rect 675146 783079 675152 783091
rect 675472 783079 675478 783091
rect 675530 783079 675536 783131
rect 672592 782931 672598 782983
rect 672650 782971 672656 782983
rect 675376 782971 675382 782983
rect 672650 782943 675382 782971
rect 672650 782931 672656 782943
rect 675376 782931 675382 782943
rect 675434 782931 675440 782983
rect 672400 782487 672406 782539
rect 672458 782527 672464 782539
rect 674224 782527 674230 782539
rect 672458 782499 674230 782527
rect 672458 782487 672464 782499
rect 674224 782487 674230 782499
rect 674282 782527 674288 782539
rect 675472 782527 675478 782539
rect 674282 782499 675478 782527
rect 674282 782487 674288 782499
rect 675472 782487 675478 782499
rect 675530 782487 675536 782539
rect 663856 780489 663862 780541
rect 663914 780529 663920 780541
rect 675088 780529 675094 780541
rect 663914 780501 675094 780529
rect 663914 780489 663920 780501
rect 675088 780489 675094 780501
rect 675146 780489 675152 780541
rect 42736 780415 42742 780467
rect 42794 780455 42800 780467
rect 47728 780455 47734 780467
rect 42794 780427 47734 780455
rect 42794 780415 42800 780427
rect 47728 780415 47734 780427
rect 47786 780415 47792 780467
rect 672880 779897 672886 779949
rect 672938 779937 672944 779949
rect 675376 779937 675382 779949
rect 672938 779909 675382 779937
rect 672938 779897 672944 779909
rect 675376 779897 675382 779909
rect 675434 779897 675440 779949
rect 42736 779675 42742 779727
rect 42794 779715 42800 779727
rect 50416 779715 50422 779727
rect 42794 779687 50422 779715
rect 42794 779675 42800 779687
rect 50416 779675 50422 779687
rect 50474 779675 50480 779727
rect 42736 778861 42742 778913
rect 42794 778901 42800 778913
rect 53296 778901 53302 778913
rect 42794 778873 53302 778901
rect 42794 778861 42800 778873
rect 53296 778861 53302 778873
rect 53354 778861 53360 778913
rect 672976 778565 672982 778617
rect 673034 778605 673040 778617
rect 675376 778605 675382 778617
rect 673034 778577 675382 778605
rect 673034 778565 673040 778577
rect 675376 778565 675382 778577
rect 675434 778565 675440 778617
rect 675088 777011 675094 777063
rect 675146 777051 675152 777063
rect 675376 777051 675382 777063
rect 675146 777023 675382 777051
rect 675146 777011 675152 777023
rect 675376 777011 675382 777023
rect 675434 777011 675440 777063
rect 654064 774717 654070 774769
rect 654122 774757 654128 774769
rect 666928 774757 666934 774769
rect 654122 774729 666934 774757
rect 654122 774717 654128 774729
rect 666928 774717 666934 774729
rect 666986 774717 666992 774769
rect 53488 771831 53494 771883
rect 53546 771871 53552 771883
rect 59536 771871 59542 771883
rect 53546 771843 59542 771871
rect 53546 771831 53552 771843
rect 59536 771831 59542 771843
rect 59594 771831 59600 771883
rect 660976 767465 660982 767517
rect 661034 767505 661040 767517
rect 674416 767505 674422 767517
rect 661034 767477 674422 767505
rect 661034 767465 661040 767477
rect 674416 767465 674422 767477
rect 674474 767465 674480 767517
rect 666736 766873 666742 766925
rect 666794 766913 666800 766925
rect 674608 766913 674614 766925
rect 666794 766885 674614 766913
rect 666794 766873 666800 766885
rect 674608 766873 674614 766885
rect 674666 766873 674672 766925
rect 42928 765985 42934 766037
rect 42986 766025 42992 766037
rect 43792 766025 43798 766037
rect 42986 765997 43798 766025
rect 42986 765985 42992 765997
rect 43792 765985 43798 765997
rect 43850 765985 43856 766037
rect 663952 765837 663958 765889
rect 664010 765877 664016 765889
rect 674416 765877 674422 765889
rect 664010 765849 674422 765877
rect 664010 765837 664016 765849
rect 674416 765837 674422 765849
rect 674474 765837 674480 765889
rect 672112 763469 672118 763521
rect 672170 763509 672176 763521
rect 674416 763509 674422 763521
rect 672170 763481 674422 763509
rect 672170 763469 672176 763481
rect 674416 763469 674422 763481
rect 674474 763469 674480 763521
rect 653968 763247 653974 763299
rect 654026 763287 654032 763299
rect 661168 763287 661174 763299
rect 654026 763259 661174 763287
rect 654026 763247 654032 763259
rect 661168 763247 661174 763259
rect 661226 763247 661232 763299
rect 672688 763247 672694 763299
rect 672746 763287 672752 763299
rect 673840 763287 673846 763299
rect 672746 763259 673846 763287
rect 672746 763247 672752 763259
rect 673840 763247 673846 763259
rect 673898 763247 673904 763299
rect 42160 761915 42166 761967
rect 42218 761955 42224 761967
rect 53296 761955 53302 761967
rect 42218 761927 53302 761955
rect 42218 761915 42224 761927
rect 53296 761915 53302 761927
rect 53354 761915 53360 761967
rect 672208 760361 672214 760413
rect 672266 760401 672272 760413
rect 673840 760401 673846 760413
rect 672266 760373 673846 760401
rect 672266 760361 672272 760373
rect 673840 760361 673846 760373
rect 673898 760361 673904 760413
rect 38992 760287 38998 760339
rect 39050 760327 39056 760339
rect 43024 760327 43030 760339
rect 39050 760299 43030 760327
rect 39050 760287 39056 760299
rect 43024 760287 43030 760299
rect 43082 760287 43088 760339
rect 43216 757475 43222 757527
rect 43274 757515 43280 757527
rect 45040 757515 45046 757527
rect 43274 757487 45046 757515
rect 43274 757475 43280 757487
rect 45040 757475 45046 757487
rect 45098 757475 45104 757527
rect 53680 757475 53686 757527
rect 53738 757515 53744 757527
rect 59536 757515 59542 757527
rect 53738 757487 59542 757515
rect 53738 757475 53744 757487
rect 59536 757475 59542 757487
rect 59594 757475 59600 757527
rect 41488 757401 41494 757453
rect 41546 757441 41552 757453
rect 43696 757441 43702 757453
rect 41546 757413 43702 757441
rect 41546 757401 41552 757413
rect 43696 757401 43702 757413
rect 43754 757401 43760 757453
rect 41392 757327 41398 757379
rect 41450 757367 41456 757379
rect 43600 757367 43606 757379
rect 41450 757339 43606 757367
rect 41450 757327 41456 757339
rect 43600 757327 43606 757339
rect 43658 757327 43664 757379
rect 41680 757253 41686 757305
rect 41738 757293 41744 757305
rect 43504 757293 43510 757305
rect 41738 757265 43510 757293
rect 41738 757253 41744 757265
rect 43504 757253 43510 757265
rect 43562 757253 43568 757305
rect 41872 756957 41878 757009
rect 41930 756957 41936 757009
rect 41890 756787 41918 756957
rect 41872 756735 41878 756787
rect 41930 756735 41936 756787
rect 42064 754885 42070 754937
rect 42122 754925 42128 754937
rect 43024 754925 43030 754937
rect 42122 754897 43030 754925
rect 42122 754885 42128 754897
rect 43024 754885 43030 754897
rect 43082 754885 43088 754937
rect 42160 754071 42166 754123
rect 42218 754111 42224 754123
rect 43216 754111 43222 754123
rect 42218 754083 43222 754111
rect 42218 754071 42224 754083
rect 43216 754071 43222 754083
rect 43274 754071 43280 754123
rect 43696 751851 43702 751903
rect 43754 751851 43760 751903
rect 43120 751777 43126 751829
rect 43178 751817 43184 751829
rect 43408 751817 43414 751829
rect 43178 751789 43414 751817
rect 43178 751777 43184 751789
rect 43408 751777 43414 751789
rect 43466 751777 43472 751829
rect 43024 751703 43030 751755
rect 43082 751743 43088 751755
rect 43714 751743 43742 751851
rect 43082 751715 43742 751743
rect 43082 751703 43088 751715
rect 42928 751629 42934 751681
rect 42986 751669 42992 751681
rect 43216 751669 43222 751681
rect 42986 751641 43222 751669
rect 42986 751629 42992 751641
rect 43216 751629 43222 751641
rect 43274 751629 43280 751681
rect 42160 750371 42166 750423
rect 42218 750411 42224 750423
rect 43120 750411 43126 750423
rect 42218 750383 43126 750411
rect 42218 750371 42224 750383
rect 43120 750371 43126 750383
rect 43178 750371 43184 750423
rect 43120 750223 43126 750275
rect 43178 750263 43184 750275
rect 43792 750263 43798 750275
rect 43178 750235 43798 750263
rect 43178 750223 43184 750235
rect 43792 750223 43798 750235
rect 43850 750223 43856 750275
rect 42064 749779 42070 749831
rect 42122 749819 42128 749831
rect 43024 749819 43030 749831
rect 42122 749791 43030 749819
rect 42122 749779 42128 749791
rect 43024 749779 43030 749791
rect 43082 749779 43088 749831
rect 42448 749261 42454 749313
rect 42506 749301 42512 749313
rect 43600 749301 43606 749313
rect 42506 749273 43606 749301
rect 42506 749261 42512 749273
rect 43600 749261 43606 749273
rect 43658 749261 43664 749313
rect 649648 748817 649654 748869
rect 649706 748857 649712 748869
rect 679792 748857 679798 748869
rect 649706 748829 679798 748857
rect 649706 748817 649712 748829
rect 679792 748817 679798 748829
rect 679850 748817 679856 748869
rect 672784 748743 672790 748795
rect 672842 748783 672848 748795
rect 673840 748783 673846 748795
rect 672842 748755 673846 748783
rect 672842 748743 672848 748755
rect 673840 748743 673846 748755
rect 673898 748743 673904 748795
rect 42160 746893 42166 746945
rect 42218 746933 42224 746945
rect 42928 746933 42934 746945
rect 42218 746905 42934 746933
rect 42218 746893 42224 746905
rect 42928 746893 42934 746905
rect 42986 746893 42992 746945
rect 42064 746079 42070 746131
rect 42122 746119 42128 746131
rect 42448 746119 42454 746131
rect 42122 746091 42454 746119
rect 42122 746079 42128 746091
rect 42448 746079 42454 746091
rect 42506 746079 42512 746131
rect 42160 745487 42166 745539
rect 42218 745527 42224 745539
rect 42448 745527 42454 745539
rect 42218 745499 42454 745527
rect 42218 745487 42224 745499
rect 42448 745487 42454 745499
rect 42506 745487 42512 745539
rect 42160 743785 42166 743837
rect 42218 743825 42224 743837
rect 43120 743825 43126 743837
rect 42218 743797 43126 743825
rect 42218 743785 42224 743797
rect 43120 743785 43126 743797
rect 43178 743785 43184 743837
rect 42064 743045 42070 743097
rect 42122 743085 42128 743097
rect 43024 743085 43030 743097
rect 42122 743057 43030 743085
rect 42122 743045 42128 743057
rect 43024 743045 43030 743057
rect 43082 743045 43088 743097
rect 53584 743045 53590 743097
rect 53642 743085 53648 743097
rect 59536 743085 59542 743097
rect 53642 743057 59542 743085
rect 53642 743045 53648 743057
rect 59536 743045 59542 743057
rect 59594 743045 59600 743097
rect 672400 742971 672406 743023
rect 672458 743011 672464 743023
rect 675088 743011 675094 743023
rect 672458 742983 675094 743011
rect 672458 742971 672464 742983
rect 675088 742971 675094 742983
rect 675146 742971 675152 743023
rect 42160 742601 42166 742653
rect 42218 742641 42224 742653
rect 42928 742641 42934 742653
rect 42218 742613 42934 742641
rect 42218 742601 42224 742613
rect 42928 742601 42934 742613
rect 42986 742601 42992 742653
rect 653968 740159 653974 740211
rect 654026 740199 654032 740211
rect 672400 740199 672406 740211
rect 654026 740171 672406 740199
rect 654026 740159 654032 740171
rect 672400 740159 672406 740171
rect 672458 740159 672464 740211
rect 674704 738013 674710 738065
rect 674762 738053 674768 738065
rect 675376 738053 675382 738065
rect 674762 738025 675382 738053
rect 674762 738013 674768 738025
rect 675376 738013 675382 738025
rect 675434 738013 675440 738065
rect 673840 737421 673846 737473
rect 673898 737461 673904 737473
rect 675472 737461 675478 737473
rect 673898 737433 675478 737461
rect 673898 737421 673904 737433
rect 675472 737421 675478 737433
rect 675530 737421 675536 737473
rect 660976 737273 660982 737325
rect 661034 737313 661040 737325
rect 674512 737313 674518 737325
rect 661034 737285 674518 737313
rect 661034 737273 661040 737285
rect 674512 737273 674518 737285
rect 674570 737273 674576 737325
rect 42832 737199 42838 737251
rect 42890 737239 42896 737251
rect 53488 737239 53494 737251
rect 42890 737211 53494 737239
rect 42890 737199 42896 737211
rect 53488 737199 53494 737211
rect 53546 737199 53552 737251
rect 42160 736681 42166 736733
rect 42218 736721 42224 736733
rect 53680 736721 53686 736733
rect 42218 736693 53686 736721
rect 42218 736681 42224 736693
rect 53680 736681 53686 736693
rect 53738 736681 53744 736733
rect 674608 736607 674614 736659
rect 674666 736647 674672 736659
rect 675088 736647 675094 736659
rect 674666 736619 675094 736647
rect 674666 736607 674672 736619
rect 675088 736607 675094 736619
rect 675146 736647 675152 736659
rect 675376 736647 675382 736659
rect 675146 736619 675382 736647
rect 675146 736607 675152 736619
rect 675376 736607 675382 736619
rect 675434 736607 675440 736659
rect 42832 735645 42838 735697
rect 42890 735685 42896 735697
rect 47536 735685 47542 735697
rect 42890 735657 47542 735685
rect 42890 735645 42896 735657
rect 47536 735645 47542 735657
rect 47594 735645 47600 735697
rect 675088 735423 675094 735475
rect 675146 735463 675152 735475
rect 675472 735463 675478 735475
rect 675146 735435 675478 735463
rect 675146 735423 675152 735435
rect 675472 735423 675478 735435
rect 675530 735423 675536 735475
rect 673360 734757 673366 734809
rect 673418 734797 673424 734809
rect 675376 734797 675382 734809
rect 673418 734769 675382 734797
rect 673418 734757 673424 734769
rect 675376 734757 675382 734769
rect 675434 734757 675440 734809
rect 672016 734387 672022 734439
rect 672074 734427 672080 734439
rect 675376 734427 675382 734439
rect 672074 734399 675382 734427
rect 672074 734387 672080 734399
rect 675376 734387 675382 734399
rect 675434 734387 675440 734439
rect 673168 733573 673174 733625
rect 673226 733613 673232 733625
rect 675472 733613 675478 733625
rect 673226 733585 675478 733613
rect 673226 733573 673232 733585
rect 675472 733573 675478 733585
rect 675530 733573 675536 733625
rect 672784 732315 672790 732367
rect 672842 732355 672848 732367
rect 675472 732355 675478 732367
rect 672842 732327 675478 732355
rect 672842 732315 672848 732327
rect 675472 732315 675478 732327
rect 675530 732315 675536 732367
rect 674512 732019 674518 732071
rect 674570 732059 674576 732071
rect 675376 732059 675382 732071
rect 674570 732031 675382 732059
rect 674570 732019 674576 732031
rect 675376 732019 675382 732031
rect 675434 732019 675440 732071
rect 674512 730465 674518 730517
rect 674570 730505 674576 730517
rect 675472 730505 675478 730517
rect 674570 730477 675478 730505
rect 674570 730465 674576 730477
rect 675472 730465 675478 730477
rect 675530 730465 675536 730517
rect 47536 728615 47542 728667
rect 47594 728655 47600 728667
rect 59536 728655 59542 728667
rect 47594 728627 59542 728655
rect 47594 728615 47600 728627
rect 59536 728615 59542 728627
rect 59594 728615 59600 728667
rect 674224 728615 674230 728667
rect 674282 728655 674288 728667
rect 675472 728655 675478 728667
rect 674282 728627 675478 728655
rect 674282 728615 674288 728627
rect 675472 728615 675478 728627
rect 675530 728615 675536 728667
rect 675088 727875 675094 727927
rect 675146 727915 675152 727927
rect 675568 727915 675574 727927
rect 675146 727887 675574 727915
rect 675146 727875 675152 727887
rect 675568 727875 675574 727887
rect 675626 727875 675632 727927
rect 663760 722473 663766 722525
rect 663818 722513 663824 722525
rect 674416 722513 674422 722525
rect 663818 722485 674422 722513
rect 663818 722473 663824 722485
rect 674416 722473 674422 722485
rect 674474 722473 674480 722525
rect 660880 721881 660886 721933
rect 660938 721921 660944 721933
rect 674704 721921 674710 721933
rect 660938 721893 674710 721921
rect 660938 721881 660944 721893
rect 674704 721881 674710 721893
rect 674762 721881 674768 721933
rect 661072 720845 661078 720897
rect 661130 720885 661136 720897
rect 674416 720885 674422 720897
rect 661130 720857 674422 720885
rect 661130 720845 661136 720857
rect 674416 720845 674422 720857
rect 674474 720845 674480 720897
rect 672688 720253 672694 720305
rect 672746 720293 672752 720305
rect 674704 720293 674710 720305
rect 672746 720265 674710 720293
rect 672746 720253 672752 720265
rect 674704 720253 674710 720265
rect 674762 720253 674768 720305
rect 672688 718995 672694 719047
rect 672746 719035 672752 719047
rect 674704 719035 674710 719047
rect 672746 719007 674710 719035
rect 672746 718995 672752 719007
rect 674704 718995 674710 719007
rect 674762 718995 674768 719047
rect 42448 718699 42454 718751
rect 42506 718739 42512 718751
rect 53488 718739 53494 718751
rect 42506 718711 53494 718739
rect 42506 718699 42512 718711
rect 53488 718699 53494 718711
rect 53546 718699 53552 718751
rect 654256 717145 654262 717197
rect 654314 717185 654320 717197
rect 663952 717185 663958 717197
rect 654314 717157 663958 717185
rect 654314 717145 654320 717157
rect 663952 717145 663958 717157
rect 664010 717145 664016 717197
rect 40240 717071 40246 717123
rect 40298 717111 40304 717123
rect 42448 717111 42454 717123
rect 40298 717083 42454 717111
rect 40298 717071 40304 717083
rect 42448 717071 42454 717083
rect 42506 717071 42512 717123
rect 672208 716997 672214 717049
rect 672266 717037 672272 717049
rect 673936 717037 673942 717049
rect 672266 717009 673942 717037
rect 672266 716997 672272 717009
rect 673936 716997 673942 717009
rect 673994 716997 674000 717049
rect 43504 714259 43510 714311
rect 43562 714299 43568 714311
rect 44944 714299 44950 714311
rect 43562 714271 44950 714299
rect 43562 714259 43568 714271
rect 44944 714259 44950 714271
rect 45002 714259 45008 714311
rect 50416 714259 50422 714311
rect 50474 714299 50480 714311
rect 59536 714299 59542 714311
rect 50474 714271 59542 714299
rect 50474 714259 50480 714271
rect 59536 714259 59542 714271
rect 59594 714259 59600 714311
rect 41584 714037 41590 714089
rect 41642 714077 41648 714089
rect 43696 714077 43702 714089
rect 41642 714049 43702 714077
rect 41642 714037 41648 714049
rect 43696 714037 43702 714049
rect 43754 714037 43760 714089
rect 41968 713889 41974 713941
rect 42026 713929 42032 713941
rect 43408 713929 43414 713941
rect 42026 713901 43414 713929
rect 42026 713889 42032 713901
rect 43408 713889 43414 713901
rect 43466 713889 43472 713941
rect 41872 713815 41878 713867
rect 41930 713815 41936 713867
rect 42064 713815 42070 713867
rect 42122 713855 42128 713867
rect 43312 713855 43318 713867
rect 42122 713827 43318 713855
rect 42122 713815 42128 713827
rect 43312 713815 43318 713827
rect 43370 713815 43376 713867
rect 41890 713571 41918 713815
rect 41872 713519 41878 713571
rect 41930 713519 41936 713571
rect 42448 713223 42454 713275
rect 42506 713263 42512 713275
rect 42506 713235 42590 713263
rect 42506 713223 42512 713235
rect 41872 711669 41878 711721
rect 41930 711709 41936 711721
rect 42562 711709 42590 713235
rect 41930 711681 42590 711709
rect 41930 711669 41936 711681
rect 672304 711521 672310 711573
rect 672362 711561 672368 711573
rect 674704 711561 674710 711573
rect 672362 711533 674710 711561
rect 672362 711521 672368 711533
rect 674704 711521 674710 711533
rect 674762 711521 674768 711573
rect 43120 711447 43126 711499
rect 43178 711487 43184 711499
rect 43600 711487 43606 711499
rect 43178 711459 43606 711487
rect 43178 711447 43184 711459
rect 43600 711447 43606 711459
rect 43658 711447 43664 711499
rect 43408 711373 43414 711425
rect 43466 711413 43472 711425
rect 43696 711413 43702 711425
rect 43466 711385 43702 711413
rect 43466 711373 43472 711385
rect 43696 711373 43702 711385
rect 43754 711373 43760 711425
rect 42160 710855 42166 710907
rect 42218 710895 42224 710907
rect 43504 710895 43510 710907
rect 42218 710867 43510 710895
rect 42218 710855 42224 710867
rect 43504 710855 43510 710867
rect 43562 710855 43568 710907
rect 671920 710485 671926 710537
rect 671978 710525 671984 710537
rect 674416 710525 674422 710537
rect 671978 710497 674422 710525
rect 671978 710485 671984 710497
rect 674416 710485 674422 710497
rect 674474 710485 674480 710537
rect 42160 709893 42166 709945
rect 42218 709933 42224 709945
rect 43120 709933 43126 709945
rect 42218 709905 43126 709933
rect 42218 709893 42224 709905
rect 43120 709893 43126 709905
rect 43178 709893 43184 709945
rect 672592 708413 672598 708465
rect 672650 708453 672656 708465
rect 674704 708453 674710 708465
rect 672650 708425 674710 708453
rect 672650 708413 672656 708425
rect 674704 708413 674710 708425
rect 674762 708413 674768 708465
rect 42160 707377 42166 707429
rect 42218 707417 42224 707429
rect 43312 707417 43318 707429
rect 42218 707389 43318 707417
rect 42218 707377 42224 707389
rect 43312 707377 43318 707389
rect 43370 707377 43376 707429
rect 672880 707377 672886 707429
rect 672938 707417 672944 707429
rect 674416 707417 674422 707429
rect 672938 707389 674422 707417
rect 672938 707377 672944 707389
rect 674416 707377 674422 707389
rect 674474 707377 674480 707429
rect 672976 706785 672982 706837
rect 673034 706825 673040 706837
rect 674704 706825 674710 706837
rect 673034 706797 674710 706825
rect 673034 706785 673040 706797
rect 674704 706785 674710 706797
rect 674762 706785 674768 706837
rect 42160 704269 42166 704321
rect 42218 704309 42224 704321
rect 43024 704309 43030 704321
rect 42218 704281 43030 704309
rect 42218 704269 42224 704281
rect 43024 704269 43030 704281
rect 43082 704269 43088 704321
rect 43024 704121 43030 704173
rect 43082 704161 43088 704173
rect 43408 704161 43414 704173
rect 43082 704133 43414 704161
rect 43082 704121 43088 704133
rect 43408 704121 43414 704133
rect 43466 704121 43472 704173
rect 42064 703529 42070 703581
rect 42122 703569 42128 703581
rect 43120 703569 43126 703581
rect 42122 703541 43126 703569
rect 42122 703529 42128 703541
rect 43120 703529 43126 703541
rect 43178 703529 43184 703581
rect 43120 703381 43126 703433
rect 43178 703421 43184 703433
rect 43600 703421 43606 703433
rect 43178 703393 43606 703421
rect 43178 703381 43184 703393
rect 43600 703381 43606 703393
rect 43658 703381 43664 703433
rect 42160 702863 42166 702915
rect 42218 702903 42224 702915
rect 43024 702903 43030 702915
rect 42218 702875 43030 702903
rect 42218 702863 42224 702875
rect 43024 702863 43030 702875
rect 43082 702863 43088 702915
rect 649744 702715 649750 702767
rect 649802 702755 649808 702767
rect 679792 702755 679798 702767
rect 649802 702727 679798 702755
rect 649802 702715 649808 702727
rect 679792 702715 679798 702727
rect 679850 702715 679856 702767
rect 673840 702641 673846 702693
rect 673898 702681 673904 702693
rect 674704 702681 674710 702693
rect 673898 702653 674710 702681
rect 673898 702641 673904 702653
rect 674704 702641 674710 702653
rect 674762 702641 674768 702693
rect 42160 702419 42166 702471
rect 42218 702459 42224 702471
rect 42736 702459 42742 702471
rect 42218 702431 42742 702459
rect 42218 702419 42224 702431
rect 42736 702419 42742 702431
rect 42794 702419 42800 702471
rect 42064 700421 42070 700473
rect 42122 700461 42128 700473
rect 43120 700461 43126 700473
rect 42122 700433 43126 700461
rect 42122 700421 42128 700433
rect 43120 700421 43126 700433
rect 43178 700421 43184 700473
rect 42160 700051 42166 700103
rect 42218 700091 42224 700103
rect 42448 700091 42454 700103
rect 42218 700063 42454 700091
rect 42218 700051 42224 700063
rect 42448 700051 42454 700063
rect 42506 700051 42512 700103
rect 42448 699829 42454 699881
rect 42506 699869 42512 699881
rect 59536 699869 59542 699881
rect 42506 699841 59542 699869
rect 42506 699829 42512 699841
rect 59536 699829 59542 699841
rect 59594 699829 59600 699881
rect 42160 699163 42166 699215
rect 42218 699203 42224 699215
rect 43024 699203 43030 699215
rect 42218 699175 43030 699203
rect 42218 699163 42224 699175
rect 43024 699163 43030 699175
rect 43082 699163 43088 699215
rect 674320 698941 674326 698993
rect 674378 698981 674384 698993
rect 675568 698981 675574 698993
rect 674378 698953 675574 698981
rect 674378 698941 674384 698953
rect 675568 698941 675574 698953
rect 675626 698941 675632 698993
rect 654448 694057 654454 694109
rect 654506 694097 654512 694109
rect 669808 694097 669814 694109
rect 654506 694069 669814 694097
rect 654506 694057 654512 694069
rect 669808 694057 669814 694069
rect 669866 694057 669872 694109
rect 42832 693983 42838 694035
rect 42890 694023 42896 694035
rect 50416 694023 50422 694035
rect 42890 693995 50422 694023
rect 42890 693983 42896 693995
rect 50416 693983 50422 693995
rect 50474 693983 50480 694035
rect 672304 692873 672310 692925
rect 672362 692913 672368 692925
rect 675376 692913 675382 692925
rect 672362 692885 675382 692913
rect 672362 692873 672368 692885
rect 675376 692873 675382 692885
rect 675434 692873 675440 692925
rect 42448 692725 42454 692777
rect 42506 692765 42512 692777
rect 47536 692765 47542 692777
rect 42506 692737 47542 692765
rect 42506 692725 42512 692737
rect 47536 692725 47542 692737
rect 47594 692725 47600 692777
rect 672976 692429 672982 692481
rect 673034 692469 673040 692481
rect 674704 692469 674710 692481
rect 673034 692441 674710 692469
rect 673034 692429 673040 692441
rect 674704 692429 674710 692441
rect 674762 692469 674768 692481
rect 675472 692469 675478 692481
rect 674762 692441 675478 692469
rect 674762 692429 674768 692441
rect 675472 692429 675478 692441
rect 675530 692429 675536 692481
rect 674608 692281 674614 692333
rect 674666 692321 674672 692333
rect 675376 692321 675382 692333
rect 674666 692293 675382 692321
rect 674666 692281 674672 692293
rect 675376 692281 675382 692293
rect 675434 692281 675440 692333
rect 674800 690653 674806 690705
rect 674858 690693 674864 690705
rect 675472 690693 675478 690705
rect 674858 690665 675478 690693
rect 674858 690653 674864 690665
rect 675472 690653 675478 690665
rect 675530 690653 675536 690705
rect 674896 689765 674902 689817
rect 674954 689805 674960 689817
rect 675376 689805 675382 689817
rect 674954 689777 675382 689805
rect 674954 689765 674960 689777
rect 675376 689765 675382 689777
rect 675434 689765 675440 689817
rect 673072 688581 673078 688633
rect 673130 688621 673136 688633
rect 675472 688621 675478 688633
rect 673130 688593 675478 688621
rect 673130 688581 673136 688593
rect 675472 688581 675478 688593
rect 675530 688581 675536 688633
rect 674896 687323 674902 687375
rect 674954 687363 674960 687375
rect 675472 687363 675478 687375
rect 674954 687335 675478 687363
rect 674954 687323 674960 687335
rect 675472 687323 675478 687335
rect 675530 687323 675536 687375
rect 669616 686213 669622 686265
rect 669674 686253 669680 686265
rect 675376 686253 675382 686265
rect 669674 686225 675382 686253
rect 669674 686213 669680 686225
rect 675376 686213 675382 686225
rect 675434 686213 675440 686265
rect 47536 685473 47542 685525
rect 47594 685513 47600 685525
rect 59536 685513 59542 685525
rect 47594 685485 59542 685513
rect 47594 685473 47600 685485
rect 59536 685473 59542 685485
rect 59594 685473 59600 685525
rect 674416 685473 674422 685525
rect 674474 685513 674480 685525
rect 675472 685513 675478 685525
rect 674474 685485 675478 685513
rect 674474 685473 674480 685485
rect 675472 685473 675478 685485
rect 675530 685473 675536 685525
rect 674032 683623 674038 683675
rect 674090 683663 674096 683675
rect 675472 683663 675478 683675
rect 674090 683635 675478 683663
rect 674090 683623 674096 683635
rect 675472 683623 675478 683635
rect 675530 683623 675536 683675
rect 674896 681921 674902 681973
rect 674954 681961 674960 681973
rect 675472 681961 675478 681973
rect 674954 681933 675478 681961
rect 674954 681921 674960 681933
rect 675472 681921 675478 681933
rect 675530 681921 675536 681973
rect 672112 681329 672118 681381
rect 672170 681369 672176 681381
rect 673744 681369 673750 681381
rect 672170 681341 673750 681369
rect 672170 681329 672176 681341
rect 673744 681329 673750 681341
rect 673802 681329 673808 681381
rect 672496 677481 672502 677533
rect 672554 677521 672560 677533
rect 674704 677521 674710 677533
rect 672554 677493 674710 677521
rect 672554 677481 672560 677493
rect 674704 677481 674710 677493
rect 674762 677481 674768 677533
rect 672688 676741 672694 676793
rect 672746 676781 672752 676793
rect 673840 676781 673846 676793
rect 672746 676753 673846 676781
rect 672746 676741 672752 676753
rect 673840 676741 673846 676753
rect 673898 676741 673904 676793
rect 669712 676667 669718 676719
rect 669770 676707 669776 676719
rect 674704 676707 674710 676719
rect 669770 676679 674710 676707
rect 669770 676667 669776 676679
rect 674704 676667 674710 676679
rect 674762 676667 674768 676719
rect 674704 676001 674710 676053
rect 674762 676041 674768 676053
rect 674992 676041 674998 676053
rect 674762 676013 674998 676041
rect 674762 676001 674768 676013
rect 674992 676001 674998 676013
rect 675050 676001 675056 676053
rect 664048 675853 664054 675905
rect 664106 675893 664112 675905
rect 674704 675893 674710 675905
rect 664106 675865 674710 675893
rect 664106 675853 664112 675865
rect 674704 675853 674710 675865
rect 674762 675853 674768 675905
rect 42448 675779 42454 675831
rect 42506 675819 42512 675831
rect 53680 675819 53686 675831
rect 42506 675791 53686 675819
rect 42506 675779 42512 675791
rect 53680 675779 53686 675791
rect 53738 675779 53744 675831
rect 42160 674965 42166 675017
rect 42218 675005 42224 675017
rect 42448 675005 42454 675017
rect 42218 674977 42454 675005
rect 42218 674965 42224 674977
rect 42448 674965 42454 674977
rect 42506 674965 42512 675017
rect 41776 674521 41782 674573
rect 41834 674561 41840 674573
rect 41968 674561 41974 674573
rect 41834 674533 41974 674561
rect 41834 674521 41840 674533
rect 41968 674521 41974 674533
rect 42026 674521 42032 674573
rect 43600 673707 43606 673759
rect 43658 673747 43664 673759
rect 44848 673747 44854 673759
rect 43658 673719 44854 673747
rect 43658 673707 43664 673719
rect 44848 673707 44854 673719
rect 44906 673707 44912 673759
rect 40144 672227 40150 672279
rect 40202 672267 40208 672279
rect 41776 672267 41782 672279
rect 40202 672239 41782 672267
rect 40202 672227 40208 672239
rect 41776 672227 41782 672239
rect 41834 672227 41840 672279
rect 50416 671043 50422 671095
rect 50474 671083 50480 671095
rect 59536 671083 59542 671095
rect 50474 671055 59542 671083
rect 50474 671043 50480 671055
rect 59536 671043 59542 671055
rect 59594 671043 59600 671095
rect 654448 671043 654454 671095
rect 654506 671083 654512 671095
rect 661072 671083 661078 671095
rect 654506 671055 661078 671083
rect 654506 671043 654512 671055
rect 661072 671043 661078 671055
rect 661130 671043 661136 671095
rect 40912 670895 40918 670947
rect 40970 670935 40976 670947
rect 43312 670935 43318 670947
rect 40970 670907 43318 670935
rect 40970 670895 40976 670907
rect 43312 670895 43318 670907
rect 43370 670895 43376 670947
rect 41680 670821 41686 670873
rect 41738 670861 41744 670873
rect 42160 670861 42166 670873
rect 41738 670833 42166 670861
rect 41738 670821 41744 670833
rect 42160 670821 42166 670833
rect 42218 670821 42224 670873
rect 41872 670673 41878 670725
rect 41930 670713 41936 670725
rect 43024 670713 43030 670725
rect 41930 670685 43030 670713
rect 41930 670673 41936 670685
rect 43024 670673 43030 670685
rect 43082 670673 43088 670725
rect 41776 670599 41782 670651
rect 41834 670639 41840 670651
rect 43120 670639 43126 670651
rect 41834 670611 43126 670639
rect 41834 670599 41840 670611
rect 43120 670599 43126 670611
rect 43178 670599 43184 670651
rect 42448 670081 42454 670133
rect 42506 670121 42512 670133
rect 43408 670121 43414 670133
rect 42506 670093 43414 670121
rect 42506 670081 42512 670093
rect 43408 670081 43414 670093
rect 43466 670081 43472 670133
rect 43024 668937 43030 668949
rect 42754 668909 43030 668937
rect 42754 668727 42782 668909
rect 43024 668897 43030 668909
rect 43082 668897 43088 668949
rect 42736 668675 42742 668727
rect 42794 668675 42800 668727
rect 42832 668675 42838 668727
rect 42890 668715 42896 668727
rect 43312 668715 43318 668727
rect 42890 668687 43318 668715
rect 42890 668675 42896 668687
rect 43312 668675 43318 668687
rect 43370 668675 43376 668727
rect 42160 668527 42166 668579
rect 42218 668567 42224 668579
rect 43120 668567 43126 668579
rect 42218 668539 43126 668567
rect 42218 668527 42224 668539
rect 43120 668527 43126 668539
rect 43178 668527 43184 668579
rect 42160 667861 42166 667913
rect 42218 667901 42224 667913
rect 43696 667901 43702 667913
rect 42218 667873 43702 667901
rect 42218 667861 42224 667873
rect 43696 667861 43702 667873
rect 43754 667861 43760 667913
rect 42160 666677 42166 666729
rect 42218 666717 42224 666729
rect 43120 666717 43126 666729
rect 42218 666689 43126 666717
rect 42218 666677 42224 666689
rect 43120 666677 43126 666689
rect 43178 666677 43184 666729
rect 43600 665271 43606 665323
rect 43658 665311 43664 665323
rect 43888 665311 43894 665323
rect 43658 665283 43894 665311
rect 43658 665271 43664 665283
rect 43888 665271 43894 665283
rect 43946 665271 43952 665323
rect 672784 665197 672790 665249
rect 672842 665237 672848 665249
rect 673840 665237 673846 665249
rect 672842 665209 673846 665237
rect 672842 665197 672848 665209
rect 673840 665197 673846 665209
rect 673898 665197 673904 665249
rect 674032 665197 674038 665249
rect 674090 665237 674096 665249
rect 674320 665237 674326 665249
rect 674090 665209 674326 665237
rect 674090 665197 674096 665209
rect 674320 665197 674326 665209
rect 674378 665197 674384 665249
rect 42160 664827 42166 664879
rect 42218 664867 42224 664879
rect 43600 664867 43606 664879
rect 42218 664839 43606 664867
rect 42218 664827 42224 664839
rect 43600 664827 43606 664839
rect 43658 664827 43664 664879
rect 672016 664309 672022 664361
rect 672074 664349 672080 664361
rect 673840 664349 673846 664361
rect 672074 664321 673846 664349
rect 672074 664309 672080 664321
rect 673840 664309 673846 664321
rect 673898 664309 673904 664361
rect 42064 664161 42070 664213
rect 42122 664201 42128 664213
rect 43120 664201 43126 664213
rect 42122 664173 43126 664201
rect 42122 664161 42128 664173
rect 43120 664161 43126 664173
rect 43178 664161 43184 664213
rect 42160 663495 42166 663547
rect 42218 663535 42224 663547
rect 42832 663535 42838 663547
rect 42218 663507 42838 663535
rect 42218 663495 42224 663507
rect 42832 663495 42838 663507
rect 42890 663495 42896 663547
rect 674608 660905 674614 660957
rect 674666 660945 674672 660957
rect 674992 660945 674998 660957
rect 674666 660917 674998 660945
rect 674666 660905 674672 660917
rect 674992 660905 674998 660917
rect 675050 660905 675056 660957
rect 42064 660831 42070 660883
rect 42122 660871 42128 660883
rect 42736 660871 42742 660883
rect 42122 660843 42742 660871
rect 42122 660831 42128 660843
rect 42736 660831 42742 660843
rect 42794 660831 42800 660883
rect 42160 659647 42166 659699
rect 42218 659687 42224 659699
rect 42832 659687 42838 659699
rect 42218 659659 42838 659687
rect 42218 659647 42224 659659
rect 42832 659647 42838 659659
rect 42890 659647 42896 659699
rect 42064 657353 42070 657405
rect 42122 657393 42128 657405
rect 42448 657393 42454 657405
rect 42122 657365 42454 657393
rect 42122 657353 42128 657365
rect 42448 657353 42454 657365
rect 42506 657353 42512 657405
rect 674896 656761 674902 656813
rect 674954 656801 674960 656813
rect 675472 656801 675478 656813
rect 674954 656773 675478 656801
rect 674954 656761 674960 656773
rect 675472 656761 675478 656773
rect 675530 656761 675536 656813
rect 42448 656687 42454 656739
rect 42506 656727 42512 656739
rect 59536 656727 59542 656739
rect 42506 656699 59542 656727
rect 42506 656687 42512 656699
rect 59536 656687 59542 656699
rect 59594 656687 59600 656739
rect 649840 656687 649846 656739
rect 649898 656727 649904 656739
rect 679696 656727 679702 656739
rect 649898 656699 679702 656727
rect 649898 656687 649904 656699
rect 679696 656687 679702 656699
rect 679754 656687 679760 656739
rect 42160 656169 42166 656221
rect 42218 656209 42224 656221
rect 43120 656209 43126 656221
rect 42218 656181 43126 656209
rect 42218 656169 42224 656181
rect 43120 656169 43126 656181
rect 43178 656169 43184 656221
rect 672976 653727 672982 653779
rect 673034 653767 673040 653779
rect 674224 653767 674230 653779
rect 673034 653739 674230 653767
rect 673034 653727 673040 653739
rect 674224 653727 674230 653739
rect 674282 653727 674288 653779
rect 42448 649731 42454 649783
rect 42506 649771 42512 649783
rect 51856 649771 51862 649783
rect 42506 649743 51862 649771
rect 42506 649731 42512 649743
rect 51856 649731 51862 649743
rect 51914 649731 51920 649783
rect 42448 649509 42454 649561
rect 42506 649549 42512 649561
rect 50416 649549 50422 649561
rect 42506 649521 50422 649549
rect 42506 649509 42512 649521
rect 50416 649509 50422 649521
rect 50474 649509 50480 649561
rect 673360 648251 673366 648303
rect 673418 648291 673424 648303
rect 675376 648291 675382 648303
rect 673418 648263 675382 648291
rect 673418 648251 673424 648263
rect 675376 648251 675382 648263
rect 675434 648251 675440 648303
rect 654256 648029 654262 648081
rect 654314 648069 654320 648081
rect 672592 648069 672598 648081
rect 654314 648041 672598 648069
rect 654314 648029 654320 648041
rect 672592 648029 672598 648041
rect 672650 648029 672656 648081
rect 672208 647955 672214 648007
rect 672266 647995 672272 648007
rect 675376 647995 675382 648007
rect 672266 647967 675382 647995
rect 672266 647955 672272 647967
rect 675376 647955 675382 647967
rect 675434 647955 675440 648007
rect 674224 647067 674230 647119
rect 674282 647107 674288 647119
rect 675376 647107 675382 647119
rect 674282 647079 675382 647107
rect 674282 647067 674288 647079
rect 675376 647067 675382 647079
rect 675434 647067 675440 647119
rect 674800 646401 674806 646453
rect 674858 646441 674864 646453
rect 675376 646441 675382 646453
rect 674858 646413 675382 646441
rect 674858 646401 674864 646413
rect 675376 646401 675382 646413
rect 675434 646401 675440 646453
rect 672784 644551 672790 644603
rect 672842 644591 672848 644603
rect 675472 644591 675478 644603
rect 672842 644563 675478 644591
rect 672842 644551 672848 644563
rect 675472 644551 675478 644563
rect 675530 644551 675536 644603
rect 51856 644477 51862 644529
rect 51914 644517 51920 644529
rect 59248 644517 59254 644529
rect 51914 644489 59254 644517
rect 51914 644477 51920 644489
rect 59248 644477 59254 644489
rect 59306 644477 59312 644529
rect 672688 644033 672694 644085
rect 672746 644073 672752 644085
rect 675472 644073 675478 644085
rect 672746 644045 675478 644073
rect 672746 644033 672752 644045
rect 675472 644033 675478 644045
rect 675530 644033 675536 644085
rect 672880 643367 672886 643419
rect 672938 643407 672944 643419
rect 675376 643407 675382 643419
rect 672938 643379 675382 643407
rect 672938 643367 672944 643379
rect 675376 643367 675382 643379
rect 675434 643367 675440 643419
rect 672496 642257 672502 642309
rect 672554 642297 672560 642309
rect 675472 642297 675478 642309
rect 672554 642269 675478 642297
rect 672554 642257 672560 642269
rect 675472 642257 675478 642269
rect 675530 642257 675536 642309
rect 666736 641073 666742 641125
rect 666794 641113 666800 641125
rect 675472 641113 675478 641125
rect 666794 641085 675478 641113
rect 666794 641073 666800 641085
rect 675472 641073 675478 641085
rect 675530 641073 675536 641125
rect 674800 638187 674806 638239
rect 674858 638227 674864 638239
rect 675568 638227 675574 638239
rect 674858 638199 675574 638227
rect 674858 638187 674864 638199
rect 675568 638187 675574 638199
rect 675626 638187 675632 638239
rect 674704 638113 674710 638165
rect 674762 638153 674768 638165
rect 675376 638153 675382 638165
rect 674762 638125 675382 638153
rect 674762 638113 674768 638125
rect 675376 638113 675382 638125
rect 675434 638113 675440 638165
rect 666928 632489 666934 632541
rect 666986 632529 666992 632541
rect 674512 632529 674518 632541
rect 666986 632501 674518 632529
rect 666986 632489 666992 632501
rect 674512 632489 674518 632501
rect 674570 632489 674576 632541
rect 666832 631749 666838 631801
rect 666890 631789 666896 631801
rect 674512 631789 674518 631801
rect 666890 631761 674518 631789
rect 666890 631749 666896 631761
rect 674512 631749 674518 631761
rect 674570 631749 674576 631801
rect 43120 630787 43126 630839
rect 43178 630827 43184 630839
rect 43696 630827 43702 630839
rect 43178 630799 43702 630827
rect 43178 630787 43184 630799
rect 43696 630787 43702 630799
rect 43754 630787 43760 630839
rect 42448 630713 42454 630765
rect 42506 630753 42512 630765
rect 56080 630753 56086 630765
rect 42506 630725 56086 630753
rect 42506 630713 42512 630725
rect 56080 630713 56086 630725
rect 56138 630713 56144 630765
rect 661168 630639 661174 630691
rect 661226 630679 661232 630691
rect 674128 630679 674134 630691
rect 661226 630651 674134 630679
rect 661226 630639 661232 630651
rect 674128 630639 674134 630651
rect 674186 630639 674192 630691
rect 43408 627901 43414 627953
rect 43466 627941 43472 627953
rect 44752 627941 44758 627953
rect 43466 627913 44758 627941
rect 43466 627901 43472 627913
rect 44752 627901 44758 627913
rect 44810 627901 44816 627953
rect 671920 627901 671926 627953
rect 671978 627941 671984 627953
rect 673744 627941 673750 627953
rect 671978 627913 673750 627941
rect 671978 627901 671984 627913
rect 673744 627901 673750 627913
rect 673802 627901 673808 627953
rect 39856 627827 39862 627879
rect 39914 627867 39920 627879
rect 43024 627867 43030 627879
rect 39914 627839 43030 627867
rect 39914 627827 39920 627839
rect 43024 627827 43030 627839
rect 43082 627827 43088 627879
rect 43120 627827 43126 627879
rect 43178 627867 43184 627879
rect 43312 627867 43318 627879
rect 43178 627839 43318 627867
rect 43178 627827 43184 627839
rect 43312 627827 43318 627839
rect 43370 627827 43376 627879
rect 50416 627827 50422 627879
rect 50474 627867 50480 627879
rect 59536 627867 59542 627879
rect 50474 627839 59542 627867
rect 50474 627827 50480 627839
rect 59536 627827 59542 627839
rect 59594 627827 59600 627879
rect 672016 627827 672022 627879
rect 672074 627867 672080 627879
rect 673840 627867 673846 627879
rect 672074 627839 673846 627867
rect 672074 627827 672080 627839
rect 673840 627827 673846 627839
rect 673898 627827 673904 627879
rect 41488 627753 41494 627805
rect 41546 627793 41552 627805
rect 43504 627793 43510 627805
rect 41546 627765 43510 627793
rect 41546 627753 41552 627765
rect 43504 627753 43510 627765
rect 43562 627753 43568 627805
rect 673264 627753 673270 627805
rect 673322 627793 673328 627805
rect 675376 627793 675382 627805
rect 673322 627765 675382 627793
rect 673322 627753 673328 627765
rect 675376 627753 675382 627765
rect 675434 627753 675440 627805
rect 41680 627679 41686 627731
rect 41738 627719 41744 627731
rect 43120 627719 43126 627731
rect 41738 627691 43126 627719
rect 41738 627679 41744 627691
rect 43120 627679 43126 627691
rect 43178 627679 43184 627731
rect 41872 627383 41878 627435
rect 41930 627383 41936 627435
rect 41968 627383 41974 627435
rect 42026 627423 42032 627435
rect 42928 627423 42934 627435
rect 42026 627395 42934 627423
rect 42026 627383 42032 627395
rect 42928 627383 42934 627395
rect 42986 627383 42992 627435
rect 41890 627213 41918 627383
rect 41872 627161 41878 627213
rect 41930 627161 41936 627213
rect 42160 625311 42166 625363
rect 42218 625351 42224 625363
rect 43024 625351 43030 625363
rect 42218 625323 43030 625351
rect 42218 625311 42224 625323
rect 43024 625311 43030 625323
rect 43082 625311 43088 625363
rect 43024 625163 43030 625215
rect 43082 625203 43088 625215
rect 43312 625203 43318 625215
rect 43082 625175 43318 625203
rect 43082 625163 43088 625175
rect 43312 625163 43318 625175
rect 43370 625163 43376 625215
rect 42160 624645 42166 624697
rect 42218 624685 42224 624697
rect 43408 624685 43414 624697
rect 42218 624657 43414 624685
rect 42218 624645 42224 624657
rect 43408 624645 43414 624657
rect 43466 624645 43472 624697
rect 674896 623757 674902 623809
rect 674954 623797 674960 623809
rect 675376 623797 675382 623809
rect 674954 623769 675382 623797
rect 674954 623757 674960 623769
rect 675376 623757 675382 623769
rect 675434 623757 675440 623809
rect 42160 623461 42166 623513
rect 42218 623501 42224 623513
rect 42928 623501 42934 623513
rect 42218 623473 42934 623501
rect 42218 623461 42224 623473
rect 42928 623461 42934 623473
rect 42986 623461 42992 623513
rect 42928 623313 42934 623365
rect 42986 623353 42992 623365
rect 43504 623353 43510 623365
rect 42986 623325 43510 623353
rect 42986 623313 42992 623325
rect 43504 623313 43510 623325
rect 43562 623313 43568 623365
rect 42160 622203 42166 622255
rect 42218 622243 42224 622255
rect 43024 622243 43030 622255
rect 42218 622215 43030 622243
rect 42218 622203 42224 622215
rect 43024 622203 43030 622215
rect 43082 622203 43088 622255
rect 654352 622055 654358 622107
rect 654410 622095 654416 622107
rect 669712 622095 669718 622107
rect 654410 622067 669718 622095
rect 654410 622055 654416 622067
rect 669712 622055 669718 622067
rect 669770 622055 669776 622107
rect 42160 620353 42166 620405
rect 42218 620393 42224 620405
rect 43120 620393 43126 620405
rect 42218 620365 43126 620393
rect 42218 620353 42224 620365
rect 43120 620353 43126 620365
rect 43178 620353 43184 620405
rect 672304 617985 672310 618037
rect 672362 618025 672368 618037
rect 674416 618025 674422 618037
rect 672362 617997 674422 618025
rect 672362 617985 672368 617997
rect 674416 617985 674422 617997
rect 674474 617985 674480 618037
rect 42160 617319 42166 617371
rect 42218 617359 42224 617371
rect 43312 617359 43318 617371
rect 42218 617331 43318 617359
rect 42218 617319 42224 617331
rect 43312 617319 43318 617331
rect 43370 617319 43376 617371
rect 42160 615839 42166 615891
rect 42218 615879 42224 615891
rect 43120 615879 43126 615891
rect 42218 615851 43126 615879
rect 42218 615839 42224 615851
rect 43120 615839 43126 615851
rect 43178 615839 43184 615891
rect 42160 614137 42166 614189
rect 42218 614177 42224 614189
rect 43696 614177 43702 614189
rect 42218 614149 43702 614177
rect 42218 614137 42224 614149
rect 43696 614137 43702 614149
rect 43754 614137 43760 614189
rect 42736 613471 42742 613523
rect 42794 613511 42800 613523
rect 59536 613511 59542 613523
rect 42794 613483 59542 613511
rect 42794 613471 42800 613483
rect 59536 613471 59542 613483
rect 59594 613471 59600 613523
rect 649936 613471 649942 613523
rect 649994 613511 650000 613523
rect 679696 613511 679702 613523
rect 649994 613483 679702 613511
rect 649994 613471 650000 613483
rect 679696 613471 679702 613483
rect 679754 613471 679760 613523
rect 654352 613397 654358 613449
rect 654410 613437 654416 613449
rect 669520 613437 669526 613449
rect 654410 613409 669526 613437
rect 654410 613397 654416 613409
rect 669520 613397 669526 613409
rect 669578 613397 669584 613449
rect 674992 613397 674998 613449
rect 675050 613437 675056 613449
rect 675568 613437 675574 613449
rect 675050 613409 675574 613437
rect 675050 613397 675056 613409
rect 675568 613397 675574 613409
rect 675626 613397 675632 613449
rect 674224 613323 674230 613375
rect 674282 613363 674288 613375
rect 675088 613363 675094 613375
rect 674282 613335 675094 613363
rect 674282 613323 674288 613335
rect 675088 613323 675094 613335
rect 675146 613323 675152 613375
rect 42160 607847 42166 607899
rect 42218 607887 42224 607899
rect 42736 607887 42742 607899
rect 42218 607859 42742 607887
rect 42218 607847 42224 607859
rect 42736 607847 42742 607859
rect 42794 607847 42800 607899
rect 42736 607699 42742 607751
rect 42794 607739 42800 607751
rect 51856 607739 51862 607751
rect 42794 607711 51862 607739
rect 42794 607699 42800 607711
rect 51856 607699 51862 607711
rect 51914 607699 51920 607751
rect 42736 606811 42742 606863
rect 42794 606851 42800 606863
rect 53872 606851 53878 606863
rect 42794 606823 53878 606851
rect 42794 606811 42800 606823
rect 53872 606811 53878 606823
rect 53930 606811 53936 606863
rect 672976 604073 672982 604125
rect 673034 604113 673040 604125
rect 675472 604113 675478 604125
rect 673034 604085 675478 604113
rect 673034 604073 673040 604085
rect 675472 604073 675478 604085
rect 675530 604073 675536 604125
rect 673072 603259 673078 603311
rect 673130 603299 673136 603311
rect 675376 603299 675382 603311
rect 673130 603271 675382 603299
rect 673130 603259 673136 603271
rect 675376 603259 675382 603271
rect 675434 603259 675440 603311
rect 673744 603037 673750 603089
rect 673802 603077 673808 603089
rect 675088 603077 675094 603089
rect 673802 603049 675094 603077
rect 673802 603037 673808 603049
rect 675088 603037 675094 603049
rect 675146 603077 675152 603089
rect 675376 603077 675382 603089
rect 675146 603049 675382 603077
rect 675146 603037 675152 603049
rect 675376 603037 675382 603049
rect 675434 603037 675440 603089
rect 671632 602889 671638 602941
rect 671690 602929 671696 602941
rect 675472 602929 675478 602941
rect 671690 602901 675478 602929
rect 671690 602889 671696 602901
rect 675472 602889 675478 602901
rect 675530 602889 675536 602941
rect 672304 602445 672310 602497
rect 672362 602485 672368 602497
rect 674992 602485 674998 602497
rect 672362 602457 674998 602485
rect 672362 602445 672368 602457
rect 674992 602445 674998 602457
rect 675050 602485 675056 602497
rect 675376 602485 675382 602497
rect 675050 602457 675382 602485
rect 675050 602445 675056 602457
rect 675376 602445 675382 602457
rect 675434 602445 675440 602497
rect 663760 601927 663766 601979
rect 663818 601967 663824 601979
rect 674416 601967 674422 601979
rect 663818 601939 674422 601967
rect 663818 601927 663824 601939
rect 674416 601927 674422 601939
rect 674474 601927 674480 601979
rect 51856 601853 51862 601905
rect 51914 601893 51920 601905
rect 59536 601893 59542 601905
rect 51914 601865 59542 601893
rect 51914 601853 51920 601865
rect 59536 601853 59542 601865
rect 59594 601853 59600 601905
rect 673552 599559 673558 599611
rect 673610 599599 673616 599611
rect 675376 599599 675382 599611
rect 673610 599571 675382 599599
rect 673610 599559 673616 599571
rect 675376 599559 675382 599571
rect 675434 599559 675440 599611
rect 671824 599263 671830 599315
rect 671882 599303 671888 599315
rect 675376 599303 675382 599315
rect 671882 599275 675382 599303
rect 671882 599263 671888 599275
rect 675376 599263 675382 599275
rect 675434 599263 675440 599315
rect 654448 599041 654454 599093
rect 654506 599081 654512 599093
rect 666832 599081 666838 599093
rect 654506 599053 666838 599081
rect 654506 599041 654512 599053
rect 666832 599041 666838 599053
rect 666890 599041 666896 599093
rect 673168 598375 673174 598427
rect 673226 598415 673232 598427
rect 675472 598415 675478 598427
rect 673226 598387 675478 598415
rect 673226 598375 673232 598387
rect 675472 598375 675478 598387
rect 675530 598375 675536 598427
rect 672112 597117 672118 597169
rect 672170 597157 672176 597169
rect 675472 597157 675478 597169
rect 672170 597129 675478 597157
rect 672170 597117 672176 597129
rect 675472 597117 675478 597129
rect 675530 597117 675536 597169
rect 674416 596821 674422 596873
rect 674474 596861 674480 596873
rect 675376 596861 675382 596873
rect 674474 596833 675382 596861
rect 674474 596821 674480 596833
rect 675376 596821 675382 596833
rect 675434 596821 675440 596873
rect 674896 595267 674902 595319
rect 674954 595307 674960 595319
rect 675472 595307 675478 595319
rect 674954 595279 675478 595307
rect 674954 595267 674960 595279
rect 675472 595267 675478 595279
rect 675530 595267 675536 595319
rect 53872 587423 53878 587475
rect 53930 587463 53936 587475
rect 58192 587463 58198 587475
rect 53930 587435 58198 587463
rect 53930 587423 53936 587435
rect 58192 587423 58198 587435
rect 58250 587423 58256 587475
rect 672400 587423 672406 587475
rect 672458 587463 672464 587475
rect 673840 587463 673846 587475
rect 672458 587435 673846 587463
rect 672458 587423 672464 587435
rect 673840 587423 673846 587435
rect 673898 587423 673904 587475
rect 672016 586165 672022 586217
rect 672074 586205 672080 586217
rect 673840 586205 673846 586217
rect 672074 586177 673846 586205
rect 672074 586165 672080 586177
rect 673840 586165 673846 586177
rect 673898 586165 673904 586217
rect 41872 586091 41878 586143
rect 41930 586131 41936 586143
rect 42736 586131 42742 586143
rect 41930 586103 42742 586131
rect 41930 586091 41936 586103
rect 42736 586091 42742 586103
rect 42794 586091 42800 586143
rect 40048 585943 40054 585995
rect 40106 585983 40112 585995
rect 41872 585983 41878 585995
rect 40106 585955 41878 585983
rect 40106 585943 40112 585955
rect 41872 585943 41878 585955
rect 41930 585943 41936 585995
rect 663952 585425 663958 585477
rect 664010 585465 664016 585477
rect 674416 585465 674422 585477
rect 664010 585437 674422 585465
rect 664010 585425 664016 585437
rect 674416 585425 674422 585437
rect 674474 585425 674480 585477
rect 655216 584759 655222 584811
rect 655274 584799 655280 584811
rect 674608 584799 674614 584811
rect 655274 584771 674614 584799
rect 655274 584759 655280 584771
rect 674608 584759 674614 584771
rect 674666 584759 674672 584811
rect 43120 584685 43126 584737
rect 43178 584725 43184 584737
rect 47632 584725 47638 584737
rect 43178 584697 47638 584725
rect 43178 584685 43184 584697
rect 47632 584685 47638 584697
rect 47690 584685 47696 584737
rect 41776 584241 41782 584293
rect 41834 584281 41840 584293
rect 43216 584281 43222 584293
rect 41834 584253 43222 584281
rect 41834 584241 41840 584253
rect 43216 584241 43222 584253
rect 43274 584241 43280 584293
rect 41968 584167 41974 584219
rect 42026 584167 42032 584219
rect 42160 584167 42166 584219
rect 42218 584207 42224 584219
rect 43312 584207 43318 584219
rect 42218 584179 43318 584207
rect 42218 584167 42224 584179
rect 43312 584167 43318 584179
rect 43370 584167 43376 584219
rect 41986 583997 42014 584167
rect 41968 583945 41974 583997
rect 42026 583945 42032 583997
rect 671728 583353 671734 583405
rect 671786 583393 671792 583405
rect 671920 583393 671926 583405
rect 671786 583365 671926 583393
rect 671786 583353 671792 583365
rect 671920 583353 671926 583365
rect 671978 583393 671984 583405
rect 674608 583393 674614 583405
rect 671978 583365 674614 583393
rect 671978 583353 671984 583365
rect 674608 583353 674614 583365
rect 674666 583353 674672 583405
rect 672016 581873 672022 581925
rect 672074 581913 672080 581925
rect 673264 581913 673270 581925
rect 672074 581885 673270 581913
rect 672074 581873 672080 581885
rect 673264 581873 673270 581885
rect 673322 581873 673328 581925
rect 671920 581799 671926 581851
rect 671978 581839 671984 581851
rect 673840 581839 673846 581851
rect 671978 581811 673846 581839
rect 671978 581799 671984 581811
rect 673840 581799 673846 581811
rect 673898 581799 673904 581851
rect 43024 581503 43030 581555
rect 43082 581543 43088 581555
rect 43312 581543 43318 581555
rect 43082 581515 43318 581543
rect 43082 581503 43088 581515
rect 43312 581503 43318 581515
rect 43370 581503 43376 581555
rect 42064 581429 42070 581481
rect 42122 581469 42128 581481
rect 43120 581469 43126 581481
rect 42122 581441 43126 581469
rect 42122 581429 42128 581441
rect 43120 581429 43126 581441
rect 43178 581429 43184 581481
rect 42928 578395 42934 578447
rect 42986 578395 42992 578447
rect 42064 578247 42070 578299
rect 42122 578287 42128 578299
rect 42946 578287 42974 578395
rect 42122 578259 42974 578287
rect 42122 578247 42128 578259
rect 42160 577655 42166 577707
rect 42218 577695 42224 577707
rect 43024 577695 43030 577707
rect 42218 577667 43030 577695
rect 42218 577655 42224 577667
rect 43024 577655 43030 577667
rect 43082 577655 43088 577707
rect 654448 576027 654454 576079
rect 654506 576067 654512 576079
rect 672400 576067 672406 576079
rect 654506 576039 672406 576067
rect 654506 576027 654512 576039
rect 672400 576027 672406 576039
rect 672458 576027 672464 576079
rect 672688 575953 672694 576005
rect 672746 575993 672752 576005
rect 673840 575993 673846 576005
rect 672746 575965 673846 575993
rect 672746 575953 672752 575965
rect 673840 575953 673846 575965
rect 673898 575953 673904 576005
rect 672496 574325 672502 574377
rect 672554 574365 672560 574377
rect 674416 574365 674422 574377
rect 672554 574337 674422 574365
rect 672554 574325 672560 574337
rect 674416 574325 674422 574337
rect 674474 574325 674480 574377
rect 42160 574103 42166 574155
rect 42218 574143 42224 574155
rect 43120 574143 43126 574155
rect 42218 574115 43126 574143
rect 42218 574103 42224 574115
rect 43120 574103 43126 574115
rect 43178 574103 43184 574155
rect 42064 573215 42070 573267
rect 42122 573255 42128 573267
rect 42448 573255 42454 573267
rect 42122 573227 42454 573255
rect 42122 573215 42128 573227
rect 42448 573215 42454 573227
rect 42506 573215 42512 573267
rect 672880 573067 672886 573119
rect 672938 573107 672944 573119
rect 673840 573107 673846 573119
rect 672938 573079 673846 573107
rect 672938 573067 672944 573079
rect 673840 573067 673846 573079
rect 673898 573067 673904 573119
rect 672208 572845 672214 572897
rect 672266 572885 672272 572897
rect 674416 572885 674422 572897
rect 672266 572857 674422 572885
rect 672266 572845 672272 572857
rect 674416 572845 674422 572857
rect 674474 572845 674480 572897
rect 42160 572771 42166 572823
rect 42218 572811 42224 572823
rect 42928 572811 42934 572823
rect 42218 572783 42934 572811
rect 42218 572771 42224 572783
rect 42928 572771 42934 572783
rect 42986 572771 42992 572823
rect 42448 572623 42454 572675
rect 42506 572663 42512 572675
rect 42928 572663 42934 572675
rect 42506 572635 42934 572663
rect 42506 572623 42512 572635
rect 42928 572623 42934 572635
rect 42986 572623 42992 572675
rect 672784 571957 672790 572009
rect 672842 571997 672848 572009
rect 674416 571997 674422 572009
rect 672842 571969 674422 571997
rect 672842 571957 672848 571969
rect 674416 571957 674422 571969
rect 674474 571957 674480 572009
rect 42160 570995 42166 571047
rect 42218 571035 42224 571047
rect 43024 571035 43030 571047
rect 42218 571007 43030 571035
rect 42218 570995 42224 571007
rect 43024 570995 43030 571007
rect 43082 570995 43088 571047
rect 42160 570329 42166 570381
rect 42218 570369 42224 570381
rect 43120 570369 43126 570381
rect 42218 570341 43126 570369
rect 42218 570329 42224 570341
rect 43120 570329 43126 570341
rect 43178 570329 43184 570381
rect 42832 570255 42838 570307
rect 42890 570295 42896 570307
rect 59536 570295 59542 570307
rect 42890 570267 59542 570295
rect 42890 570255 42896 570267
rect 59536 570255 59542 570267
rect 59594 570255 59600 570307
rect 42064 569737 42070 569789
rect 42122 569777 42128 569789
rect 42928 569777 42934 569789
rect 42122 569749 42934 569777
rect 42122 569737 42128 569749
rect 42928 569737 42934 569749
rect 42986 569737 42992 569789
rect 650032 567369 650038 567421
rect 650090 567409 650096 567421
rect 679792 567409 679798 567421
rect 650090 567381 679798 567409
rect 650090 567369 650096 567381
rect 679792 567369 679798 567381
rect 679850 567369 679856 567421
rect 654352 567295 654358 567347
rect 654410 567335 654416 567347
rect 666640 567335 666646 567347
rect 654410 567307 666646 567335
rect 654410 567295 654416 567307
rect 666640 567295 666646 567307
rect 666698 567295 666704 567347
rect 34480 564483 34486 564535
rect 34538 564523 34544 564535
rect 51856 564523 51862 564535
rect 34538 564495 51862 564523
rect 34538 564483 34544 564495
rect 51856 564483 51862 564495
rect 51914 564483 51920 564535
rect 673744 564113 673750 564165
rect 673802 564153 673808 564165
rect 675088 564153 675094 564165
rect 673802 564125 675094 564153
rect 673802 564113 673808 564125
rect 675088 564113 675094 564125
rect 675146 564113 675152 564165
rect 42160 563447 42166 563499
rect 42218 563487 42224 563499
rect 48880 563487 48886 563499
rect 42218 563459 48886 563487
rect 42218 563447 42224 563459
rect 48880 563447 48886 563459
rect 48938 563447 48944 563499
rect 672304 563447 672310 563499
rect 672362 563487 672368 563499
rect 674992 563487 674998 563499
rect 672362 563459 674998 563487
rect 672362 563447 672368 563459
rect 674992 563447 674998 563459
rect 675050 563447 675056 563499
rect 51856 561523 51862 561575
rect 51914 561563 51920 561575
rect 59440 561563 59446 561575
rect 51914 561535 59446 561563
rect 51914 561523 51920 561535
rect 59440 561523 59446 561535
rect 59498 561523 59504 561575
rect 674704 559525 674710 559577
rect 674762 559565 674768 559577
rect 675376 559565 675382 559577
rect 674762 559537 675382 559565
rect 674762 559525 674768 559537
rect 675376 559525 675382 559537
rect 675434 559525 675440 559577
rect 675088 557823 675094 557875
rect 675146 557863 675152 557875
rect 675376 557863 675382 557875
rect 675146 557835 675382 557863
rect 675146 557823 675152 557835
rect 675376 557823 675382 557835
rect 675434 557823 675440 557875
rect 675088 557083 675094 557135
rect 675146 557123 675152 557135
rect 675472 557123 675478 557135
rect 675146 557095 675478 557123
rect 675146 557083 675152 557095
rect 675472 557083 675478 557095
rect 675530 557083 675536 557135
rect 660880 555825 660886 555877
rect 660938 555865 660944 555877
rect 674992 555865 674998 555877
rect 660938 555837 674998 555865
rect 660938 555825 660944 555837
rect 674992 555825 674998 555837
rect 675050 555825 675056 555877
rect 674224 555233 674230 555285
rect 674282 555273 674288 555285
rect 675472 555273 675478 555285
rect 674282 555245 675478 555273
rect 674282 555233 674288 555245
rect 675472 555233 675478 555245
rect 675530 555233 675536 555285
rect 674416 553753 674422 553805
rect 674474 553793 674480 553805
rect 675472 553793 675478 553805
rect 674474 553765 675478 553793
rect 674474 553753 674480 553765
rect 675472 553753 675478 553765
rect 675530 553753 675536 553805
rect 673744 553161 673750 553213
rect 673802 553201 673808 553213
rect 675376 553201 675382 553213
rect 673802 553173 675382 553201
rect 673802 553161 673808 553173
rect 675376 553161 675382 553173
rect 675434 553161 675440 553213
rect 654448 552939 654454 552991
rect 654506 552979 654512 552991
rect 663952 552979 663958 552991
rect 654506 552951 663958 552979
rect 654506 552939 654512 552951
rect 663952 552939 663958 552951
rect 664010 552939 664016 552991
rect 674320 551903 674326 551955
rect 674378 551943 674384 551955
rect 675472 551943 675478 551955
rect 674378 551915 675478 551943
rect 674378 551903 674384 551915
rect 675472 551903 675478 551915
rect 675530 551903 675536 551955
rect 674992 551607 674998 551659
rect 675050 551647 675056 551659
rect 675376 551647 675382 551659
rect 675050 551619 675382 551647
rect 675050 551607 675056 551619
rect 675376 551607 675382 551619
rect 675434 551607 675440 551659
rect 674992 550053 674998 550105
rect 675050 550093 675056 550105
rect 675472 550093 675478 550105
rect 675050 550065 675478 550093
rect 675050 550053 675056 550065
rect 675472 550053 675478 550065
rect 675530 550053 675536 550105
rect 674512 548203 674518 548255
rect 674570 548243 674576 548255
rect 675472 548243 675478 548255
rect 674570 548215 675478 548243
rect 674570 548203 674576 548215
rect 675472 548203 675478 548215
rect 675530 548203 675536 548255
rect 674032 546353 674038 546405
rect 674090 546393 674096 546405
rect 674320 546393 674326 546405
rect 674090 546365 674326 546393
rect 674090 546353 674096 546365
rect 674320 546353 674326 546365
rect 674378 546353 674384 546405
rect 43312 544799 43318 544851
rect 43370 544839 43376 544851
rect 44560 544839 44566 544851
rect 43370 544811 44566 544839
rect 43370 544799 43376 544811
rect 44560 544799 44566 544811
rect 44618 544799 44624 544851
rect 48880 544651 48886 544703
rect 48938 544691 48944 544703
rect 59536 544691 59542 544703
rect 48938 544663 59542 544691
rect 48938 544651 48944 544663
rect 59536 544651 59542 544663
rect 59594 544651 59600 544703
rect 41872 544503 41878 544555
rect 41930 544543 41936 544555
rect 42160 544543 42166 544555
rect 41930 544515 42166 544543
rect 41930 544503 41936 544515
rect 42160 544503 42166 544515
rect 42218 544503 42224 544555
rect 42160 544355 42166 544407
rect 42218 544395 42224 544407
rect 42448 544395 42454 544407
rect 42218 544367 42454 544395
rect 42218 544355 42224 544367
rect 42448 544355 42454 544367
rect 42506 544355 42512 544407
rect 40240 544207 40246 544259
rect 40298 544247 40304 544259
rect 41008 544247 41014 544259
rect 40298 544219 41014 544247
rect 40298 544207 40304 544219
rect 41008 544207 41014 544219
rect 41066 544207 41072 544259
rect 42928 541617 42934 541669
rect 42986 541657 42992 541669
rect 43312 541657 43318 541669
rect 42986 541629 43318 541657
rect 42986 541617 42992 541629
rect 43312 541617 43318 541629
rect 43370 541617 43376 541669
rect 654160 541543 654166 541595
rect 654218 541583 654224 541595
rect 661168 541583 661174 541595
rect 654218 541555 661174 541583
rect 654218 541543 654224 541555
rect 661168 541543 661174 541555
rect 661226 541543 661232 541595
rect 42928 541469 42934 541521
rect 42986 541509 42992 541521
rect 50512 541509 50518 541521
rect 42986 541481 50518 541509
rect 42986 541469 42992 541481
rect 50512 541469 50518 541481
rect 50570 541469 50576 541521
rect 655408 541469 655414 541521
rect 655466 541509 655472 541521
rect 674320 541509 674326 541521
rect 655466 541481 674326 541509
rect 655466 541469 655472 541481
rect 674320 541469 674326 541481
rect 674378 541469 674384 541521
rect 669808 541395 669814 541447
rect 669866 541435 669872 541447
rect 674608 541435 674614 541447
rect 669866 541407 674614 541435
rect 669866 541395 669872 541407
rect 674608 541395 674614 541407
rect 674666 541395 674672 541447
rect 41392 541321 41398 541373
rect 41450 541361 41456 541373
rect 43504 541361 43510 541373
rect 41450 541333 43510 541361
rect 41450 541321 41456 541333
rect 43504 541321 43510 541333
rect 43562 541321 43568 541373
rect 41968 540951 41974 541003
rect 42026 540951 42032 541003
rect 42064 540951 42070 541003
rect 42122 540991 42128 541003
rect 42448 540991 42454 541003
rect 42122 540963 42454 540991
rect 42122 540951 42128 540963
rect 42448 540951 42454 540963
rect 42506 540951 42512 541003
rect 41986 540781 42014 540951
rect 41968 540729 41974 540781
rect 42026 540729 42032 540781
rect 661072 540729 661078 540781
rect 661130 540769 661136 540781
rect 674608 540769 674614 540781
rect 661130 540741 674614 540769
rect 661130 540729 661136 540741
rect 674608 540729 674614 540741
rect 674666 540729 674672 540781
rect 671920 539841 671926 539893
rect 671978 539881 671984 539893
rect 674608 539881 674614 539893
rect 671978 539853 674614 539881
rect 671978 539841 671984 539853
rect 674608 539841 674614 539853
rect 674666 539841 674672 539893
rect 673936 539767 673942 539819
rect 673994 539807 674000 539819
rect 674224 539807 674230 539819
rect 673994 539779 674230 539807
rect 673994 539767 674000 539779
rect 674224 539767 674230 539779
rect 674282 539767 674288 539819
rect 674512 539249 674518 539301
rect 674570 539289 674576 539301
rect 675088 539289 675094 539301
rect 674570 539261 675094 539289
rect 674570 539249 674576 539261
rect 675088 539249 675094 539261
rect 675146 539249 675152 539301
rect 42160 538287 42166 538339
rect 42218 538327 42224 538339
rect 42928 538327 42934 538339
rect 42218 538299 42934 538327
rect 42218 538287 42224 538299
rect 42928 538287 42934 538299
rect 42986 538287 42992 538339
rect 42928 538139 42934 538191
rect 42986 538179 42992 538191
rect 43312 538179 43318 538191
rect 42986 538151 43318 538179
rect 42986 538139 42992 538151
rect 43312 538139 43318 538151
rect 43370 538139 43376 538191
rect 42064 535771 42070 535823
rect 42122 535811 42128 535823
rect 43024 535811 43030 535823
rect 42122 535783 43030 535811
rect 42122 535771 42128 535783
rect 43024 535771 43030 535783
rect 43082 535771 43088 535823
rect 43024 535623 43030 535675
rect 43082 535663 43088 535675
rect 43504 535663 43510 535675
rect 43082 535635 43510 535663
rect 43082 535623 43088 535635
rect 43504 535623 43510 535635
rect 43562 535623 43568 535675
rect 672016 535623 672022 535675
rect 672074 535663 672080 535675
rect 676624 535663 676630 535675
rect 672074 535635 676630 535663
rect 672074 535623 672080 535635
rect 676624 535623 676630 535635
rect 676682 535623 676688 535675
rect 671728 535549 671734 535601
rect 671786 535589 671792 535601
rect 676528 535589 676534 535601
rect 671786 535561 676534 535589
rect 671786 535549 671792 535561
rect 676528 535549 676534 535561
rect 676586 535549 676592 535601
rect 42160 534587 42166 534639
rect 42218 534627 42224 534639
rect 42928 534627 42934 534639
rect 42218 534599 42934 534627
rect 42218 534587 42224 534599
rect 42928 534587 42934 534599
rect 42986 534587 42992 534639
rect 42160 531479 42166 531531
rect 42218 531519 42224 531531
rect 42448 531519 42454 531531
rect 42218 531491 42454 531519
rect 42218 531479 42224 531491
rect 42448 531479 42454 531491
rect 42506 531479 42512 531531
rect 672976 531109 672982 531161
rect 673034 531149 673040 531161
rect 674800 531149 674806 531161
rect 673034 531121 674806 531149
rect 673034 531109 673040 531121
rect 674800 531109 674806 531121
rect 674858 531109 674864 531161
rect 42160 530887 42166 530939
rect 42218 530927 42224 530939
rect 43024 530927 43030 530939
rect 42218 530899 43030 530927
rect 42218 530887 42224 530899
rect 43024 530887 43030 530899
rect 43082 530887 43088 530939
rect 42064 530147 42070 530199
rect 42122 530187 42128 530199
rect 42928 530187 42934 530199
rect 42122 530159 42934 530187
rect 42122 530147 42128 530159
rect 42928 530147 42934 530159
rect 42986 530147 42992 530199
rect 43024 529925 43030 529977
rect 43082 529965 43088 529977
rect 59536 529965 59542 529977
rect 43082 529937 59542 529965
rect 43082 529925 43088 529937
rect 59536 529925 59542 529937
rect 59594 529925 59600 529977
rect 654064 529925 654070 529977
rect 654122 529965 654128 529977
rect 672496 529965 672502 529977
rect 654122 529937 672502 529965
rect 654122 529925 654128 529937
rect 672496 529925 672502 529937
rect 672554 529925 672560 529977
rect 674032 529925 674038 529977
rect 674090 529965 674096 529977
rect 674416 529965 674422 529977
rect 674090 529937 674422 529965
rect 674090 529925 674096 529937
rect 674416 529925 674422 529937
rect 674474 529925 674480 529977
rect 672112 529481 672118 529533
rect 672170 529521 672176 529533
rect 674800 529521 674806 529533
rect 672170 529493 674806 529521
rect 672170 529481 672176 529493
rect 674800 529481 674806 529493
rect 674858 529481 674864 529533
rect 42160 529407 42166 529459
rect 42218 529447 42224 529459
rect 42448 529447 42454 529459
rect 42218 529419 42454 529447
rect 42218 529407 42224 529419
rect 42448 529407 42454 529419
rect 42506 529407 42512 529459
rect 671824 528889 671830 528941
rect 671882 528929 671888 528941
rect 674800 528929 674806 528941
rect 671882 528901 674806 528929
rect 671882 528889 671888 528901
rect 674800 528889 674806 528901
rect 674858 528889 674864 528941
rect 671632 528001 671638 528053
rect 671690 528041 671696 528053
rect 674800 528041 674806 528053
rect 671690 528013 674806 528041
rect 671690 528001 671696 528013
rect 674800 528001 674806 528013
rect 674858 528001 674864 528053
rect 42160 527631 42166 527683
rect 42218 527671 42224 527683
rect 43120 527671 43126 527683
rect 42218 527643 43126 527671
rect 42218 527631 42224 527643
rect 43120 527631 43126 527643
rect 43178 527631 43184 527683
rect 42064 527187 42070 527239
rect 42122 527227 42128 527239
rect 42928 527227 42934 527239
rect 42122 527199 42934 527227
rect 42122 527187 42128 527199
rect 42928 527187 42934 527199
rect 42986 527187 42992 527239
rect 650128 521267 650134 521319
rect 650186 521307 650192 521319
rect 679792 521307 679798 521319
rect 650186 521279 679798 521307
rect 650186 521267 650192 521279
rect 679792 521267 679798 521279
rect 679850 521267 679856 521319
rect 41872 519787 41878 519839
rect 41930 519827 41936 519839
rect 43024 519827 43030 519839
rect 41930 519799 43030 519827
rect 41930 519787 41936 519799
rect 43024 519787 43030 519799
rect 43082 519787 43088 519839
rect 654064 519343 654070 519395
rect 654122 519383 654128 519395
rect 663856 519383 663862 519395
rect 654122 519355 663862 519383
rect 654122 519343 654128 519355
rect 663856 519343 663862 519355
rect 663914 519343 663920 519395
rect 53872 515495 53878 515547
rect 53930 515535 53936 515547
rect 59536 515535 59542 515547
rect 53930 515507 59542 515535
rect 53930 515495 53936 515507
rect 59536 515495 59542 515507
rect 59594 515495 59600 515547
rect 656368 506911 656374 506963
rect 656426 506951 656432 506963
rect 669520 506951 669526 506963
rect 656426 506923 669526 506951
rect 656426 506911 656432 506923
rect 669520 506911 669526 506923
rect 669578 506911 669584 506963
rect 47632 501139 47638 501191
rect 47690 501179 47696 501191
rect 59536 501179 59542 501191
rect 47690 501151 59542 501179
rect 47690 501139 47696 501151
rect 59536 501139 59542 501151
rect 59594 501139 59600 501191
rect 674416 497439 674422 497491
rect 674474 497479 674480 497491
rect 674896 497479 674902 497491
rect 674474 497451 674902 497479
rect 674474 497439 674480 497451
rect 674896 497439 674902 497451
rect 674954 497439 674960 497491
rect 672592 497291 672598 497343
rect 672650 497331 672656 497343
rect 674416 497331 674422 497343
rect 672650 497303 674422 497331
rect 672650 497291 672656 497303
rect 674416 497291 674422 497303
rect 674474 497291 674480 497343
rect 669712 496477 669718 496529
rect 669770 496517 669776 496529
rect 674416 496517 674422 496529
rect 669770 496489 674422 496517
rect 669770 496477 669776 496489
rect 674416 496477 674422 496489
rect 674474 496477 674480 496529
rect 655312 495515 655318 495567
rect 655370 495555 655376 495567
rect 674704 495555 674710 495567
rect 655370 495527 674710 495555
rect 655370 495515 655376 495527
rect 674704 495515 674710 495527
rect 674762 495515 674768 495567
rect 44752 486709 44758 486761
rect 44810 486749 44816 486761
rect 58576 486749 58582 486761
rect 44810 486721 58582 486749
rect 44810 486709 44816 486721
rect 58576 486709 58582 486721
rect 58634 486709 58640 486761
rect 654256 483823 654262 483875
rect 654314 483863 654320 483875
rect 666928 483863 666934 483875
rect 654314 483835 666934 483863
rect 654314 483823 654320 483835
rect 666928 483823 666934 483835
rect 666986 483823 666992 483875
rect 650224 478125 650230 478177
rect 650282 478165 650288 478177
rect 679792 478165 679798 478177
rect 650282 478137 679798 478165
rect 650282 478125 650288 478137
rect 679792 478125 679798 478137
rect 679850 478125 679856 478177
rect 44848 472353 44854 472405
rect 44906 472393 44912 472405
rect 59536 472393 59542 472405
rect 44906 472365 59542 472393
rect 44906 472353 44912 472365
rect 59536 472353 59542 472365
rect 59594 472353 59600 472405
rect 654448 472205 654454 472257
rect 654506 472245 654512 472257
rect 660976 472245 660982 472257
rect 654506 472217 660982 472245
rect 654506 472205 654512 472217
rect 660976 472205 660982 472217
rect 661034 472205 661040 472257
rect 50512 457923 50518 457975
rect 50570 457963 50576 457975
rect 59536 457963 59542 457975
rect 50570 457935 59542 457963
rect 50570 457923 50576 457935
rect 59536 457923 59542 457935
rect 59594 457923 59600 457975
rect 654448 457923 654454 457975
rect 654506 457963 654512 457975
rect 661072 457963 661078 457975
rect 654506 457935 661078 457963
rect 654506 457923 654512 457935
rect 661072 457923 661078 457935
rect 661130 457923 661136 457975
rect 654352 446379 654358 446431
rect 654410 446419 654416 446431
rect 663856 446419 663862 446431
rect 654410 446391 663862 446419
rect 654410 446379 654416 446391
rect 663856 446379 663862 446391
rect 663914 446379 663920 446431
rect 53968 443567 53974 443619
rect 54026 443607 54032 443619
rect 59536 443607 59542 443619
rect 54026 443579 59542 443607
rect 54026 443567 54032 443579
rect 59536 443567 59542 443579
rect 59594 443567 59600 443619
rect 42256 437129 42262 437181
rect 42314 437169 42320 437181
rect 53872 437169 53878 437181
rect 42314 437141 53878 437169
rect 42314 437129 42320 437141
rect 53872 437129 53878 437141
rect 53930 437129 53936 437181
rect 42256 436241 42262 436293
rect 42314 436281 42320 436293
rect 47632 436281 47638 436293
rect 42314 436253 47638 436281
rect 42314 436241 42320 436253
rect 47632 436241 47638 436253
rect 47690 436241 47696 436293
rect 654448 434909 654454 434961
rect 654506 434949 654512 434961
rect 664048 434949 664054 434961
rect 654506 434921 664054 434949
rect 654506 434909 654512 434921
rect 664048 434909 664054 434921
rect 664106 434909 664112 434961
rect 47632 429137 47638 429189
rect 47690 429177 47696 429189
rect 59536 429177 59542 429189
rect 47690 429149 59542 429177
rect 47690 429137 47696 429149
rect 59536 429137 59542 429149
rect 59594 429137 59600 429189
rect 654448 426177 654454 426229
rect 654506 426217 654512 426229
rect 669616 426217 669622 426229
rect 654506 426189 669622 426217
rect 654506 426177 654512 426189
rect 669616 426177 669622 426189
rect 669674 426177 669680 426229
rect 42352 418407 42358 418459
rect 42410 418447 42416 418459
rect 53872 418447 53878 418459
rect 42410 418419 53878 418447
rect 42410 418407 42416 418419
rect 53872 418407 53878 418419
rect 53930 418407 53936 418459
rect 37360 416483 37366 416535
rect 37418 416523 37424 416535
rect 42448 416523 42454 416535
rect 37418 416495 42454 416523
rect 37418 416483 37424 416495
rect 42448 416483 42454 416495
rect 42506 416483 42512 416535
rect 40240 415373 40246 415425
rect 40298 415413 40304 415425
rect 42928 415413 42934 415425
rect 40298 415385 42934 415413
rect 40298 415373 40304 415385
rect 42928 415373 42934 415385
rect 42986 415373 42992 415425
rect 40144 415151 40150 415203
rect 40202 415191 40208 415203
rect 43024 415191 43030 415203
rect 40202 415163 43030 415191
rect 40202 415151 40208 415163
rect 43024 415151 43030 415163
rect 43082 415151 43088 415203
rect 43216 414855 43222 414907
rect 43274 414895 43280 414907
rect 43696 414895 43702 414907
rect 43274 414867 43702 414895
rect 43274 414855 43280 414867
rect 43696 414855 43702 414867
rect 43754 414855 43760 414907
rect 37264 414707 37270 414759
rect 37322 414747 37328 414759
rect 43216 414747 43222 414759
rect 37322 414719 43222 414747
rect 37322 414707 37328 414719
rect 43216 414707 43222 414719
rect 43274 414707 43280 414759
rect 45040 414707 45046 414759
rect 45098 414747 45104 414759
rect 58384 414747 58390 414759
rect 45098 414719 58390 414747
rect 45098 414707 45104 414719
rect 58384 414707 58390 414719
rect 58442 414707 58448 414759
rect 41776 413375 41782 413427
rect 41834 413375 41840 413427
rect 41794 413205 41822 413375
rect 41776 413153 41782 413205
rect 41834 413153 41840 413205
rect 653872 411821 653878 411873
rect 653930 411861 653936 411873
rect 669616 411861 669622 411873
rect 653930 411833 669622 411861
rect 653930 411821 653936 411833
rect 669616 411821 669622 411833
rect 669674 411821 669680 411873
rect 42352 411451 42358 411503
rect 42410 411451 42416 411503
rect 42160 411303 42166 411355
rect 42218 411343 42224 411355
rect 42370 411343 42398 411451
rect 42218 411315 42398 411343
rect 42218 411303 42224 411315
rect 42544 409823 42550 409875
rect 42602 409863 42608 409875
rect 42602 409835 42974 409863
rect 42602 409823 42608 409835
rect 42160 409675 42166 409727
rect 42218 409715 42224 409727
rect 42544 409715 42550 409727
rect 42218 409687 42550 409715
rect 42218 409675 42224 409687
rect 42544 409675 42550 409687
rect 42602 409675 42608 409727
rect 42160 409453 42166 409505
rect 42218 409493 42224 409505
rect 42352 409493 42358 409505
rect 42218 409465 42358 409493
rect 42218 409453 42224 409465
rect 42352 409453 42358 409465
rect 42410 409453 42416 409505
rect 42946 409419 42974 409835
rect 42946 409391 43070 409419
rect 42352 409305 42358 409357
rect 42410 409345 42416 409357
rect 42928 409345 42934 409357
rect 42410 409317 42934 409345
rect 42410 409305 42416 409317
rect 42928 409305 42934 409317
rect 42986 409305 42992 409357
rect 42928 409157 42934 409209
rect 42986 409197 42992 409209
rect 43042 409197 43070 409391
rect 42986 409169 43070 409197
rect 42986 409157 42992 409169
rect 666832 409157 666838 409209
rect 666890 409197 666896 409209
rect 674416 409197 674422 409209
rect 666890 409169 674422 409197
rect 666890 409157 666896 409169
rect 674416 409157 674422 409169
rect 674474 409157 674480 409209
rect 655120 409083 655126 409135
rect 655178 409123 655184 409135
rect 674704 409123 674710 409135
rect 655178 409095 674710 409123
rect 655178 409083 655184 409095
rect 674704 409083 674710 409095
rect 674762 409083 674768 409135
rect 672400 408343 672406 408395
rect 672458 408383 672464 408395
rect 674704 408383 674710 408395
rect 672458 408355 674710 408383
rect 672458 408343 672464 408355
rect 674704 408343 674710 408355
rect 674762 408343 674768 408395
rect 42160 408195 42166 408247
rect 42218 408235 42224 408247
rect 43120 408235 43126 408247
rect 42218 408207 43126 408235
rect 42218 408195 42224 408207
rect 43120 408195 43126 408207
rect 43178 408195 43184 408247
rect 42064 407455 42070 407507
rect 42122 407495 42128 407507
rect 43024 407495 43030 407507
rect 42122 407467 43030 407495
rect 42122 407455 42128 407467
rect 43024 407455 43030 407467
rect 43082 407455 43088 407507
rect 42160 407011 42166 407063
rect 42218 407051 42224 407063
rect 42352 407051 42358 407063
rect 42218 407023 42358 407051
rect 42218 407011 42224 407023
rect 42352 407011 42358 407023
rect 42410 407011 42416 407063
rect 42544 406049 42550 406101
rect 42602 406089 42608 406101
rect 53392 406089 53398 406101
rect 42602 406061 53398 406089
rect 42602 406049 42608 406061
rect 53392 406049 53398 406061
rect 53450 406049 53456 406101
rect 42160 403829 42166 403881
rect 42218 403869 42224 403881
rect 43216 403869 43222 403881
rect 42218 403841 43222 403869
rect 42218 403829 42224 403841
rect 43216 403829 43222 403841
rect 43274 403829 43280 403881
rect 42160 403311 42166 403363
rect 42218 403351 42224 403363
rect 42928 403351 42934 403363
rect 42218 403323 42934 403351
rect 42218 403311 42224 403323
rect 42928 403311 42934 403323
rect 42986 403311 42992 403363
rect 56272 400351 56278 400403
rect 56330 400391 56336 400403
rect 57616 400391 57622 400403
rect 56330 400363 57622 400391
rect 56330 400351 56336 400363
rect 57616 400351 57622 400363
rect 57674 400351 57680 400403
rect 654448 400351 654454 400403
rect 654506 400391 654512 400403
rect 666640 400391 666646 400403
rect 654506 400363 666646 400391
rect 654506 400351 654512 400363
rect 666640 400351 666646 400363
rect 666698 400351 666704 400403
rect 42352 393913 42358 393965
rect 42410 393953 42416 393965
rect 44848 393953 44854 393965
rect 42410 393925 44854 393953
rect 42410 393913 42416 393925
rect 44848 393913 44854 393925
rect 44906 393913 44912 393965
rect 42640 392877 42646 392929
rect 42698 392917 42704 392929
rect 50512 392917 50518 392929
rect 42698 392889 50518 392917
rect 42698 392877 42704 392889
rect 50512 392877 50518 392889
rect 50570 392877 50576 392929
rect 42352 392285 42358 392337
rect 42410 392325 42416 392337
rect 44752 392325 44758 392337
rect 42410 392297 44758 392325
rect 42410 392285 42416 392297
rect 44752 392285 44758 392297
rect 44810 392285 44816 392337
rect 650320 391693 650326 391745
rect 650378 391733 650384 391745
rect 679696 391733 679702 391745
rect 650378 391705 679702 391733
rect 650378 391693 650384 391705
rect 679696 391693 679702 391705
rect 679754 391693 679760 391745
rect 654448 388807 654454 388859
rect 654506 388847 654512 388859
rect 669712 388847 669718 388859
rect 654506 388819 669718 388847
rect 654506 388807 654512 388819
rect 669712 388807 669718 388819
rect 669770 388807 669776 388859
rect 675376 386365 675382 386417
rect 675434 386365 675440 386417
rect 675394 386195 675422 386365
rect 675376 386143 675382 386195
rect 675434 386143 675440 386195
rect 44944 385921 44950 385973
rect 45002 385961 45008 385973
rect 59248 385961 59254 385973
rect 45002 385933 59254 385961
rect 45002 385921 45008 385933
rect 59248 385921 59254 385933
rect 59306 385921 59312 385973
rect 675184 385403 675190 385455
rect 675242 385443 675248 385455
rect 675472 385443 675478 385455
rect 675242 385415 675478 385443
rect 675242 385403 675248 385415
rect 675472 385403 675478 385415
rect 675530 385403 675536 385455
rect 674320 385107 674326 385159
rect 674378 385147 674384 385159
rect 675184 385147 675190 385159
rect 674378 385119 675190 385147
rect 674378 385107 674384 385119
rect 675184 385107 675190 385119
rect 675242 385107 675248 385159
rect 674032 384811 674038 384863
rect 674090 384851 674096 384863
rect 675376 384851 675382 384863
rect 674090 384823 675382 384851
rect 674090 384811 674096 384823
rect 675376 384811 675382 384823
rect 675434 384811 675440 384863
rect 673936 383109 673942 383161
rect 673994 383149 674000 383161
rect 675280 383149 675286 383161
rect 673994 383121 675286 383149
rect 673994 383109 674000 383121
rect 675280 383109 675286 383121
rect 675338 383109 675344 383161
rect 674608 382443 674614 382495
rect 674666 382483 674672 382495
rect 675472 382483 675478 382495
rect 674666 382455 675478 382483
rect 674666 382443 674672 382455
rect 675472 382443 675478 382455
rect 675530 382443 675536 382495
rect 654448 380075 654454 380127
rect 654506 380115 654512 380127
rect 666736 380115 666742 380127
rect 654506 380087 666742 380115
rect 654506 380075 654512 380087
rect 666736 380075 666742 380087
rect 666794 380075 666800 380127
rect 675088 378965 675094 379017
rect 675146 379005 675152 379017
rect 675280 379005 675286 379017
rect 675146 378977 675286 379005
rect 675146 378965 675152 378977
rect 675280 378965 675286 378977
rect 675338 378965 675344 379017
rect 674992 378151 674998 378203
rect 675050 378191 675056 378203
rect 675376 378191 675382 378203
rect 675050 378163 675382 378191
rect 675050 378151 675056 378163
rect 675376 378151 675382 378163
rect 675434 378151 675440 378203
rect 674896 377559 674902 377611
rect 674954 377599 674960 377611
rect 675376 377599 675382 377611
rect 674954 377571 675382 377599
rect 674954 377559 674960 377571
rect 675376 377559 675382 377571
rect 675434 377559 675440 377611
rect 674704 376819 674710 376871
rect 674762 376859 674768 376871
rect 675472 376859 675478 376871
rect 674762 376831 675478 376859
rect 674762 376819 674768 376831
rect 675472 376819 675478 376831
rect 675530 376819 675536 376871
rect 674128 375709 674134 375761
rect 674186 375749 674192 375761
rect 675472 375749 675478 375761
rect 674186 375721 675478 375749
rect 674186 375709 674192 375721
rect 675472 375709 675478 375721
rect 675530 375709 675536 375761
rect 42256 375191 42262 375243
rect 42314 375231 42320 375243
rect 44752 375231 44758 375243
rect 42314 375203 44758 375231
rect 42314 375191 42320 375203
rect 44752 375191 44758 375203
rect 44810 375191 44816 375243
rect 37360 373193 37366 373245
rect 37418 373233 37424 373245
rect 43312 373233 43318 373245
rect 37418 373205 43318 373233
rect 37418 373193 37424 373205
rect 43312 373193 43318 373205
rect 43370 373193 43376 373245
rect 40048 373045 40054 373097
rect 40106 373085 40112 373097
rect 43024 373085 43030 373097
rect 40106 373057 43030 373085
rect 40106 373045 40112 373057
rect 43024 373045 43030 373057
rect 43082 373045 43088 373097
rect 40144 372527 40150 372579
rect 40202 372567 40208 372579
rect 42832 372567 42838 372579
rect 40202 372539 42838 372567
rect 40202 372527 40208 372539
rect 42832 372527 42838 372539
rect 42890 372527 42896 372579
rect 40240 372231 40246 372283
rect 40298 372271 40304 372283
rect 42928 372271 42934 372283
rect 40298 372243 42934 372271
rect 40298 372231 40304 372243
rect 42928 372231 42934 372243
rect 42986 372231 42992 372283
rect 37264 371565 37270 371617
rect 37322 371605 37328 371617
rect 38320 371605 38326 371617
rect 37322 371577 38326 371605
rect 37322 371565 37328 371577
rect 38320 371565 38326 371577
rect 38378 371565 38384 371617
rect 47728 371565 47734 371617
rect 47786 371605 47792 371617
rect 59536 371605 59542 371617
rect 47786 371577 59542 371605
rect 47786 371565 47792 371577
rect 59536 371565 59542 371577
rect 59594 371565 59600 371617
rect 41968 370159 41974 370211
rect 42026 370159 42032 370211
rect 41986 369829 42014 370159
rect 42160 369937 42166 369989
rect 42218 369977 42224 369989
rect 42352 369977 42358 369989
rect 42218 369949 42358 369977
rect 42218 369937 42224 369949
rect 42352 369937 42358 369949
rect 42410 369937 42416 369989
rect 42352 369829 42358 369841
rect 41986 369801 42358 369829
rect 42352 369789 42358 369801
rect 42410 369789 42416 369841
rect 42064 368087 42070 368139
rect 42122 368127 42128 368139
rect 42352 368127 42358 368139
rect 42122 368099 42358 368127
rect 42122 368087 42128 368099
rect 42352 368087 42358 368099
rect 42410 368087 42416 368139
rect 42064 367347 42070 367399
rect 42122 367387 42128 367399
rect 47440 367387 47446 367399
rect 42122 367359 47446 367387
rect 42122 367347 42128 367359
rect 47440 367347 47446 367359
rect 47498 367347 47504 367399
rect 42064 366237 42070 366289
rect 42122 366277 42128 366289
rect 42832 366277 42838 366289
rect 42122 366249 42838 366277
rect 42122 366237 42128 366249
rect 42832 366237 42838 366249
rect 42890 366237 42896 366289
rect 654448 365793 654454 365845
rect 654506 365833 654512 365845
rect 660976 365833 660982 365845
rect 654506 365805 660982 365833
rect 654506 365793 654512 365805
rect 660976 365793 660982 365805
rect 661034 365793 661040 365845
rect 42160 364979 42166 365031
rect 42218 365019 42224 365031
rect 43120 365019 43126 365031
rect 42218 364991 43126 365019
rect 42218 364979 42224 364991
rect 43120 364979 43126 364991
rect 43178 364979 43184 365031
rect 661168 364905 661174 364957
rect 661226 364945 661232 364957
rect 674704 364945 674710 364957
rect 661226 364917 674710 364945
rect 661226 364905 661232 364917
rect 674704 364905 674710 364917
rect 674762 364905 674768 364957
rect 42064 364239 42070 364291
rect 42122 364279 42128 364291
rect 43024 364279 43030 364291
rect 42122 364251 43030 364279
rect 42122 364239 42128 364251
rect 43024 364239 43030 364251
rect 43082 364239 43088 364291
rect 663952 363869 663958 363921
rect 664010 363909 664016 363921
rect 674416 363909 674422 363921
rect 664010 363881 674422 363909
rect 664010 363869 664016 363881
rect 674416 363869 674422 363881
rect 674474 363869 674480 363921
rect 42160 363647 42166 363699
rect 42218 363687 42224 363699
rect 42928 363687 42934 363699
rect 42218 363659 42934 363687
rect 42218 363647 42224 363659
rect 42928 363647 42934 363659
rect 42986 363647 42992 363699
rect 672496 363277 672502 363329
rect 672554 363317 672560 363329
rect 674704 363317 674710 363329
rect 672554 363289 674710 363317
rect 672554 363277 672560 363289
rect 674704 363277 674710 363289
rect 674762 363277 674768 363329
rect 42160 360613 42166 360665
rect 42218 360653 42224 360665
rect 43312 360653 43318 360665
rect 42218 360625 43318 360653
rect 42218 360613 42224 360625
rect 43312 360613 43318 360625
rect 43370 360613 43376 360665
rect 56176 357357 56182 357409
rect 56234 357397 56240 357409
rect 60208 357397 60214 357409
rect 56234 357369 60214 357397
rect 56234 357357 56240 357369
rect 60208 357357 60214 357369
rect 60266 357357 60272 357409
rect 42352 350697 42358 350749
rect 42410 350737 42416 350749
rect 47632 350737 47638 350749
rect 42410 350709 47638 350737
rect 42410 350697 42416 350709
rect 47632 350697 47638 350709
rect 47690 350697 47696 350749
rect 42352 349957 42358 350009
rect 42410 349997 42416 350009
rect 45040 349997 45046 350009
rect 42410 349969 45046 349997
rect 42410 349957 42416 349969
rect 45040 349957 45046 349969
rect 45098 349957 45104 350009
rect 42352 349069 42358 349121
rect 42410 349109 42416 349121
rect 53968 349109 53974 349121
rect 42410 349081 53974 349109
rect 42410 349069 42416 349081
rect 53968 349069 53974 349081
rect 54026 349069 54032 349121
rect 650416 345591 650422 345643
rect 650474 345631 650480 345643
rect 679792 345631 679798 345643
rect 650474 345603 679798 345631
rect 650474 345591 650480 345603
rect 679792 345591 679798 345603
rect 679850 345591 679856 345643
rect 674704 344407 674710 344459
rect 674762 344447 674768 344459
rect 676816 344447 676822 344459
rect 674762 344419 676822 344447
rect 674762 344407 674768 344419
rect 676816 344407 676822 344419
rect 676874 344407 676880 344459
rect 50512 342779 50518 342831
rect 50570 342819 50576 342831
rect 58384 342819 58390 342831
rect 50570 342791 58390 342819
rect 50570 342779 50576 342791
rect 58384 342779 58390 342791
rect 58442 342779 58448 342831
rect 654448 342705 654454 342757
rect 654506 342745 654512 342757
rect 666736 342745 666742 342757
rect 654506 342717 666742 342745
rect 654506 342705 654512 342717
rect 666736 342705 666742 342717
rect 666794 342705 666800 342757
rect 674608 340929 674614 340981
rect 674666 340969 674672 340981
rect 675472 340969 675478 340981
rect 674666 340941 675478 340969
rect 674666 340929 674672 340941
rect 675472 340929 675478 340941
rect 675530 340929 675536 340981
rect 673936 339523 673942 339575
rect 673994 339563 674000 339575
rect 675376 339563 675382 339575
rect 673994 339535 675382 339563
rect 673994 339523 674000 339535
rect 675376 339523 675382 339535
rect 675434 339523 675440 339575
rect 674320 336563 674326 336615
rect 674378 336603 674384 336615
rect 675376 336603 675382 336615
rect 674378 336575 675382 336603
rect 674378 336563 674384 336575
rect 675376 336563 675382 336575
rect 675434 336563 675440 336615
rect 674032 332715 674038 332767
rect 674090 332755 674096 332767
rect 675376 332755 675382 332767
rect 674090 332727 675382 332755
rect 674090 332715 674096 332727
rect 675376 332715 675382 332727
rect 675434 332715 675440 332767
rect 674224 332345 674230 332397
rect 674282 332385 674288 332397
rect 675472 332385 675478 332397
rect 674282 332357 675478 332385
rect 674282 332345 674288 332357
rect 675472 332345 675478 332357
rect 675530 332345 675536 332397
rect 654448 332271 654454 332323
rect 654506 332311 654512 332323
rect 663760 332311 663766 332323
rect 654506 332283 663766 332311
rect 654506 332271 654512 332283
rect 663760 332271 663766 332283
rect 663818 332271 663824 332323
rect 42256 331975 42262 332027
rect 42314 332015 42320 332027
rect 45040 332015 45046 332027
rect 42314 331987 45046 332015
rect 42314 331975 42320 331987
rect 45040 331975 45046 331987
rect 45098 331975 45104 332027
rect 674128 331531 674134 331583
rect 674186 331571 674192 331583
rect 675376 331571 675382 331583
rect 674186 331543 675382 331571
rect 674186 331531 674192 331543
rect 675376 331531 675382 331543
rect 675434 331531 675440 331583
rect 41872 330643 41878 330695
rect 41930 330683 41936 330695
rect 42544 330683 42550 330695
rect 41930 330655 42550 330683
rect 41930 330643 41936 330655
rect 42544 330643 42550 330655
rect 42602 330643 42608 330695
rect 674704 330495 674710 330547
rect 674762 330535 674768 330547
rect 675472 330535 675478 330547
rect 674762 330507 675478 330535
rect 674762 330495 674768 330507
rect 675472 330495 675478 330507
rect 675530 330495 675536 330547
rect 37168 329755 37174 329807
rect 37226 329795 37232 329807
rect 43120 329795 43126 329807
rect 37226 329767 43126 329795
rect 37226 329755 37232 329767
rect 43120 329755 43126 329767
rect 43178 329755 43184 329807
rect 40048 328793 40054 328845
rect 40106 328833 40112 328845
rect 42928 328833 42934 328845
rect 40106 328805 42934 328833
rect 40106 328793 40112 328805
rect 42928 328793 42934 328805
rect 42986 328793 42992 328845
rect 39952 328497 39958 328549
rect 40010 328537 40016 328549
rect 43312 328537 43318 328549
rect 40010 328509 43318 328537
rect 40010 328497 40016 328509
rect 43312 328497 43318 328509
rect 43370 328497 43376 328549
rect 37360 328423 37366 328475
rect 37418 328463 37424 328475
rect 43024 328463 43030 328475
rect 37418 328435 43030 328463
rect 37418 328423 37424 328435
rect 43024 328423 43030 328435
rect 43082 328423 43088 328475
rect 40240 328349 40246 328401
rect 40298 328389 40304 328401
rect 42832 328389 42838 328401
rect 40298 328361 42838 328389
rect 40298 328349 40304 328361
rect 42832 328349 42838 328361
rect 42890 328349 42896 328401
rect 53392 328349 53398 328401
rect 53450 328389 53456 328401
rect 57808 328389 57814 328401
rect 53450 328361 57814 328389
rect 53450 328349 53456 328361
rect 57808 328349 57814 328361
rect 57866 328349 57872 328401
rect 41776 327017 41782 327069
rect 41834 327017 41840 327069
rect 41794 326773 41822 327017
rect 41776 326721 41782 326773
rect 41834 326721 41840 326773
rect 42064 324871 42070 324923
rect 42122 324911 42128 324923
rect 42544 324911 42550 324923
rect 42122 324883 42550 324911
rect 42122 324871 42128 324883
rect 42544 324871 42550 324883
rect 42602 324871 42608 324923
rect 42160 324131 42166 324183
rect 42218 324171 42224 324183
rect 50320 324171 50326 324183
rect 42218 324143 50326 324171
rect 42218 324131 42224 324143
rect 50320 324131 50326 324143
rect 50378 324131 50384 324183
rect 42160 323095 42166 323147
rect 42218 323135 42224 323147
rect 43120 323135 43126 323147
rect 42218 323107 43126 323135
rect 42218 323095 42224 323107
rect 43120 323095 43126 323107
rect 43178 323095 43184 323147
rect 42064 321763 42070 321815
rect 42122 321803 42128 321815
rect 42544 321803 42550 321815
rect 42122 321775 42550 321803
rect 42122 321763 42128 321775
rect 42544 321763 42550 321775
rect 42602 321763 42608 321815
rect 42160 321023 42166 321075
rect 42218 321063 42224 321075
rect 42928 321063 42934 321075
rect 42218 321035 42934 321063
rect 42218 321023 42224 321035
rect 42928 321023 42934 321035
rect 42986 321023 42992 321075
rect 42928 320875 42934 320927
rect 42986 320915 42992 320927
rect 43312 320915 43318 320927
rect 42986 320887 43318 320915
rect 42986 320875 42992 320887
rect 43312 320875 43318 320887
rect 43370 320875 43376 320927
rect 42160 320579 42166 320631
rect 42218 320619 42224 320631
rect 42832 320619 42838 320631
rect 42218 320591 42838 320619
rect 42218 320579 42224 320591
rect 42832 320579 42838 320591
rect 42890 320579 42896 320631
rect 655216 319691 655222 319743
rect 655274 319731 655280 319743
rect 674416 319731 674422 319743
rect 655274 319703 674422 319731
rect 655274 319691 655280 319703
rect 674416 319691 674422 319703
rect 674474 319691 674480 319743
rect 669520 318877 669526 318929
rect 669578 318917 669584 318929
rect 674416 318917 674422 318929
rect 669578 318889 674422 318917
rect 669578 318877 669584 318889
rect 674416 318877 674422 318889
rect 674474 318877 674480 318929
rect 42256 318729 42262 318781
rect 42314 318769 42320 318781
rect 43024 318769 43030 318781
rect 42314 318741 43030 318769
rect 42314 318729 42320 318741
rect 43024 318729 43030 318741
rect 43082 318729 43088 318781
rect 666928 318285 666934 318337
rect 666986 318325 666992 318337
rect 674704 318325 674710 318337
rect 666986 318297 674710 318325
rect 666986 318285 666992 318297
rect 674704 318285 674710 318297
rect 674762 318285 674768 318337
rect 42064 316583 42070 316635
rect 42122 316623 42128 316635
rect 42928 316623 42934 316635
rect 42122 316595 42934 316623
rect 42122 316583 42128 316595
rect 42928 316583 42934 316595
rect 42986 316583 42992 316635
rect 44848 313919 44854 313971
rect 44906 313959 44912 313971
rect 58000 313959 58006 313971
rect 44906 313931 58006 313959
rect 44906 313919 44912 313931
rect 58000 313919 58006 313931
rect 58058 313919 58064 313971
rect 42352 307481 42358 307533
rect 42410 307521 42416 307533
rect 44944 307521 44950 307533
rect 42410 307493 44950 307521
rect 42410 307481 42416 307493
rect 44944 307481 44950 307493
rect 45002 307481 45008 307533
rect 42352 306741 42358 306793
rect 42410 306781 42416 306793
rect 47728 306781 47734 306793
rect 42410 306753 47734 306781
rect 42410 306741 42416 306753
rect 47728 306741 47734 306753
rect 47786 306741 47792 306793
rect 42352 305483 42358 305535
rect 42410 305523 42416 305535
rect 56272 305523 56278 305535
rect 42410 305495 56278 305523
rect 42410 305483 42416 305495
rect 56272 305483 56278 305495
rect 56330 305483 56336 305535
rect 44944 299563 44950 299615
rect 45002 299603 45008 299615
rect 59440 299603 59446 299615
rect 45002 299575 59446 299603
rect 45002 299563 45008 299575
rect 59440 299563 59446 299575
rect 59498 299563 59504 299615
rect 650512 299563 650518 299615
rect 650570 299603 650576 299615
rect 679792 299603 679798 299615
rect 650570 299575 679798 299603
rect 650570 299563 650576 299575
rect 679792 299563 679798 299575
rect 679850 299563 679856 299615
rect 674704 299489 674710 299541
rect 674762 299529 674768 299541
rect 676816 299529 676822 299541
rect 674762 299501 676822 299529
rect 674762 299489 674768 299501
rect 676816 299489 676822 299501
rect 676874 299489 676880 299541
rect 674800 299415 674806 299467
rect 674858 299455 674864 299467
rect 676912 299455 676918 299467
rect 674858 299427 676918 299455
rect 674858 299415 674864 299427
rect 676912 299415 676918 299427
rect 676970 299415 676976 299467
rect 674032 294753 674038 294805
rect 674090 294793 674096 294805
rect 675184 294793 675190 294805
rect 674090 294765 675190 294793
rect 674090 294753 674096 294765
rect 675184 294753 675190 294765
rect 675242 294753 675248 294805
rect 674224 294235 674230 294287
rect 674282 294275 674288 294287
rect 675088 294275 675094 294287
rect 674282 294247 675094 294275
rect 674282 294235 674288 294247
rect 675088 294235 675094 294247
rect 675146 294235 675152 294287
rect 673936 292903 673942 292955
rect 673994 292943 674000 292955
rect 675376 292943 675382 292955
rect 673994 292915 675382 292943
rect 673994 292903 674000 292915
rect 675376 292903 675382 292915
rect 675434 292903 675440 292955
rect 674608 291719 674614 291771
rect 674666 291759 674672 291771
rect 675088 291759 675094 291771
rect 674666 291731 675094 291759
rect 674666 291719 674672 291731
rect 675088 291719 675094 291731
rect 675146 291719 675152 291771
rect 674320 291053 674326 291105
rect 674378 291093 674384 291105
rect 675088 291093 675094 291105
rect 674378 291065 675094 291093
rect 674378 291053 674384 291065
rect 675088 291053 675094 291065
rect 675146 291053 675152 291105
rect 41776 289795 41782 289847
rect 41834 289835 41840 289847
rect 42256 289835 42262 289847
rect 41834 289807 42262 289835
rect 41834 289795 41840 289807
rect 42256 289795 42262 289807
rect 42314 289795 42320 289847
rect 674800 288537 674806 288589
rect 674858 288577 674864 288589
rect 675472 288577 675478 288589
rect 674858 288549 675478 288577
rect 674858 288537 674864 288549
rect 675472 288537 675478 288549
rect 675530 288537 675536 288589
rect 42256 288019 42262 288071
rect 42314 288059 42320 288071
rect 56272 288059 56278 288071
rect 42314 288031 56278 288059
rect 42314 288019 42320 288031
rect 56272 288019 56278 288031
rect 56330 288019 56336 288071
rect 674416 287723 674422 287775
rect 674474 287763 674480 287775
rect 675376 287763 675382 287775
rect 674474 287735 675382 287763
rect 674474 287723 674480 287735
rect 675376 287723 675382 287735
rect 675434 287723 675440 287775
rect 674704 287353 674710 287405
rect 674762 287393 674768 287405
rect 675472 287393 675478 287405
rect 674762 287365 675478 287393
rect 674762 287353 674768 287365
rect 675472 287353 675478 287365
rect 675530 287353 675536 287405
rect 37264 286761 37270 286813
rect 37322 286801 37328 286813
rect 40528 286801 40534 286813
rect 37322 286773 40534 286801
rect 37322 286761 37328 286773
rect 40528 286761 40534 286773
rect 40586 286761 40592 286813
rect 674128 286539 674134 286591
rect 674186 286579 674192 286591
rect 675376 286579 675382 286591
rect 674186 286551 675382 286579
rect 674186 286539 674192 286551
rect 675376 286539 675382 286551
rect 675434 286539 675440 286591
rect 40048 285281 40054 285333
rect 40106 285321 40112 285333
rect 42256 285321 42262 285333
rect 40106 285293 42262 285321
rect 40106 285281 40112 285293
rect 42256 285281 42262 285293
rect 42314 285281 42320 285333
rect 40144 285207 40150 285259
rect 40202 285247 40208 285259
rect 43120 285247 43126 285259
rect 40202 285219 43126 285247
rect 40202 285207 40208 285219
rect 43120 285207 43126 285219
rect 43178 285207 43184 285259
rect 40240 285133 40246 285185
rect 40298 285173 40304 285185
rect 43024 285173 43030 285185
rect 40298 285145 43030 285173
rect 40298 285133 40304 285145
rect 43024 285133 43030 285145
rect 43082 285133 43088 285185
rect 45136 285133 45142 285185
rect 45194 285173 45200 285185
rect 58096 285173 58102 285185
rect 45194 285145 58102 285173
rect 45194 285133 45200 285145
rect 58096 285133 58102 285145
rect 58154 285133 58160 285185
rect 654448 284911 654454 284963
rect 654506 284951 654512 284963
rect 660880 284951 660886 284963
rect 654506 284923 660886 284951
rect 654506 284911 654512 284923
rect 660880 284911 660886 284923
rect 660938 284911 660944 284963
rect 41776 283801 41782 283853
rect 41834 283801 41840 283853
rect 41794 283557 41822 283801
rect 41776 283505 41782 283557
rect 41834 283505 41840 283557
rect 42160 281729 42166 281781
rect 42218 281769 42224 281781
rect 42352 281769 42358 281781
rect 42218 281741 42358 281769
rect 42218 281729 42224 281741
rect 42352 281729 42358 281741
rect 42410 281729 42416 281781
rect 42064 280101 42070 280153
rect 42122 280141 42128 280153
rect 42352 280141 42358 280153
rect 42122 280113 42358 280141
rect 42122 280101 42128 280113
rect 42352 280101 42358 280113
rect 42410 280101 42416 280153
rect 350338 278633 393854 278661
rect 42160 278547 42166 278599
rect 42218 278587 42224 278599
rect 42928 278587 42934 278599
rect 42218 278559 42934 278587
rect 42218 278547 42224 278559
rect 42928 278547 42934 278559
rect 42986 278547 42992 278599
rect 64912 278547 64918 278599
rect 64970 278587 64976 278599
rect 67600 278587 67606 278599
rect 64970 278559 67606 278587
rect 64970 278547 64976 278559
rect 67600 278547 67606 278559
rect 67658 278547 67664 278599
rect 299248 278547 299254 278599
rect 299306 278587 299312 278599
rect 299488 278587 299494 278599
rect 299306 278559 299494 278587
rect 299306 278547 299312 278559
rect 299488 278547 299494 278559
rect 299546 278547 299552 278599
rect 350338 278525 350366 278633
rect 393826 278599 393854 278633
rect 407554 278633 432446 278661
rect 407554 278599 407582 278633
rect 432418 278599 432446 278633
rect 384400 278587 384406 278599
rect 350434 278559 384406 278587
rect 226672 278473 226678 278525
rect 226730 278513 226736 278525
rect 329776 278513 329782 278525
rect 226730 278485 329782 278513
rect 226730 278473 226736 278485
rect 329776 278473 329782 278485
rect 329834 278473 329840 278525
rect 350320 278473 350326 278525
rect 350378 278473 350384 278525
rect 219568 278399 219574 278451
rect 219626 278439 219632 278451
rect 326512 278439 326518 278451
rect 219626 278411 326518 278439
rect 219626 278399 219632 278411
rect 326512 278399 326518 278411
rect 326570 278399 326576 278451
rect 339856 278399 339862 278451
rect 339914 278439 339920 278451
rect 350434 278439 350462 278559
rect 384400 278547 384406 278559
rect 384458 278547 384464 278599
rect 393808 278547 393814 278599
rect 393866 278547 393872 278599
rect 407536 278547 407542 278599
rect 407594 278547 407600 278599
rect 432400 278547 432406 278599
rect 432458 278547 432464 278599
rect 351760 278473 351766 278525
rect 351818 278513 351824 278525
rect 372496 278513 372502 278525
rect 351818 278485 372502 278513
rect 351818 278473 351824 278485
rect 372496 278473 372502 278485
rect 372554 278473 372560 278525
rect 372880 278473 372886 278525
rect 372938 278513 372944 278525
rect 374608 278513 374614 278525
rect 372938 278485 374614 278513
rect 372938 278473 372944 278485
rect 374608 278473 374614 278485
rect 374666 278473 374672 278525
rect 374704 278473 374710 278525
rect 374762 278513 374768 278525
rect 374762 278485 402974 278513
rect 374762 278473 374768 278485
rect 339914 278411 350462 278439
rect 339914 278399 339920 278411
rect 366352 278399 366358 278451
rect 366410 278439 366416 278451
rect 378352 278439 378358 278451
rect 366410 278411 378358 278439
rect 366410 278399 366416 278411
rect 378352 278399 378358 278411
rect 378410 278399 378416 278451
rect 380176 278439 380182 278451
rect 378466 278411 380182 278439
rect 292048 278325 292054 278377
rect 292106 278365 292112 278377
rect 374800 278365 374806 278377
rect 292106 278337 374806 278365
rect 292106 278325 292112 278337
rect 374800 278325 374806 278337
rect 374858 278325 374864 278377
rect 375280 278325 375286 278377
rect 375338 278365 375344 278377
rect 378466 278365 378494 278411
rect 380176 278399 380182 278411
rect 380234 278399 380240 278451
rect 380272 278399 380278 278451
rect 380330 278439 380336 278451
rect 400912 278439 400918 278451
rect 380330 278411 400918 278439
rect 380330 278399 380336 278411
rect 400912 278399 400918 278411
rect 400970 278399 400976 278451
rect 402946 278439 402974 278485
rect 408112 278439 408118 278451
rect 402946 278411 408118 278439
rect 408112 278399 408118 278411
rect 408170 278399 408176 278451
rect 375338 278337 378494 278365
rect 375338 278325 375344 278337
rect 378544 278325 378550 278377
rect 378602 278365 378608 278377
rect 384688 278365 384694 278377
rect 378602 278337 384694 278365
rect 378602 278325 378608 278337
rect 384688 278325 384694 278337
rect 384746 278325 384752 278377
rect 302800 278251 302806 278303
rect 302858 278291 302864 278303
rect 460432 278291 460438 278303
rect 302858 278263 460438 278291
rect 302858 278251 302864 278263
rect 460432 278251 460438 278263
rect 460490 278251 460496 278303
rect 293200 278177 293206 278229
rect 293258 278217 293264 278229
rect 382000 278217 382006 278229
rect 293258 278189 382006 278217
rect 293258 278177 293264 278189
rect 382000 278177 382006 278189
rect 382058 278177 382064 278229
rect 382384 278177 382390 278229
rect 382442 278217 382448 278229
rect 384016 278217 384022 278229
rect 382442 278189 384022 278217
rect 382442 278177 382448 278189
rect 384016 278177 384022 278189
rect 384074 278177 384080 278229
rect 384400 278177 384406 278229
rect 384458 278217 384464 278229
rect 407536 278217 407542 278229
rect 384458 278189 407542 278217
rect 384458 278177 384464 278189
rect 407536 278177 407542 278189
rect 407594 278177 407600 278229
rect 300784 278103 300790 278155
rect 300842 278143 300848 278155
rect 446320 278143 446326 278155
rect 300842 278115 446326 278143
rect 300842 278103 300848 278115
rect 446320 278103 446326 278115
rect 446378 278103 446384 278155
rect 301840 278029 301846 278081
rect 301898 278069 301904 278081
rect 453232 278069 453238 278081
rect 301898 278041 453238 278069
rect 301898 278029 301904 278041
rect 453232 278029 453238 278041
rect 453290 278029 453296 278081
rect 291664 277955 291670 278007
rect 291722 277995 291728 278007
rect 371344 277995 371350 278007
rect 291722 277967 371350 277995
rect 291722 277955 291728 277967
rect 371344 277955 371350 277967
rect 371402 277955 371408 278007
rect 371920 277955 371926 278007
rect 371978 277995 371984 278007
rect 397360 277995 397366 278007
rect 371978 277967 397366 277995
rect 371978 277955 371984 277967
rect 397360 277955 397366 277967
rect 397418 277955 397424 278007
rect 64816 277881 64822 277933
rect 64874 277921 64880 277933
rect 191440 277921 191446 277933
rect 64874 277893 191446 277921
rect 64874 277881 64880 277893
rect 191440 277881 191446 277893
rect 191498 277881 191504 277933
rect 287728 277881 287734 277933
rect 287786 277921 287792 277933
rect 339088 277921 339094 277933
rect 287786 277893 339094 277921
rect 287786 277881 287792 277893
rect 339088 277881 339094 277893
rect 339146 277881 339152 277933
rect 352912 277881 352918 277933
rect 352970 277921 352976 277933
rect 415312 277921 415318 277933
rect 352970 277893 415318 277921
rect 352970 277881 352976 277893
rect 415312 277881 415318 277893
rect 415370 277881 415376 277933
rect 569872 277881 569878 277933
rect 569930 277921 569936 277933
rect 649456 277921 649462 277933
rect 569930 277893 649462 277921
rect 569930 277881 569936 277893
rect 649456 277881 649462 277893
rect 649514 277881 649520 277933
rect 42160 277807 42166 277859
rect 42218 277847 42224 277859
rect 43120 277847 43126 277859
rect 42218 277819 43126 277847
rect 42218 277807 42224 277819
rect 43120 277807 43126 277819
rect 43178 277807 43184 277859
rect 283792 277807 283798 277859
rect 283850 277847 283856 277859
rect 336304 277847 336310 277859
rect 283850 277819 336310 277847
rect 283850 277807 283856 277819
rect 336304 277807 336310 277819
rect 336362 277807 336368 277859
rect 354448 277807 354454 277859
rect 354506 277847 354512 277859
rect 429520 277847 429526 277859
rect 354506 277819 429526 277847
rect 354506 277807 354512 277819
rect 429520 277807 429526 277819
rect 429578 277807 429584 277859
rect 288400 277733 288406 277785
rect 288458 277773 288464 277785
rect 342736 277773 342742 277785
rect 288458 277745 342742 277773
rect 288458 277733 288464 277745
rect 342736 277733 342742 277745
rect 342794 277733 342800 277785
rect 355792 277733 355798 277785
rect 355850 277773 355856 277785
rect 443824 277773 443830 277785
rect 355850 277745 443830 277773
rect 355850 277733 355856 277745
rect 443824 277733 443830 277745
rect 443882 277733 443888 277785
rect 289264 277659 289270 277711
rect 289322 277699 289328 277711
rect 350032 277699 350038 277711
rect 289322 277671 350038 277699
rect 289322 277659 289328 277671
rect 350032 277659 350038 277671
rect 350090 277659 350096 277711
rect 358768 277659 358774 277711
rect 358826 277699 358832 277711
rect 384400 277699 384406 277711
rect 358826 277671 384406 277699
rect 358826 277659 358832 277671
rect 384400 277659 384406 277671
rect 384458 277659 384464 277711
rect 384496 277659 384502 277711
rect 384554 277699 384560 277711
rect 454768 277699 454774 277711
rect 384554 277671 454774 277699
rect 384554 277659 384560 277671
rect 454768 277659 454774 277671
rect 454826 277659 454832 277711
rect 294736 277585 294742 277637
rect 294794 277625 294800 277637
rect 396496 277625 396502 277637
rect 294794 277597 396502 277625
rect 294794 277585 294800 277597
rect 396496 277585 396502 277597
rect 396554 277585 396560 277637
rect 289936 277511 289942 277563
rect 289994 277551 290000 277563
rect 357232 277551 357238 277563
rect 289994 277523 357238 277551
rect 289994 277511 290000 277523
rect 357232 277511 357238 277523
rect 357290 277511 357296 277563
rect 368272 277511 368278 277563
rect 368330 277551 368336 277563
rect 375184 277551 375190 277563
rect 368330 277523 375190 277551
rect 368330 277511 368336 277523
rect 375184 277511 375190 277523
rect 375242 277511 375248 277563
rect 375280 277511 375286 277563
rect 375338 277551 375344 277563
rect 383824 277551 383830 277563
rect 375338 277523 383830 277551
rect 375338 277511 375344 277523
rect 383824 277511 383830 277523
rect 383882 277511 383888 277563
rect 383920 277511 383926 277563
rect 383978 277551 383984 277563
rect 384304 277551 384310 277563
rect 383978 277523 384310 277551
rect 383978 277511 383984 277523
rect 384304 277511 384310 277523
rect 384362 277511 384368 277563
rect 384400 277511 384406 277563
rect 384458 277551 384464 277563
rect 465520 277551 465526 277563
rect 384458 277523 465526 277551
rect 384458 277511 384464 277523
rect 465520 277511 465526 277523
rect 465578 277511 465584 277563
rect 295792 277437 295798 277489
rect 295850 277477 295856 277489
rect 403600 277477 403606 277489
rect 295850 277449 403606 277477
rect 295850 277437 295856 277449
rect 403600 277437 403606 277449
rect 403658 277437 403664 277489
rect 42064 277363 42070 277415
rect 42122 277403 42128 277415
rect 43024 277403 43030 277415
rect 42122 277375 43030 277403
rect 42122 277363 42128 277375
rect 43024 277363 43030 277375
rect 43082 277363 43088 277415
rect 296464 277363 296470 277415
rect 296522 277403 296528 277415
rect 410800 277403 410806 277415
rect 296522 277375 410806 277403
rect 296522 277363 296528 277375
rect 410800 277363 410806 277375
rect 410858 277363 410864 277415
rect 240688 277289 240694 277341
rect 240746 277329 240752 277341
rect 331312 277329 331318 277341
rect 240746 277301 331318 277329
rect 240746 277289 240752 277301
rect 331312 277289 331318 277301
rect 331370 277289 331376 277341
rect 351088 277289 351094 277341
rect 351146 277329 351152 277341
rect 380272 277329 380278 277341
rect 351146 277301 380278 277329
rect 351146 277289 351152 277301
rect 380272 277289 380278 277301
rect 380330 277289 380336 277341
rect 380368 277289 380374 277341
rect 380426 277329 380432 277341
rect 384112 277329 384118 277341
rect 380426 277301 384118 277329
rect 380426 277289 380432 277301
rect 384112 277289 384118 277301
rect 384170 277289 384176 277341
rect 384208 277289 384214 277341
rect 384266 277329 384272 277341
rect 479728 277329 479734 277341
rect 384266 277301 479734 277329
rect 384266 277289 384272 277301
rect 479728 277289 479734 277301
rect 479786 277289 479792 277341
rect 297520 277215 297526 277267
rect 297578 277255 297584 277267
rect 417904 277255 417910 277267
rect 297578 277227 417910 277255
rect 297578 277215 297584 277227
rect 417904 277215 417910 277227
rect 417962 277215 417968 277267
rect 317968 277141 317974 277193
rect 318026 277181 318032 277193
rect 439312 277181 439318 277193
rect 318026 277153 439318 277181
rect 318026 277141 318032 277153
rect 439312 277141 439318 277153
rect 439370 277141 439376 277193
rect 298192 277067 298198 277119
rect 298250 277107 298256 277119
rect 425008 277107 425014 277119
rect 298250 277079 425014 277107
rect 298250 277067 298256 277079
rect 425008 277067 425014 277079
rect 425066 277067 425072 277119
rect 254896 276993 254902 277045
rect 254954 277033 254960 277045
rect 332752 277033 332758 277045
rect 254954 277005 332758 277033
rect 254954 276993 254960 277005
rect 332752 276993 332758 277005
rect 332810 276993 332816 277045
rect 360496 276993 360502 277045
rect 360554 277033 360560 277045
rect 384208 277033 384214 277045
rect 360554 277005 384214 277033
rect 360554 276993 360560 277005
rect 384208 276993 384214 277005
rect 384266 276993 384272 277045
rect 384400 276993 384406 277045
rect 384458 277033 384464 277045
rect 391600 277033 391606 277045
rect 384458 277005 391606 277033
rect 384458 276993 384464 277005
rect 391600 276993 391606 277005
rect 391658 276993 391664 277045
rect 297808 276919 297814 276971
rect 297866 276959 297872 276971
rect 338128 276959 338134 276971
rect 297866 276931 338134 276959
rect 297866 276919 297872 276931
rect 338128 276919 338134 276931
rect 338186 276919 338192 276971
rect 365872 276919 365878 276971
rect 365930 276959 365936 276971
rect 365930 276931 384446 276959
rect 365930 276919 365936 276931
rect 269200 276845 269206 276897
rect 269258 276885 269264 276897
rect 334480 276885 334486 276897
rect 269258 276857 334486 276885
rect 269258 276845 269264 276857
rect 334480 276845 334486 276857
rect 334538 276845 334544 276897
rect 357712 276845 357718 276897
rect 357770 276885 357776 276897
rect 384304 276885 384310 276897
rect 357770 276857 384310 276885
rect 357770 276845 357776 276857
rect 384304 276845 384310 276857
rect 384362 276845 384368 276897
rect 384418 276885 384446 276931
rect 384496 276919 384502 276971
rect 384554 276959 384560 276971
rect 508336 276959 508342 276971
rect 384554 276931 508342 276959
rect 384554 276919 384560 276931
rect 508336 276919 508342 276931
rect 508394 276919 508400 276971
rect 398992 276885 398998 276897
rect 384418 276857 398998 276885
rect 398992 276845 398998 276857
rect 399050 276845 399056 276897
rect 262096 276771 262102 276823
rect 262154 276811 262160 276823
rect 333904 276811 333910 276823
rect 262154 276783 333910 276811
rect 262154 276771 262160 276783
rect 333904 276771 333910 276783
rect 333962 276771 333968 276823
rect 362128 276771 362134 276823
rect 362186 276811 362192 276823
rect 403216 276811 403222 276823
rect 362186 276783 403222 276811
rect 362186 276771 362192 276783
rect 403216 276771 403222 276783
rect 403274 276771 403280 276823
rect 247888 276697 247894 276749
rect 247946 276737 247952 276749
rect 332176 276737 332182 276749
rect 247946 276709 332182 276737
rect 247946 276697 247952 276709
rect 332176 276697 332182 276709
rect 332234 276697 332240 276749
rect 349168 276697 349174 276749
rect 349226 276737 349232 276749
rect 349226 276709 372926 276737
rect 349226 276697 349232 276709
rect 239440 276623 239446 276675
rect 239498 276663 239504 276675
rect 252304 276663 252310 276675
rect 239498 276635 252310 276663
rect 239498 276623 239504 276635
rect 252304 276623 252310 276635
rect 252362 276623 252368 276675
rect 290800 276623 290806 276675
rect 290858 276663 290864 276675
rect 364432 276663 364438 276675
rect 290858 276635 364438 276663
rect 290858 276623 290864 276635
rect 364432 276623 364438 276635
rect 364490 276623 364496 276675
rect 212176 276549 212182 276601
rect 212234 276589 212240 276601
rect 327376 276589 327382 276601
rect 212234 276561 327382 276589
rect 212234 276549 212240 276561
rect 327376 276549 327382 276561
rect 327434 276549 327440 276601
rect 372898 276589 372926 276709
rect 375184 276697 375190 276749
rect 375242 276737 375248 276749
rect 379984 276737 379990 276749
rect 375242 276709 379990 276737
rect 375242 276697 375248 276709
rect 379984 276697 379990 276709
rect 380042 276697 380048 276749
rect 380080 276697 380086 276749
rect 380138 276737 380144 276749
rect 381136 276737 381142 276749
rect 380138 276709 381142 276737
rect 380138 276697 380144 276709
rect 381136 276697 381142 276709
rect 381194 276697 381200 276749
rect 381232 276697 381238 276749
rect 381290 276737 381296 276749
rect 381290 276709 384638 276737
rect 381290 276697 381296 276709
rect 372976 276623 372982 276675
rect 373034 276663 373040 276675
rect 384496 276663 384502 276675
rect 373034 276635 384502 276663
rect 373034 276623 373040 276635
rect 384496 276623 384502 276635
rect 384554 276623 384560 276675
rect 384610 276663 384638 276709
rect 386224 276697 386230 276749
rect 386282 276737 386288 276749
rect 400048 276737 400054 276749
rect 386282 276709 400054 276737
rect 386282 276697 386288 276709
rect 400048 276697 400054 276709
rect 400106 276697 400112 276749
rect 384610 276635 387134 276663
rect 386992 276589 386998 276601
rect 372898 276561 386998 276589
rect 386992 276549 386998 276561
rect 387050 276549 387056 276601
rect 387106 276589 387134 276635
rect 387184 276623 387190 276675
rect 387242 276663 387248 276675
rect 615376 276663 615382 276675
rect 387242 276635 615382 276663
rect 387242 276623 387248 276635
rect 615376 276623 615382 276635
rect 615434 276623 615440 276675
rect 640336 276589 640342 276601
rect 387106 276561 640342 276589
rect 640336 276549 640342 276561
rect 640394 276549 640400 276601
rect 194320 276475 194326 276527
rect 194378 276515 194384 276527
rect 325744 276515 325750 276527
rect 194378 276487 325750 276515
rect 194378 276475 194384 276487
rect 325744 276475 325750 276487
rect 325802 276475 325808 276527
rect 374320 276475 374326 276527
rect 374378 276515 374384 276527
rect 639088 276515 639094 276527
rect 374378 276487 639094 276515
rect 374378 276475 374384 276487
rect 639088 276475 639094 276487
rect 639146 276475 639152 276527
rect 42352 276401 42358 276453
rect 42410 276441 42416 276453
rect 53584 276441 53590 276453
rect 42410 276413 53590 276441
rect 42410 276401 42416 276413
rect 53584 276401 53590 276413
rect 53642 276401 53648 276453
rect 231760 276401 231766 276453
rect 231818 276441 231824 276453
rect 334576 276441 334582 276453
rect 231818 276413 334582 276441
rect 231818 276401 231824 276413
rect 334576 276401 334582 276413
rect 334634 276401 334640 276453
rect 365008 276401 365014 276453
rect 365066 276441 365072 276453
rect 369136 276441 369142 276453
rect 365066 276413 369142 276441
rect 365066 276401 365072 276413
rect 369136 276401 369142 276413
rect 369194 276401 369200 276453
rect 371344 276401 371350 276453
rect 371402 276441 371408 276453
rect 374128 276441 374134 276453
rect 371402 276413 374134 276441
rect 371402 276401 371408 276413
rect 374128 276401 374134 276413
rect 374186 276401 374192 276453
rect 374224 276401 374230 276453
rect 374282 276441 374288 276453
rect 375472 276441 375478 276453
rect 374282 276413 375478 276441
rect 374282 276401 374288 276413
rect 375472 276401 375478 276413
rect 375530 276401 375536 276453
rect 375664 276401 375670 276453
rect 375722 276441 375728 276453
rect 384112 276441 384118 276453
rect 375722 276413 384118 276441
rect 375722 276401 375728 276413
rect 384112 276401 384118 276413
rect 384170 276401 384176 276453
rect 384208 276401 384214 276453
rect 384266 276441 384272 276453
rect 384880 276441 384886 276453
rect 384266 276413 384886 276441
rect 384266 276401 384272 276413
rect 384880 276401 384886 276413
rect 384938 276401 384944 276453
rect 385072 276401 385078 276453
rect 385130 276441 385136 276453
rect 561808 276441 561814 276453
rect 385130 276413 561814 276441
rect 385130 276401 385136 276413
rect 561808 276401 561814 276413
rect 561866 276401 561872 276453
rect 232336 276327 232342 276379
rect 232394 276367 232400 276379
rect 341776 276367 341782 276379
rect 232394 276339 341782 276367
rect 232394 276327 232400 276339
rect 341776 276327 341782 276339
rect 341834 276327 341840 276379
rect 372496 276327 372502 276379
rect 372554 276367 372560 276379
rect 374704 276367 374710 276379
rect 372554 276339 374710 276367
rect 372554 276327 372560 276339
rect 374704 276327 374710 276339
rect 374762 276327 374768 276379
rect 375568 276327 375574 276379
rect 375626 276367 375632 276379
rect 391696 276367 391702 276379
rect 375626 276339 391702 276367
rect 375626 276327 375632 276339
rect 391696 276327 391702 276339
rect 391754 276327 391760 276379
rect 395056 276327 395062 276379
rect 395114 276367 395120 276379
rect 568912 276367 568918 276379
rect 395114 276339 568918 276367
rect 395114 276327 395120 276339
rect 568912 276327 568918 276339
rect 568970 276327 568976 276379
rect 244720 276253 244726 276305
rect 244778 276293 244784 276305
rect 441712 276293 441718 276305
rect 244778 276265 441718 276293
rect 244778 276253 244784 276265
rect 441712 276253 441718 276265
rect 441770 276253 441776 276305
rect 245392 276179 245398 276231
rect 245450 276219 245456 276231
rect 448816 276219 448822 276231
rect 245450 276191 448822 276219
rect 245450 276179 245456 276191
rect 448816 276179 448822 276191
rect 448874 276179 448880 276231
rect 233392 276105 233398 276157
rect 233450 276145 233456 276157
rect 348976 276145 348982 276157
rect 233450 276117 348982 276145
rect 233450 276105 233456 276117
rect 348976 276105 348982 276117
rect 349034 276105 349040 276157
rect 367504 276105 367510 276157
rect 367562 276145 367568 276157
rect 375376 276145 375382 276157
rect 367562 276117 375382 276145
rect 367562 276105 367568 276117
rect 375376 276105 375382 276117
rect 375434 276105 375440 276157
rect 376336 276105 376342 276157
rect 376394 276145 376400 276157
rect 383920 276145 383926 276157
rect 376394 276117 383926 276145
rect 376394 276105 376400 276117
rect 383920 276105 383926 276117
rect 383978 276105 383984 276157
rect 384688 276105 384694 276157
rect 384746 276145 384752 276157
rect 576112 276145 576118 276157
rect 384746 276117 576118 276145
rect 384746 276105 384752 276117
rect 576112 276105 576118 276117
rect 576170 276105 576176 276157
rect 246352 276031 246358 276083
rect 246410 276071 246416 276083
rect 455920 276071 455926 276083
rect 246410 276043 455926 276071
rect 246410 276031 246416 276043
rect 455920 276031 455926 276043
rect 455978 276031 455984 276083
rect 234064 275957 234070 276009
rect 234122 275997 234128 276009
rect 356080 275997 356086 276009
rect 234122 275969 356086 275997
rect 234122 275957 234128 275969
rect 356080 275957 356086 275969
rect 356138 275957 356144 276009
rect 368080 275957 368086 276009
rect 368138 275997 368144 276009
rect 375664 275997 375670 276009
rect 368138 275969 375670 275997
rect 368138 275957 368144 275969
rect 375664 275957 375670 275969
rect 375722 275957 375728 276009
rect 375760 275957 375766 276009
rect 375818 275997 375824 276009
rect 379888 275997 379894 276009
rect 375818 275969 379894 275997
rect 375818 275957 375824 275969
rect 379888 275957 379894 275969
rect 379946 275957 379952 276009
rect 379984 275957 379990 276009
rect 380042 275997 380048 276009
rect 383536 275997 383542 276009
rect 380042 275969 383542 275997
rect 380042 275957 380048 275969
rect 383536 275957 383542 275969
rect 383594 275957 383600 276009
rect 384304 275957 384310 276009
rect 384362 275997 384368 276009
rect 583216 275997 583222 276009
rect 384362 275969 583222 275997
rect 384362 275957 384368 275969
rect 583216 275957 583222 275969
rect 583274 275957 583280 276009
rect 247408 275883 247414 275935
rect 247466 275923 247472 275935
rect 463120 275923 463126 275935
rect 247466 275895 463126 275923
rect 247466 275883 247472 275895
rect 463120 275883 463126 275895
rect 463178 275883 463184 275935
rect 204976 275809 204982 275861
rect 205034 275849 205040 275861
rect 317584 275849 317590 275861
rect 205034 275821 317590 275849
rect 205034 275809 205040 275821
rect 317584 275809 317590 275821
rect 317642 275809 317648 275861
rect 317680 275809 317686 275861
rect 317738 275849 317744 275861
rect 324016 275849 324022 275861
rect 317738 275821 324022 275849
rect 317738 275809 317744 275821
rect 324016 275809 324022 275821
rect 324074 275809 324080 275861
rect 324496 275809 324502 275861
rect 324554 275849 324560 275861
rect 374320 275849 374326 275861
rect 324554 275821 374326 275849
rect 324554 275809 324560 275821
rect 374320 275809 374326 275821
rect 374378 275809 374384 275861
rect 374608 275809 374614 275861
rect 374666 275849 374672 275861
rect 377968 275849 377974 275861
rect 374666 275821 377974 275849
rect 374666 275809 374672 275821
rect 377968 275809 377974 275821
rect 378026 275809 378032 275861
rect 378064 275809 378070 275861
rect 378122 275849 378128 275861
rect 384304 275849 384310 275861
rect 378122 275821 384310 275849
rect 378122 275809 378128 275821
rect 384304 275809 384310 275821
rect 384362 275809 384368 275861
rect 384400 275809 384406 275861
rect 384458 275849 384464 275861
rect 590320 275849 590326 275861
rect 384458 275821 590326 275849
rect 384458 275809 384464 275821
rect 590320 275809 590326 275821
rect 590378 275809 590384 275861
rect 248080 275735 248086 275787
rect 248138 275775 248144 275787
rect 470224 275775 470230 275787
rect 248138 275747 470230 275775
rect 248138 275735 248144 275747
rect 470224 275735 470230 275747
rect 470282 275735 470288 275787
rect 235024 275661 235030 275713
rect 235082 275701 235088 275713
rect 363184 275701 363190 275713
rect 235082 275673 363190 275701
rect 235082 275661 235088 275673
rect 363184 275661 363190 275673
rect 363242 275661 363248 275713
rect 364240 275661 364246 275713
rect 364298 275701 364304 275713
rect 372976 275701 372982 275713
rect 364298 275673 372982 275701
rect 364298 275661 364304 275673
rect 372976 275661 372982 275673
rect 373034 275661 373040 275713
rect 374032 275661 374038 275713
rect 374090 275701 374096 275713
rect 384400 275701 384406 275713
rect 374090 275673 384406 275701
rect 374090 275661 374096 275673
rect 384400 275661 384406 275673
rect 384458 275661 384464 275713
rect 384784 275661 384790 275713
rect 384842 275701 384848 275713
rect 385072 275701 385078 275713
rect 384842 275673 385078 275701
rect 384842 275661 384848 275673
rect 385072 275661 385078 275673
rect 385130 275661 385136 275713
rect 385168 275661 385174 275713
rect 385226 275701 385232 275713
rect 604624 275701 604630 275713
rect 385226 275673 604630 275701
rect 385226 275661 385232 275673
rect 604624 275661 604630 275673
rect 604682 275661 604688 275713
rect 235984 275587 235990 275639
rect 236042 275627 236048 275639
rect 370288 275627 370294 275639
rect 236042 275599 370294 275627
rect 236042 275587 236048 275599
rect 370288 275587 370294 275599
rect 370346 275587 370352 275639
rect 377776 275587 377782 275639
rect 377834 275627 377840 275639
rect 390544 275627 390550 275639
rect 377834 275599 390550 275627
rect 377834 275587 377840 275599
rect 390544 275587 390550 275599
rect 390602 275587 390608 275639
rect 398896 275587 398902 275639
rect 398954 275627 398960 275639
rect 618832 275627 618838 275639
rect 398954 275599 618838 275627
rect 398954 275587 398960 275599
rect 618832 275587 618838 275599
rect 618890 275587 618896 275639
rect 226288 275513 226294 275565
rect 226346 275553 226352 275565
rect 291856 275553 291862 275565
rect 226346 275525 291862 275553
rect 226346 275513 226352 275525
rect 291856 275513 291862 275525
rect 291914 275513 291920 275565
rect 317584 275513 317590 275565
rect 317642 275553 317648 275565
rect 326992 275553 326998 275565
rect 317642 275525 326998 275553
rect 317642 275513 317648 275525
rect 326992 275513 326998 275525
rect 327050 275513 327056 275565
rect 327088 275513 327094 275565
rect 327146 275553 327152 275565
rect 557008 275553 557014 275565
rect 327146 275525 557014 275553
rect 327146 275513 327152 275525
rect 557008 275513 557014 275525
rect 557066 275513 557072 275565
rect 227440 275439 227446 275491
rect 227498 275479 227504 275491
rect 298960 275479 298966 275491
rect 227498 275451 298966 275479
rect 227498 275439 227504 275451
rect 298960 275439 298966 275451
rect 299018 275439 299024 275491
rect 315376 275439 315382 275491
rect 315434 275479 315440 275491
rect 564208 275479 564214 275491
rect 315434 275451 564214 275479
rect 315434 275439 315440 275451
rect 564208 275439 564214 275451
rect 564266 275439 564272 275491
rect 200176 275365 200182 275417
rect 200234 275405 200240 275417
rect 267664 275405 267670 275417
rect 200234 275377 267670 275405
rect 200234 275365 200240 275377
rect 267664 275365 267670 275377
rect 267722 275365 267728 275417
rect 267760 275365 267766 275417
rect 267818 275405 267824 275417
rect 270256 275405 270262 275417
rect 267818 275377 270262 275405
rect 267818 275365 267824 275377
rect 270256 275365 270262 275377
rect 270314 275365 270320 275417
rect 315952 275365 315958 275417
rect 316010 275405 316016 275417
rect 571312 275405 571318 275417
rect 316010 275377 571318 275405
rect 316010 275365 316016 275377
rect 571312 275365 571318 275377
rect 571370 275365 571376 275417
rect 236752 275291 236758 275343
rect 236810 275331 236816 275343
rect 377488 275331 377494 275343
rect 236810 275303 377494 275331
rect 236810 275291 236816 275303
rect 377488 275291 377494 275303
rect 377546 275291 377552 275343
rect 377584 275291 377590 275343
rect 377642 275331 377648 275343
rect 385168 275331 385174 275343
rect 377642 275303 385174 275331
rect 377642 275291 377648 275303
rect 385168 275291 385174 275303
rect 385226 275291 385232 275343
rect 385264 275291 385270 275343
rect 385322 275331 385328 275343
rect 394480 275331 394486 275343
rect 385322 275303 394486 275331
rect 385322 275291 385328 275303
rect 394480 275291 394486 275303
rect 394538 275291 394544 275343
rect 398800 275291 398806 275343
rect 398858 275331 398864 275343
rect 636688 275331 636694 275343
rect 398858 275303 636694 275331
rect 398858 275291 398864 275303
rect 636688 275291 636694 275303
rect 636746 275291 636752 275343
rect 196720 275217 196726 275269
rect 196778 275257 196784 275269
rect 257584 275257 257590 275269
rect 196778 275229 257590 275257
rect 196778 275217 196784 275229
rect 257584 275217 257590 275229
rect 257642 275217 257648 275269
rect 317584 275217 317590 275269
rect 317642 275257 317648 275269
rect 578512 275257 578518 275269
rect 317642 275229 578518 275257
rect 317642 275217 317648 275229
rect 578512 275217 578518 275229
rect 578570 275217 578576 275269
rect 228016 275143 228022 275195
rect 228074 275183 228080 275195
rect 257488 275183 257494 275195
rect 228074 275155 257494 275183
rect 228074 275143 228080 275155
rect 257488 275143 257494 275155
rect 257546 275143 257552 275195
rect 257872 275143 257878 275195
rect 257930 275183 257936 275195
rect 306064 275183 306070 275195
rect 257930 275155 306070 275183
rect 257930 275143 257936 275155
rect 306064 275143 306070 275155
rect 306122 275143 306128 275195
rect 314320 275143 314326 275195
rect 314378 275183 314384 275195
rect 317680 275183 317686 275195
rect 314378 275155 317686 275183
rect 314378 275143 314384 275155
rect 317680 275143 317686 275155
rect 317738 275143 317744 275195
rect 318640 275143 318646 275195
rect 318698 275183 318704 275195
rect 318698 275155 338366 275183
rect 318698 275143 318704 275155
rect 193072 275069 193078 275121
rect 193130 275109 193136 275121
rect 257584 275109 257590 275121
rect 193130 275081 257590 275109
rect 193130 275069 193136 275081
rect 257584 275069 257590 275081
rect 257642 275069 257648 275121
rect 257776 275069 257782 275121
rect 257834 275109 257840 275121
rect 267664 275109 267670 275121
rect 257834 275081 267670 275109
rect 257834 275069 257840 275081
rect 267664 275069 267670 275081
rect 267722 275069 267728 275121
rect 267760 275069 267766 275121
rect 267818 275109 267824 275121
rect 272464 275109 272470 275121
rect 267818 275081 272470 275109
rect 267818 275069 267824 275081
rect 272464 275069 272470 275081
rect 272522 275069 272528 275121
rect 284944 275069 284950 275121
rect 285002 275109 285008 275121
rect 314416 275109 314422 275121
rect 285002 275081 314422 275109
rect 285002 275069 285008 275081
rect 314416 275069 314422 275081
rect 314474 275069 314480 275121
rect 319792 275069 319798 275121
rect 319850 275109 319856 275121
rect 338338 275109 338366 275155
rect 338416 275143 338422 275195
rect 338474 275183 338480 275195
rect 585616 275183 585622 275195
rect 338474 275155 585622 275183
rect 338474 275143 338480 275155
rect 585616 275143 585622 275155
rect 585674 275143 585680 275195
rect 592720 275109 592726 275121
rect 319850 275081 338270 275109
rect 338338 275081 592726 275109
rect 319850 275069 319856 275081
rect 229072 274995 229078 275047
rect 229130 275035 229136 275047
rect 313264 275035 313270 275047
rect 229130 275007 313270 275035
rect 229130 274995 229136 275007
rect 313264 274995 313270 275007
rect 313322 274995 313328 275047
rect 318160 274995 318166 275047
rect 318218 275035 318224 275047
rect 330160 275035 330166 275047
rect 318218 275007 330166 275035
rect 318218 274995 318224 275007
rect 330160 274995 330166 275007
rect 330218 274995 330224 275047
rect 338242 275035 338270 275081
rect 592720 275069 592726 275081
rect 592778 275069 592784 275121
rect 599824 275035 599830 275047
rect 338242 275007 599830 275035
rect 599824 274995 599830 275007
rect 599882 274995 599888 275047
rect 243760 274921 243766 274973
rect 243818 274961 243824 274973
rect 434512 274961 434518 274973
rect 243818 274933 434518 274961
rect 243818 274921 243824 274933
rect 434512 274921 434518 274933
rect 434570 274921 434576 274973
rect 663856 274921 663862 274973
rect 663914 274961 663920 274973
rect 674704 274961 674710 274973
rect 663914 274933 674710 274961
rect 663914 274921 663920 274933
rect 674704 274921 674710 274933
rect 674762 274921 674768 274973
rect 242992 274847 242998 274899
rect 243050 274887 243056 274899
rect 427408 274887 427414 274899
rect 243050 274859 427414 274887
rect 243050 274847 243056 274859
rect 427408 274847 427414 274859
rect 427466 274847 427472 274899
rect 233488 274773 233494 274825
rect 233546 274813 233552 274825
rect 318160 274813 318166 274825
rect 233546 274785 318166 274813
rect 233546 274773 233552 274785
rect 318160 274773 318166 274785
rect 318218 274773 318224 274825
rect 318256 274773 318262 274825
rect 318314 274813 318320 274825
rect 335632 274813 335638 274825
rect 318314 274785 335638 274813
rect 318314 274773 318320 274785
rect 335632 274773 335638 274785
rect 335690 274773 335696 274825
rect 362704 274773 362710 274825
rect 362762 274813 362768 274825
rect 375760 274813 375766 274825
rect 362762 274785 375766 274813
rect 362762 274773 362768 274785
rect 375760 274773 375766 274785
rect 375818 274773 375824 274825
rect 377872 274773 377878 274825
rect 377930 274813 377936 274825
rect 554704 274813 554710 274825
rect 377930 274785 554710 274813
rect 377930 274773 377936 274785
rect 554704 274773 554710 274785
rect 554762 274773 554768 274825
rect 242224 274699 242230 274751
rect 242282 274739 242288 274751
rect 420208 274739 420214 274751
rect 242282 274711 420214 274739
rect 242282 274699 242288 274711
rect 420208 274699 420214 274711
rect 420266 274699 420272 274751
rect 241072 274625 241078 274677
rect 241130 274665 241136 274677
rect 413200 274665 413206 274677
rect 241130 274637 413206 274665
rect 241130 274625 241136 274637
rect 413200 274625 413206 274637
rect 413258 274625 413264 274677
rect 429232 274625 429238 274677
rect 429290 274665 429296 274677
rect 449104 274665 449110 274677
rect 429290 274637 449110 274665
rect 429290 274625 429296 274637
rect 449104 274625 449110 274637
rect 449162 274625 449168 274677
rect 153808 274551 153814 274603
rect 153866 274591 153872 274603
rect 161200 274591 161206 274603
rect 153866 274563 161206 274591
rect 153866 274551 153872 274563
rect 161200 274551 161206 274563
rect 161258 274551 161264 274603
rect 240496 274551 240502 274603
rect 240554 274591 240560 274603
rect 406000 274591 406006 274603
rect 240554 274563 406006 274591
rect 240554 274551 240560 274563
rect 406000 274551 406006 274563
rect 406058 274551 406064 274603
rect 619120 274551 619126 274603
rect 619178 274591 619184 274603
rect 627280 274591 627286 274603
rect 619178 274563 627286 274591
rect 619178 274551 619184 274563
rect 627280 274551 627286 274563
rect 627338 274551 627344 274603
rect 239344 274477 239350 274529
rect 239402 274517 239408 274529
rect 398608 274517 398614 274529
rect 239402 274489 398614 274517
rect 239402 274477 239408 274489
rect 398608 274477 398614 274489
rect 398666 274477 398672 274529
rect 238480 274403 238486 274455
rect 238538 274443 238544 274455
rect 375568 274443 375574 274455
rect 238538 274415 375574 274443
rect 238538 274403 238544 274415
rect 375568 274403 375574 274415
rect 375626 274403 375632 274455
rect 375760 274403 375766 274455
rect 375818 274443 375824 274455
rect 377584 274443 377590 274455
rect 375818 274415 377590 274443
rect 375818 274403 375824 274415
rect 377584 274403 377590 274415
rect 377642 274403 377648 274455
rect 379120 274443 379126 274455
rect 377698 274415 379126 274443
rect 237808 274329 237814 274381
rect 237866 274369 237872 274381
rect 376336 274369 376342 274381
rect 237866 274341 376342 274369
rect 237866 274329 237872 274341
rect 376336 274329 376342 274341
rect 376394 274329 376400 274381
rect 377296 274329 377302 274381
rect 377354 274369 377360 274381
rect 377698 274369 377726 274415
rect 379120 274403 379126 274415
rect 379178 274403 379184 274455
rect 379216 274403 379222 274455
rect 379274 274443 379280 274455
rect 385072 274443 385078 274455
rect 379274 274415 385078 274443
rect 379274 274403 379280 274415
rect 385072 274403 385078 274415
rect 385130 274403 385136 274455
rect 593296 274403 593302 274455
rect 593354 274443 593360 274455
rect 613360 274443 613366 274455
rect 593354 274415 613366 274443
rect 593354 274403 593360 274415
rect 613360 274403 613366 274415
rect 613418 274403 613424 274455
rect 377354 274341 377726 274369
rect 377354 274329 377360 274341
rect 378544 274329 378550 274381
rect 378602 274369 378608 274381
rect 383728 274369 383734 274381
rect 378602 274341 383734 274369
rect 378602 274329 378608 274341
rect 383728 274329 383734 274341
rect 383786 274329 383792 274381
rect 383824 274329 383830 274381
rect 383882 274369 383888 274381
rect 384400 274369 384406 274381
rect 383882 274341 384406 274369
rect 383882 274329 383888 274341
rect 384400 274329 384406 274341
rect 384458 274329 384464 274381
rect 384496 274329 384502 274381
rect 384554 274369 384560 274381
rect 394384 274369 394390 274381
rect 384554 274341 394390 274369
rect 384554 274329 384560 274341
rect 394384 274329 394390 274341
rect 394442 274329 394448 274381
rect 394480 274329 394486 274381
rect 394538 274369 394544 274381
rect 398800 274369 398806 274381
rect 394538 274341 398806 274369
rect 394538 274329 394544 274341
rect 398800 274329 398806 274341
rect 398858 274329 398864 274381
rect 230224 274255 230230 274307
rect 230282 274295 230288 274307
rect 323632 274295 323638 274307
rect 230282 274267 323638 274295
rect 230282 274255 230288 274267
rect 323632 274255 323638 274267
rect 323690 274255 323696 274307
rect 324016 274255 324022 274307
rect 324074 274295 324080 274307
rect 327088 274295 327094 274307
rect 324074 274267 327094 274295
rect 324074 274255 324080 274267
rect 327088 274255 327094 274267
rect 327146 274255 327152 274307
rect 338416 274295 338422 274307
rect 327586 274267 338422 274295
rect 230608 274181 230614 274233
rect 230666 274221 230672 274233
rect 327472 274221 327478 274233
rect 230666 274193 327478 274221
rect 230666 274181 230672 274193
rect 327472 274181 327478 274193
rect 327530 274181 327536 274233
rect 207376 274107 207382 274159
rect 207434 274147 207440 274159
rect 271312 274147 271318 274159
rect 207434 274119 271318 274147
rect 207434 274107 207440 274119
rect 271312 274107 271318 274119
rect 271370 274107 271376 274159
rect 276400 274107 276406 274159
rect 276458 274147 276464 274159
rect 318256 274147 318262 274159
rect 276458 274119 318262 274147
rect 276458 274107 276464 274119
rect 318256 274107 318262 274119
rect 318314 274107 318320 274159
rect 318448 274107 318454 274159
rect 318506 274147 318512 274159
rect 327586 274147 327614 274267
rect 338416 274255 338422 274267
rect 338474 274255 338480 274307
rect 368464 274255 368470 274307
rect 368522 274295 368528 274307
rect 368848 274295 368854 274307
rect 368522 274267 368854 274295
rect 368522 274255 368528 274267
rect 368848 274255 368854 274267
rect 368906 274255 368912 274307
rect 369616 274255 369622 274307
rect 369674 274295 369680 274307
rect 377872 274295 377878 274307
rect 369674 274267 377878 274295
rect 369674 274255 369680 274267
rect 377872 274255 377878 274267
rect 377930 274255 377936 274307
rect 377968 274255 377974 274307
rect 378026 274295 378032 274307
rect 383920 274295 383926 274307
rect 378026 274267 383926 274295
rect 378026 274255 378032 274267
rect 383920 274255 383926 274267
rect 383978 274255 383984 274307
rect 472624 274295 472630 274307
rect 384418 274267 472630 274295
rect 359728 274181 359734 274233
rect 359786 274221 359792 274233
rect 384418 274221 384446 274267
rect 472624 274255 472630 274267
rect 472682 274255 472688 274307
rect 359786 274193 384446 274221
rect 359786 274181 359792 274193
rect 384496 274181 384502 274233
rect 384554 274221 384560 274233
rect 458320 274221 458326 274233
rect 384554 274193 458326 274221
rect 384554 274181 384560 274193
rect 458320 274181 458326 274193
rect 458378 274181 458384 274233
rect 469552 274181 469558 274233
rect 469610 274221 469616 274233
rect 477616 274221 477622 274233
rect 469610 274193 477622 274221
rect 469610 274181 469616 274193
rect 477616 274181 477622 274193
rect 477674 274181 477680 274233
rect 552976 274181 552982 274233
rect 553034 274221 553040 274233
rect 573040 274221 573046 274233
rect 553034 274193 573046 274221
rect 553034 274181 553040 274193
rect 573040 274181 573046 274193
rect 573098 274181 573104 274233
rect 318506 274119 327614 274147
rect 318506 274107 318512 274119
rect 355696 274107 355702 274159
rect 355754 274147 355760 274159
rect 440464 274147 440470 274159
rect 355754 274119 440470 274147
rect 355754 274107 355760 274119
rect 440464 274107 440470 274119
rect 440522 274107 440528 274159
rect 214576 274033 214582 274085
rect 214634 274073 214640 274085
rect 252208 274073 252214 274085
rect 214634 274045 252214 274073
rect 214634 274033 214640 274045
rect 252208 274033 252214 274045
rect 252266 274033 252272 274085
rect 252304 274033 252310 274085
rect 252362 274073 252368 274085
rect 275248 274073 275254 274085
rect 252362 274045 275254 274073
rect 252362 274033 252368 274045
rect 275248 274033 275254 274045
rect 275306 274033 275312 274085
rect 287056 274033 287062 274085
rect 287114 274073 287120 274085
rect 336688 274073 336694 274085
rect 287114 274045 336694 274073
rect 287114 274033 287120 274045
rect 336688 274033 336694 274045
rect 336746 274033 336752 274085
rect 353488 274033 353494 274085
rect 353546 274073 353552 274085
rect 422608 274073 422614 274085
rect 353546 274045 422614 274073
rect 353546 274033 353552 274045
rect 422608 274033 422614 274045
rect 422666 274033 422672 274085
rect 661072 274033 661078 274085
rect 661130 274073 661136 274085
rect 674704 274073 674710 274085
rect 661130 274045 674710 274073
rect 661130 274033 661136 274045
rect 674704 274033 674710 274045
rect 674762 274033 674768 274085
rect 225424 273959 225430 274011
rect 225482 273999 225488 274011
rect 284656 273999 284662 274011
rect 225482 273971 284662 273999
rect 225482 273959 225488 273971
rect 284656 273959 284662 273971
rect 284714 273959 284720 274011
rect 317008 273959 317014 274011
rect 317066 273999 317072 274011
rect 335440 273999 335446 274011
rect 317066 273971 335446 273999
rect 317066 273959 317072 273971
rect 335440 273959 335446 273971
rect 335498 273959 335504 274011
rect 358096 273959 358102 274011
rect 358154 273999 358160 274011
rect 384496 273999 384502 274011
rect 358154 273971 384502 273999
rect 358154 273959 358160 273971
rect 384496 273959 384502 273971
rect 384554 273959 384560 274011
rect 384592 273959 384598 274011
rect 384650 273999 384656 274011
rect 392848 273999 392854 274011
rect 384650 273971 392854 273999
rect 384650 273959 384656 273971
rect 392848 273959 392854 273971
rect 392906 273959 392912 274011
rect 225232 273885 225238 273937
rect 225290 273925 225296 273937
rect 281104 273925 281110 273937
rect 225290 273897 281110 273925
rect 225290 273885 225296 273897
rect 281104 273885 281110 273897
rect 281162 273885 281168 273937
rect 301264 273885 301270 273937
rect 301322 273925 301328 273937
rect 338704 273925 338710 273937
rect 301322 273897 338710 273925
rect 301322 273885 301328 273897
rect 338704 273885 338710 273897
rect 338762 273885 338768 273937
rect 370960 273885 370966 273937
rect 371018 273925 371024 273937
rect 396112 273925 396118 273937
rect 371018 273897 396118 273925
rect 371018 273885 371024 273897
rect 396112 273885 396118 273897
rect 396170 273885 396176 273937
rect 224080 273811 224086 273863
rect 224138 273851 224144 273863
rect 274000 273851 274006 273863
rect 224138 273823 274006 273851
rect 224138 273811 224144 273823
rect 274000 273811 274006 273823
rect 274058 273811 274064 273863
rect 274096 273811 274102 273863
rect 274154 273851 274160 273863
rect 274154 273823 286142 273851
rect 274154 273811 274160 273823
rect 223024 273737 223030 273789
rect 223082 273777 223088 273789
rect 223082 273749 252062 273777
rect 223082 273737 223088 273749
rect 158800 273663 158806 273715
rect 158858 273703 158864 273715
rect 178288 273703 178294 273715
rect 158858 273675 178294 273703
rect 158858 273663 158864 273675
rect 178288 273663 178294 273675
rect 178346 273663 178352 273715
rect 252034 273703 252062 273749
rect 252208 273737 252214 273789
rect 252266 273777 252272 273789
rect 267760 273777 267766 273789
rect 252266 273749 267766 273777
rect 252266 273737 252272 273749
rect 267760 273737 267766 273749
rect 267818 273737 267824 273789
rect 269392 273737 269398 273789
rect 269450 273777 269456 273789
rect 286000 273777 286006 273789
rect 269450 273749 286006 273777
rect 269450 273737 269456 273749
rect 286000 273737 286006 273749
rect 286058 273737 286064 273789
rect 286114 273777 286142 273823
rect 286672 273811 286678 273863
rect 286730 273851 286736 273863
rect 328720 273851 328726 273863
rect 286730 273823 328726 273851
rect 286730 273811 286736 273823
rect 328720 273811 328726 273823
rect 328778 273811 328784 273863
rect 343120 273811 343126 273863
rect 343178 273851 343184 273863
rect 359632 273851 359638 273863
rect 343178 273823 359638 273851
rect 343178 273811 343184 273823
rect 359632 273811 359638 273823
rect 359690 273811 359696 273863
rect 361936 273811 361942 273863
rect 361994 273851 362000 273863
rect 400336 273851 400342 273863
rect 361994 273823 400342 273851
rect 361994 273811 362000 273823
rect 400336 273811 400342 273823
rect 400394 273811 400400 273863
rect 370384 273777 370390 273789
rect 286114 273749 370390 273777
rect 370384 273737 370390 273749
rect 370442 273737 370448 273789
rect 373360 273737 373366 273789
rect 373418 273777 373424 273789
rect 378064 273777 378070 273789
rect 373418 273749 378070 273777
rect 373418 273737 373424 273749
rect 378064 273737 378070 273749
rect 378122 273737 378128 273789
rect 378160 273737 378166 273789
rect 378218 273777 378224 273789
rect 383632 273777 383638 273789
rect 378218 273749 383638 273777
rect 378218 273737 378224 273749
rect 383632 273737 383638 273749
rect 383690 273737 383696 273789
rect 383728 273737 383734 273789
rect 383786 273777 383792 273789
rect 398896 273777 398902 273789
rect 383786 273749 398902 273777
rect 383786 273737 383792 273749
rect 398896 273737 398902 273749
rect 398954 273737 398960 273789
rect 263344 273703 263350 273715
rect 252034 273675 263350 273703
rect 263344 273663 263350 273675
rect 263402 273663 263408 273715
rect 267184 273663 267190 273715
rect 267242 273703 267248 273715
rect 372400 273703 372406 273715
rect 267242 273675 372406 273703
rect 267242 273663 267248 273675
rect 372400 273663 372406 273675
rect 372458 273663 372464 273715
rect 372496 273663 372502 273715
rect 372554 273703 372560 273715
rect 377680 273703 377686 273715
rect 372554 273675 377686 273703
rect 372554 273663 372560 273675
rect 377680 273663 377686 273675
rect 377738 273663 377744 273715
rect 378832 273703 378838 273715
rect 378562 273675 378838 273703
rect 143152 273589 143158 273641
rect 143210 273629 143216 273641
rect 160720 273629 160726 273641
rect 143210 273601 160726 273629
rect 143210 273589 143216 273601
rect 160720 273589 160726 273601
rect 160778 273589 160784 273641
rect 267856 273589 267862 273641
rect 267914 273629 267920 273641
rect 270736 273629 270742 273641
rect 267914 273601 270742 273629
rect 267914 273589 267920 273601
rect 270736 273589 270742 273601
rect 270794 273589 270800 273641
rect 270832 273589 270838 273641
rect 270890 273629 270896 273641
rect 274096 273629 274102 273641
rect 270890 273601 274102 273629
rect 270890 273589 270896 273601
rect 274096 273589 274102 273601
rect 274154 273589 274160 273641
rect 285442 273601 285950 273629
rect 102640 273515 102646 273567
rect 102698 273555 102704 273567
rect 211600 273555 211606 273567
rect 102698 273527 211606 273555
rect 102698 273515 102704 273527
rect 211600 273515 211606 273527
rect 211658 273515 211664 273567
rect 228784 273515 228790 273567
rect 228842 273555 228848 273567
rect 274192 273555 274198 273567
rect 228842 273527 274198 273555
rect 228842 273515 228848 273527
rect 274192 273515 274198 273527
rect 274250 273515 274256 273567
rect 275152 273515 275158 273567
rect 275210 273555 275216 273567
rect 279664 273555 279670 273567
rect 275210 273527 279670 273555
rect 275210 273515 275216 273527
rect 279664 273515 279670 273527
rect 279722 273515 279728 273567
rect 67024 273441 67030 273493
rect 67082 273481 67088 273493
rect 209680 273481 209686 273493
rect 67082 273453 209686 273481
rect 67082 273441 67088 273453
rect 209680 273441 209686 273453
rect 209738 273441 209744 273493
rect 209776 273441 209782 273493
rect 209834 273481 209840 273493
rect 216112 273481 216118 273493
rect 209834 273453 216118 273481
rect 209834 273441 209840 273453
rect 216112 273441 216118 273453
rect 216170 273441 216176 273493
rect 218224 273441 218230 273493
rect 218282 273481 218288 273493
rect 223984 273481 223990 273493
rect 218282 273453 223990 273481
rect 218282 273441 218288 273453
rect 223984 273441 223990 273453
rect 224042 273441 224048 273493
rect 224560 273441 224566 273493
rect 224618 273481 224624 273493
rect 277552 273481 277558 273493
rect 224618 273453 277558 273481
rect 224618 273441 224624 273453
rect 277552 273441 277558 273453
rect 277610 273441 277616 273493
rect 278800 273441 278806 273493
rect 278858 273481 278864 273493
rect 280048 273481 280054 273493
rect 278858 273453 280054 273481
rect 278858 273441 278864 273453
rect 280048 273441 280054 273453
rect 280106 273441 280112 273493
rect 280720 273441 280726 273493
rect 280778 273481 280784 273493
rect 282352 273481 282358 273493
rect 280778 273453 282358 273481
rect 280778 273441 280784 273453
rect 282352 273441 282358 273453
rect 282410 273441 282416 273493
rect 284464 273441 284470 273493
rect 284522 273481 284528 273493
rect 285442 273481 285470 273601
rect 285922 273555 285950 273601
rect 286000 273589 286006 273641
rect 286058 273629 286064 273641
rect 378562 273629 378590 273675
rect 378832 273663 378838 273675
rect 378890 273663 378896 273715
rect 378928 273663 378934 273715
rect 378986 273703 378992 273715
rect 379696 273703 379702 273715
rect 378986 273675 379702 273703
rect 378986 273663 378992 273675
rect 379696 273663 379702 273675
rect 379754 273663 379760 273715
rect 380080 273663 380086 273715
rect 380138 273703 380144 273715
rect 394480 273703 394486 273715
rect 380138 273675 394486 273703
rect 380138 273663 380144 273675
rect 394480 273663 394486 273675
rect 394538 273663 394544 273715
rect 286058 273601 378590 273629
rect 286058 273589 286064 273601
rect 378640 273589 378646 273641
rect 378698 273629 378704 273641
rect 379024 273629 379030 273641
rect 378698 273601 379030 273629
rect 378698 273589 378704 273601
rect 379024 273589 379030 273601
rect 379082 273589 379088 273641
rect 379120 273589 379126 273641
rect 379178 273629 379184 273641
rect 387184 273629 387190 273641
rect 379178 273601 387190 273629
rect 379178 273589 379184 273601
rect 387184 273589 387190 273601
rect 387242 273589 387248 273641
rect 388624 273589 388630 273641
rect 388682 273629 388688 273641
rect 391216 273629 391222 273641
rect 388682 273601 391222 273629
rect 388682 273589 388688 273601
rect 391216 273589 391222 273601
rect 391274 273589 391280 273641
rect 310864 273555 310870 273567
rect 285922 273527 310870 273555
rect 310864 273515 310870 273527
rect 310922 273515 310928 273567
rect 319120 273515 319126 273567
rect 319178 273555 319184 273567
rect 323728 273555 323734 273567
rect 319178 273527 323734 273555
rect 319178 273515 319184 273527
rect 323728 273515 323734 273527
rect 323786 273515 323792 273567
rect 323824 273515 323830 273567
rect 323882 273555 323888 273567
rect 553456 273555 553462 273567
rect 323882 273527 553462 273555
rect 323882 273515 323888 273527
rect 553456 273515 553462 273527
rect 553514 273515 553520 273567
rect 284522 273453 285470 273481
rect 284522 273441 284528 273453
rect 285520 273441 285526 273493
rect 285578 273481 285584 273493
rect 321520 273481 321526 273493
rect 285578 273453 321526 273481
rect 285578 273441 285584 273453
rect 321520 273441 321526 273453
rect 321578 273441 321584 273493
rect 321616 273441 321622 273493
rect 321674 273481 321680 273493
rect 334096 273481 334102 273493
rect 321674 273453 334102 273481
rect 321674 273441 321680 273453
rect 334096 273441 334102 273453
rect 334154 273441 334160 273493
rect 336976 273441 336982 273493
rect 337034 273481 337040 273493
rect 343024 273481 343030 273493
rect 337034 273453 343030 273481
rect 337034 273441 337040 273453
rect 343024 273441 343030 273453
rect 343082 273441 343088 273493
rect 347440 273441 347446 273493
rect 347498 273481 347504 273493
rect 349840 273481 349846 273493
rect 347498 273453 349846 273481
rect 347498 273441 347504 273453
rect 349840 273441 349846 273453
rect 349898 273441 349904 273493
rect 351184 273441 351190 273493
rect 351242 273481 351248 273493
rect 362032 273481 362038 273493
rect 351242 273453 362038 273481
rect 351242 273441 351248 273453
rect 362032 273441 362038 273453
rect 362090 273441 362096 273493
rect 368656 273441 368662 273493
rect 368714 273481 368720 273493
rect 369136 273481 369142 273493
rect 368714 273453 369142 273481
rect 368714 273441 368720 273453
rect 369136 273441 369142 273453
rect 369194 273441 369200 273493
rect 370000 273441 370006 273493
rect 370058 273481 370064 273493
rect 378640 273481 378646 273493
rect 370058 273453 378646 273481
rect 370058 273441 370064 273453
rect 378640 273441 378646 273453
rect 378698 273441 378704 273493
rect 379120 273441 379126 273493
rect 379178 273481 379184 273493
rect 379178 273453 389150 273481
rect 379178 273441 379184 273453
rect 161008 273367 161014 273419
rect 161066 273407 161072 273419
rect 377968 273407 377974 273419
rect 161066 273379 377974 273407
rect 161066 273367 161072 273379
rect 377968 273367 377974 273379
rect 378026 273367 378032 273419
rect 378352 273367 378358 273419
rect 378410 273407 378416 273419
rect 389008 273407 389014 273419
rect 378410 273379 389014 273407
rect 378410 273367 378416 273379
rect 389008 273367 389014 273379
rect 389066 273367 389072 273419
rect 389122 273407 389150 273453
rect 391216 273441 391222 273493
rect 391274 273481 391280 273493
rect 622480 273481 622486 273493
rect 391274 273453 622486 273481
rect 391274 273441 391280 273453
rect 622480 273441 622486 273453
rect 622538 273441 622544 273493
rect 393616 273407 393622 273419
rect 389122 273379 393622 273407
rect 393616 273367 393622 273379
rect 393674 273367 393680 273419
rect 393712 273367 393718 273419
rect 393770 273407 393776 273419
rect 402544 273407 402550 273419
rect 393770 273379 402550 273407
rect 393770 273367 393776 273379
rect 402544 273367 402550 273379
rect 402602 273367 402608 273419
rect 403216 273367 403222 273419
rect 403274 273407 403280 273419
rect 494032 273407 494038 273419
rect 403274 273379 494038 273407
rect 403274 273367 403280 273379
rect 494032 273367 494038 273379
rect 494090 273367 494096 273419
rect 144400 273293 144406 273345
rect 144458 273333 144464 273345
rect 146800 273333 146806 273345
rect 144458 273305 146806 273333
rect 144458 273293 144464 273305
rect 146800 273293 146806 273305
rect 146858 273293 146864 273345
rect 157456 273293 157462 273345
rect 157514 273333 157520 273345
rect 404080 273333 404086 273345
rect 157514 273305 404086 273333
rect 157514 273293 157520 273305
rect 404080 273293 404086 273305
rect 404138 273293 404144 273345
rect 664048 273293 664054 273345
rect 664106 273333 664112 273345
rect 674704 273333 674710 273345
rect 664106 273305 674710 273333
rect 664106 273293 664112 273305
rect 674704 273293 674710 273305
rect 674762 273293 674768 273345
rect 65872 273219 65878 273271
rect 65930 273259 65936 273271
rect 212368 273259 212374 273271
rect 65930 273231 212374 273259
rect 65930 273219 65936 273231
rect 212368 273219 212374 273231
rect 212426 273219 212432 273271
rect 213328 273219 213334 273271
rect 213386 273259 213392 273271
rect 216688 273259 216694 273271
rect 213386 273231 216694 273259
rect 213386 273219 213392 273231
rect 216688 273219 216694 273231
rect 216746 273219 216752 273271
rect 217552 273219 217558 273271
rect 217610 273259 217616 273271
rect 220432 273259 220438 273271
rect 217610 273231 220438 273259
rect 217610 273219 217616 273231
rect 220432 273219 220438 273231
rect 220490 273219 220496 273271
rect 229744 273219 229750 273271
rect 229802 273259 229808 273271
rect 320368 273259 320374 273271
rect 229802 273231 320374 273259
rect 229802 273219 229808 273231
rect 320368 273219 320374 273231
rect 320426 273219 320432 273271
rect 320464 273219 320470 273271
rect 320522 273259 320528 273271
rect 323632 273259 323638 273271
rect 320522 273231 323638 273259
rect 320522 273219 320528 273231
rect 323632 273219 323638 273231
rect 323690 273219 323696 273271
rect 323728 273219 323734 273271
rect 323786 273259 323792 273271
rect 340528 273259 340534 273271
rect 323786 273231 340534 273259
rect 323786 273219 323792 273231
rect 340528 273219 340534 273231
rect 340586 273219 340592 273271
rect 340624 273219 340630 273271
rect 340682 273259 340688 273271
rect 343504 273259 343510 273271
rect 340682 273231 343510 273259
rect 340682 273219 340688 273231
rect 343504 273219 343510 273231
rect 343562 273219 343568 273271
rect 344656 273219 344662 273271
rect 344714 273259 344720 273271
rect 347728 273259 347734 273271
rect 344714 273231 347734 273259
rect 344714 273219 344720 273231
rect 347728 273219 347734 273231
rect 347786 273219 347792 273271
rect 347920 273219 347926 273271
rect 347978 273259 347984 273271
rect 349744 273259 349750 273271
rect 347978 273231 349750 273259
rect 347978 273219 347984 273231
rect 349744 273219 349750 273231
rect 349802 273219 349808 273271
rect 349840 273219 349846 273271
rect 349898 273259 349904 273271
rect 372688 273259 372694 273271
rect 349898 273231 372694 273259
rect 349898 273219 349904 273231
rect 372688 273219 372694 273231
rect 372746 273219 372752 273271
rect 374416 273219 374422 273271
rect 374474 273259 374480 273271
rect 376240 273259 376246 273271
rect 374474 273231 376246 273259
rect 374474 273219 374480 273231
rect 376240 273219 376246 273231
rect 376298 273219 376304 273271
rect 376336 273219 376342 273271
rect 376394 273259 376400 273271
rect 379312 273259 379318 273271
rect 376394 273231 379318 273259
rect 376394 273219 376400 273231
rect 379312 273219 379318 273231
rect 379370 273219 379376 273271
rect 379408 273219 379414 273271
rect 379466 273259 379472 273271
rect 388624 273259 388630 273271
rect 379466 273231 388630 273259
rect 379466 273219 379472 273231
rect 388624 273219 388630 273231
rect 388682 273219 388688 273271
rect 388720 273219 388726 273271
rect 388778 273259 388784 273271
rect 395344 273259 395350 273271
rect 388778 273231 395350 273259
rect 388778 273219 388784 273231
rect 395344 273219 395350 273231
rect 395402 273219 395408 273271
rect 396016 273219 396022 273271
rect 396074 273259 396080 273271
rect 396074 273231 398846 273259
rect 396074 273219 396080 273231
rect 161296 273145 161302 273197
rect 161354 273185 161360 273197
rect 161354 273157 164222 273185
rect 161354 273145 161360 273157
rect 147952 273071 147958 273123
rect 148010 273111 148016 273123
rect 149680 273111 149686 273123
rect 148010 273083 149686 273111
rect 148010 273071 148016 273083
rect 149680 273071 149686 273083
rect 149738 273071 149744 273123
rect 152656 273071 152662 273123
rect 152714 273111 152720 273123
rect 155344 273111 155350 273123
rect 152714 273083 155350 273111
rect 152714 273071 152720 273083
rect 155344 273071 155350 273083
rect 155402 273071 155408 273123
rect 156208 273071 156214 273123
rect 156266 273111 156272 273123
rect 158320 273111 158326 273123
rect 156266 273083 158326 273111
rect 156266 273071 156272 273083
rect 158320 273071 158326 273083
rect 158378 273071 158384 273123
rect 162160 273071 162166 273123
rect 162218 273111 162224 273123
rect 164080 273111 164086 273123
rect 162218 273083 164086 273111
rect 162218 273071 162224 273083
rect 164080 273071 164086 273083
rect 164138 273071 164144 273123
rect 164194 273111 164222 273157
rect 164272 273145 164278 273197
rect 164330 273185 164336 273197
rect 378352 273185 378358 273197
rect 164330 273157 378358 273185
rect 164330 273145 164336 273157
rect 378352 273145 378358 273157
rect 378410 273145 378416 273197
rect 378736 273145 378742 273197
rect 378794 273185 378800 273197
rect 397072 273185 397078 273197
rect 378794 273157 397078 273185
rect 378794 273145 378800 273157
rect 397072 273145 397078 273157
rect 397130 273145 397136 273197
rect 397360 273145 397366 273197
rect 397418 273185 397424 273197
rect 398704 273185 398710 273197
rect 397418 273157 398710 273185
rect 397418 273145 397424 273157
rect 398704 273145 398710 273157
rect 398762 273145 398768 273197
rect 398818 273185 398846 273231
rect 398896 273219 398902 273271
rect 398954 273259 398960 273271
rect 629680 273259 629686 273271
rect 398954 273231 629686 273259
rect 398954 273219 398960 273231
rect 629680 273219 629686 273231
rect 629738 273219 629744 273271
rect 399856 273185 399862 273197
rect 398818 273157 399862 273185
rect 399856 273145 399862 273157
rect 399914 273145 399920 273197
rect 400336 273145 400342 273197
rect 400394 273185 400400 273197
rect 490480 273185 490486 273197
rect 400394 273157 490486 273185
rect 400394 273145 400400 273157
rect 490480 273145 490486 273157
rect 490538 273145 490544 273197
rect 362992 273111 362998 273123
rect 164194 273083 362998 273111
rect 362992 273071 362998 273083
rect 363050 273071 363056 273123
rect 363376 273071 363382 273123
rect 363434 273111 363440 273123
rect 403312 273111 403318 273123
rect 363434 273083 403318 273111
rect 363434 273071 363440 273083
rect 403312 273071 403318 273083
rect 403370 273071 403376 273123
rect 501232 273071 501238 273123
rect 501290 273111 501296 273123
rect 617680 273111 617686 273123
rect 501290 273083 617686 273111
rect 501290 273071 501296 273083
rect 617680 273071 617686 273083
rect 617738 273071 617744 273123
rect 139600 272997 139606 273049
rect 139658 273037 139664 273049
rect 139658 273009 146654 273037
rect 139658 272997 139664 273009
rect 68176 272849 68182 272901
rect 68234 272889 68240 272901
rect 69040 272889 69046 272901
rect 68234 272861 69046 272889
rect 68234 272849 68240 272861
rect 69040 272849 69046 272861
rect 69098 272849 69104 272901
rect 75376 272849 75382 272901
rect 75434 272889 75440 272901
rect 77680 272889 77686 272901
rect 75434 272861 77686 272889
rect 75434 272849 75440 272861
rect 77680 272849 77686 272861
rect 77738 272849 77744 272901
rect 98032 272849 98038 272901
rect 98090 272889 98096 272901
rect 100720 272889 100726 272901
rect 98090 272861 100726 272889
rect 98090 272849 98096 272861
rect 100720 272849 100726 272861
rect 100778 272849 100784 272901
rect 101488 272849 101494 272901
rect 101546 272889 101552 272901
rect 103600 272889 103606 272901
rect 101546 272861 103606 272889
rect 101546 272849 101552 272861
rect 103600 272849 103606 272861
rect 103658 272849 103664 272901
rect 115792 272849 115798 272901
rect 115850 272889 115856 272901
rect 118000 272889 118006 272901
rect 115850 272861 118006 272889
rect 115850 272849 115856 272861
rect 118000 272849 118006 272861
rect 118058 272849 118064 272901
rect 119344 272849 119350 272901
rect 119402 272889 119408 272901
rect 120880 272889 120886 272901
rect 119402 272861 120886 272889
rect 119402 272849 119408 272861
rect 120880 272849 120886 272861
rect 120938 272849 120944 272901
rect 122896 272849 122902 272901
rect 122954 272889 122960 272901
rect 123760 272889 123766 272901
rect 122954 272861 123766 272889
rect 122954 272849 122960 272861
rect 123760 272849 123766 272861
rect 123818 272849 123824 272901
rect 130096 272849 130102 272901
rect 130154 272889 130160 272901
rect 132400 272889 132406 272901
rect 130154 272861 132406 272889
rect 130154 272849 130160 272861
rect 132400 272849 132406 272861
rect 132458 272849 132464 272901
rect 133552 272849 133558 272901
rect 133610 272889 133616 272901
rect 135280 272889 135286 272901
rect 133610 272861 135286 272889
rect 133610 272849 133616 272861
rect 135280 272849 135286 272861
rect 135338 272849 135344 272901
rect 137200 272849 137206 272901
rect 137258 272889 137264 272901
rect 138160 272889 138166 272901
rect 137258 272861 138166 272889
rect 137258 272849 137264 272861
rect 138160 272849 138166 272861
rect 138218 272849 138224 272901
rect 138352 272849 138358 272901
rect 138410 272889 138416 272901
rect 140944 272889 140950 272901
rect 138410 272861 140950 272889
rect 138410 272849 138416 272861
rect 140944 272849 140950 272861
rect 141002 272849 141008 272901
rect 142000 272849 142006 272901
rect 142058 272889 142064 272901
rect 143920 272889 143926 272901
rect 142058 272861 143926 272889
rect 142058 272849 142064 272861
rect 143920 272849 143926 272861
rect 143978 272849 143984 272901
rect 146626 272889 146654 273009
rect 178480 272997 178486 273049
rect 178538 273037 178544 273049
rect 302416 273037 302422 273049
rect 178538 273009 302422 273037
rect 178538 272997 178544 273009
rect 302416 272997 302422 273009
rect 302474 272997 302480 273049
rect 322480 272997 322486 273049
rect 322538 273037 322544 273049
rect 339568 273037 339574 273049
rect 322538 273009 339574 273037
rect 322538 272997 322544 273009
rect 339568 272997 339574 273009
rect 339626 272997 339632 273049
rect 339760 272997 339766 273049
rect 339818 273037 339824 273049
rect 362896 273037 362902 273049
rect 339818 273009 362902 273037
rect 339818 272997 339824 273009
rect 362896 272997 362902 273009
rect 362954 272997 362960 273049
rect 379504 273037 379510 273049
rect 363106 273009 379510 273037
rect 146704 272923 146710 272975
rect 146762 272963 146768 272975
rect 158800 272963 158806 272975
rect 146762 272935 158806 272963
rect 146762 272923 146768 272935
rect 158800 272923 158806 272935
rect 158858 272923 158864 272975
rect 279376 272963 279382 272975
rect 158914 272935 279382 272963
rect 158914 272889 158942 272935
rect 279376 272923 279382 272935
rect 279434 272923 279440 272975
rect 279568 272923 279574 272975
rect 279626 272963 279632 272975
rect 363106 272963 363134 273009
rect 379504 272997 379510 273009
rect 379562 272997 379568 273049
rect 379600 272997 379606 273049
rect 379658 273037 379664 273049
rect 398608 273037 398614 273049
rect 379658 273009 398614 273037
rect 379658 272997 379664 273009
rect 398608 272997 398614 273009
rect 398666 272997 398672 273049
rect 540400 273037 540406 273049
rect 398914 273009 540406 273037
rect 279626 272935 363134 272963
rect 279626 272923 279632 272935
rect 363184 272923 363190 272975
rect 363242 272963 363248 272975
rect 363242 272935 378302 272963
rect 363242 272923 363248 272935
rect 146626 272861 158942 272889
rect 161200 272849 161206 272901
rect 161258 272889 161264 272901
rect 378160 272889 378166 272901
rect 161258 272861 378166 272889
rect 161258 272849 161264 272861
rect 378160 272849 378166 272861
rect 378218 272849 378224 272901
rect 378274 272889 378302 272935
rect 378736 272923 378742 272975
rect 378794 272963 378800 272975
rect 394192 272963 394198 272975
rect 378794 272935 394198 272963
rect 378794 272923 378800 272935
rect 394192 272923 394198 272935
rect 394250 272923 394256 272975
rect 394384 272923 394390 272975
rect 394442 272963 394448 272975
rect 398914 272963 398942 273009
rect 540400 272997 540406 273009
rect 540458 272997 540464 273049
rect 394442 272935 398942 272963
rect 394442 272923 394448 272935
rect 398992 272923 398998 272975
rect 399050 272963 399056 272975
rect 407632 272963 407638 272975
rect 399050 272935 407638 272963
rect 399050 272923 399056 272935
rect 407632 272923 407638 272935
rect 407690 272923 407696 272975
rect 407728 272923 407734 272975
rect 407786 272963 407792 272975
rect 533200 272963 533206 272975
rect 407786 272935 533206 272963
rect 407786 272923 407792 272935
rect 533200 272923 533206 272935
rect 533258 272923 533264 272975
rect 378928 272889 378934 272901
rect 378274 272861 378934 272889
rect 378928 272849 378934 272861
rect 378986 272849 378992 272901
rect 379138 272861 379262 272889
rect 135952 272775 135958 272827
rect 136010 272815 136016 272827
rect 370384 272815 370390 272827
rect 136010 272787 370390 272815
rect 136010 272775 136016 272787
rect 370384 272775 370390 272787
rect 370442 272775 370448 272827
rect 373072 272775 373078 272827
rect 373130 272815 373136 272827
rect 379138 272815 379166 272861
rect 373130 272787 378686 272815
rect 373130 272775 373136 272787
rect 128944 272701 128950 272753
rect 129002 272741 129008 272753
rect 160528 272741 160534 272753
rect 129002 272713 160534 272741
rect 129002 272701 129008 272713
rect 160528 272701 160534 272713
rect 160586 272701 160592 272753
rect 161200 272701 161206 272753
rect 161258 272741 161264 272753
rect 378544 272741 378550 272753
rect 161258 272713 378550 272741
rect 161258 272701 161264 272713
rect 378544 272701 378550 272713
rect 378602 272701 378608 272753
rect 378658 272741 378686 272787
rect 378946 272787 379166 272815
rect 379234 272815 379262 272861
rect 379312 272849 379318 272901
rect 379370 272889 379376 272901
rect 388720 272889 388726 272901
rect 379370 272861 388726 272889
rect 379370 272849 379376 272861
rect 388720 272849 388726 272861
rect 388778 272849 388784 272901
rect 388816 272849 388822 272901
rect 388874 272889 388880 272901
rect 388874 272861 392606 272889
rect 388874 272849 388880 272861
rect 392464 272815 392470 272827
rect 379234 272787 392470 272815
rect 378946 272741 378974 272787
rect 392464 272775 392470 272787
rect 392522 272775 392528 272827
rect 392578 272815 392606 272861
rect 394480 272849 394486 272901
rect 394538 272889 394544 272901
rect 518992 272889 518998 272901
rect 394538 272861 518998 272889
rect 394538 272849 394544 272861
rect 518992 272849 518998 272861
rect 519050 272849 519056 272901
rect 407536 272815 407542 272827
rect 392578 272787 407542 272815
rect 407536 272775 407542 272787
rect 407594 272775 407600 272827
rect 407632 272775 407638 272827
rect 407690 272815 407696 272827
rect 522544 272815 522550 272827
rect 407690 272787 522550 272815
rect 407690 272775 407696 272787
rect 522544 272775 522550 272787
rect 522602 272775 522608 272827
rect 391696 272741 391702 272753
rect 378658 272713 378974 272741
rect 379042 272713 391702 272741
rect 105040 272627 105046 272679
rect 105098 272667 105104 272679
rect 106480 272667 106486 272679
rect 105098 272639 106486 272667
rect 105098 272627 105104 272639
rect 106480 272627 106486 272639
rect 106538 272627 106544 272679
rect 114640 272627 114646 272679
rect 114698 272667 114704 272679
rect 114698 272639 118046 272667
rect 114698 272627 114704 272639
rect 111088 272479 111094 272531
rect 111146 272519 111152 272531
rect 118018 272519 118046 272639
rect 125296 272627 125302 272679
rect 125354 272667 125360 272679
rect 377968 272667 377974 272679
rect 125354 272639 377974 272667
rect 125354 272627 125360 272639
rect 377968 272627 377974 272639
rect 378026 272627 378032 272679
rect 378352 272627 378358 272679
rect 378410 272667 378416 272679
rect 378410 272639 378782 272667
rect 378410 272627 378416 272639
rect 118096 272553 118102 272605
rect 118154 272593 118160 272605
rect 378640 272593 378646 272605
rect 118154 272565 378646 272593
rect 118154 272553 118160 272565
rect 378640 272553 378646 272565
rect 378698 272553 378704 272605
rect 378754 272593 378782 272639
rect 378832 272627 378838 272679
rect 378890 272667 378896 272679
rect 379042 272667 379070 272713
rect 391696 272701 391702 272713
rect 391754 272701 391760 272753
rect 391792 272701 391798 272753
rect 391850 272741 391856 272753
rect 396016 272741 396022 272753
rect 391850 272713 396022 272741
rect 391850 272701 391856 272713
rect 396016 272701 396022 272713
rect 396074 272701 396080 272753
rect 396112 272701 396118 272753
rect 396170 272741 396176 272753
rect 504688 272741 504694 272753
rect 396170 272713 504694 272741
rect 396170 272701 396176 272713
rect 504688 272701 504694 272713
rect 504746 272701 504752 272753
rect 402352 272667 402358 272679
rect 378890 272639 379070 272667
rect 379138 272639 402358 272667
rect 378890 272627 378896 272639
rect 379138 272593 379166 272639
rect 402352 272627 402358 272639
rect 402410 272627 402416 272679
rect 418960 272627 418966 272679
rect 419018 272667 419024 272679
rect 501136 272667 501142 272679
rect 419018 272639 501142 272667
rect 419018 272627 419024 272639
rect 501136 272627 501142 272639
rect 501194 272627 501200 272679
rect 505264 272627 505270 272679
rect 505322 272667 505328 272679
rect 621232 272667 621238 272679
rect 505322 272639 621238 272667
rect 505322 272627 505328 272639
rect 621232 272627 621238 272639
rect 621290 272627 621296 272679
rect 390928 272593 390934 272605
rect 378754 272565 379166 272593
rect 379234 272565 390934 272593
rect 379024 272519 379030 272531
rect 111146 272491 117854 272519
rect 118018 272491 379030 272519
rect 111146 272479 111152 272491
rect 103888 272405 103894 272457
rect 103946 272445 103952 272457
rect 117826 272445 117854 272491
rect 379024 272479 379030 272491
rect 379082 272479 379088 272531
rect 373072 272445 373078 272457
rect 103946 272417 116606 272445
rect 117826 272417 373078 272445
rect 103946 272405 103952 272417
rect 116578 272371 116606 272417
rect 373072 272405 373078 272417
rect 373130 272405 373136 272457
rect 373168 272405 373174 272457
rect 373226 272445 373232 272457
rect 378352 272445 378358 272457
rect 373226 272417 378358 272445
rect 373226 272405 373232 272417
rect 378352 272405 378358 272417
rect 378410 272405 378416 272457
rect 379234 272445 379262 272565
rect 390928 272553 390934 272565
rect 390986 272553 390992 272605
rect 404944 272593 404950 272605
rect 391042 272565 404950 272593
rect 379312 272479 379318 272531
rect 379370 272519 379376 272531
rect 389872 272519 389878 272531
rect 379370 272491 389878 272519
rect 379370 272479 379376 272491
rect 389872 272479 389878 272491
rect 389930 272479 389936 272531
rect 389968 272479 389974 272531
rect 390026 272519 390032 272531
rect 391042 272519 391070 272565
rect 404944 272553 404950 272565
rect 405002 272553 405008 272605
rect 405040 272553 405046 272605
rect 405098 272593 405104 272605
rect 497584 272593 497590 272605
rect 405098 272565 497590 272593
rect 405098 272553 405104 272565
rect 497584 272553 497590 272565
rect 497642 272553 497648 272605
rect 497680 272553 497686 272605
rect 497738 272593 497744 272605
rect 614224 272593 614230 272605
rect 497738 272565 614230 272593
rect 497738 272553 497744 272565
rect 614224 272553 614230 272565
rect 614282 272553 614288 272605
rect 390026 272491 391070 272519
rect 390026 272479 390032 272491
rect 393136 272479 393142 272531
rect 393194 272519 393200 272531
rect 526096 272519 526102 272531
rect 393194 272491 526102 272519
rect 393194 272479 393200 272491
rect 526096 272479 526102 272491
rect 526154 272479 526160 272531
rect 378562 272417 379262 272445
rect 378562 272371 378590 272417
rect 379792 272405 379798 272457
rect 379850 272445 379856 272457
rect 398800 272445 398806 272457
rect 379850 272417 398806 272445
rect 379850 272405 379856 272417
rect 398800 272405 398806 272417
rect 398858 272405 398864 272457
rect 529744 272445 529750 272457
rect 398914 272417 529750 272445
rect 116578 272343 378590 272371
rect 378658 272343 391934 272371
rect 107440 272257 107446 272309
rect 107498 272297 107504 272309
rect 107498 272269 370334 272297
rect 107498 272257 107504 272269
rect 99184 272183 99190 272235
rect 99242 272223 99248 272235
rect 370192 272223 370198 272235
rect 99242 272195 370198 272223
rect 99242 272183 99248 272195
rect 370192 272183 370198 272195
rect 370250 272183 370256 272235
rect 370306 272223 370334 272269
rect 370384 272257 370390 272309
rect 370442 272297 370448 272309
rect 378658 272297 378686 272343
rect 370442 272269 378686 272297
rect 378754 272269 379358 272297
rect 370442 272257 370448 272269
rect 378544 272223 378550 272235
rect 370306 272195 378550 272223
rect 378544 272183 378550 272195
rect 378602 272183 378608 272235
rect 378640 272183 378646 272235
rect 378698 272223 378704 272235
rect 378754 272223 378782 272269
rect 378698 272195 378782 272223
rect 378698 272183 378704 272195
rect 378928 272183 378934 272235
rect 378986 272223 378992 272235
rect 379330 272223 379358 272269
rect 379504 272257 379510 272309
rect 379562 272297 379568 272309
rect 391906 272297 391934 272343
rect 391984 272331 391990 272383
rect 392042 272371 392048 272383
rect 398914 272371 398942 272417
rect 529744 272405 529750 272417
rect 529802 272405 529808 272457
rect 392042 272343 398942 272371
rect 392042 272331 392048 272343
rect 398992 272331 398998 272383
rect 399050 272371 399056 272383
rect 399050 272343 401534 272371
rect 399050 272331 399056 272343
rect 399184 272297 399190 272309
rect 379562 272269 391262 272297
rect 391906 272269 399190 272297
rect 379562 272257 379568 272269
rect 391234 272223 391262 272269
rect 399184 272257 399190 272269
rect 399242 272257 399248 272309
rect 399856 272257 399862 272309
rect 399914 272297 399920 272309
rect 399914 272269 401438 272297
rect 399914 272257 399920 272269
rect 399664 272223 399670 272235
rect 378986 272195 379262 272223
rect 379330 272195 390782 272223
rect 391234 272195 399670 272223
rect 378986 272183 378992 272195
rect 84880 272109 84886 272161
rect 84938 272149 84944 272161
rect 86320 272149 86326 272161
rect 84938 272121 86326 272149
rect 84938 272109 84944 272121
rect 86320 272109 86326 272121
rect 86378 272109 86384 272161
rect 100336 272109 100342 272161
rect 100394 272149 100400 272161
rect 379120 272149 379126 272161
rect 100394 272121 379126 272149
rect 100394 272109 100400 272121
rect 379120 272109 379126 272121
rect 379178 272109 379184 272161
rect 379234 272149 379262 272195
rect 390754 272149 390782 272195
rect 399664 272183 399670 272195
rect 399722 272183 399728 272235
rect 400624 272149 400630 272161
rect 379234 272121 390686 272149
rect 390754 272121 400630 272149
rect 89584 272035 89590 272087
rect 89642 272075 89648 272087
rect 92080 272075 92086 272087
rect 89642 272047 92086 272075
rect 89642 272035 89648 272047
rect 92080 272035 92086 272047
rect 92138 272035 92144 272087
rect 145552 272035 145558 272087
rect 145610 272075 145616 272087
rect 146704 272075 146710 272087
rect 145610 272047 146710 272075
rect 145610 272035 145616 272047
rect 146704 272035 146710 272047
rect 146762 272035 146768 272087
rect 150256 272035 150262 272087
rect 150314 272075 150320 272087
rect 164272 272075 164278 272087
rect 150314 272047 164278 272075
rect 150314 272035 150320 272047
rect 164272 272035 164278 272047
rect 164330 272035 164336 272087
rect 165808 272035 165814 272087
rect 165866 272075 165872 272087
rect 166960 272075 166966 272087
rect 165866 272047 166966 272075
rect 165866 272035 165872 272047
rect 166960 272035 166966 272047
rect 167018 272035 167024 272087
rect 170512 272035 170518 272087
rect 170570 272075 170576 272087
rect 172720 272075 172726 272087
rect 170570 272047 172726 272075
rect 170570 272035 170576 272047
rect 172720 272035 172726 272047
rect 172778 272035 172784 272087
rect 174064 272035 174070 272087
rect 174122 272075 174128 272087
rect 175504 272075 175510 272087
rect 174122 272047 175510 272075
rect 174122 272035 174128 272047
rect 175504 272035 175510 272047
rect 175562 272035 175568 272087
rect 177616 272035 177622 272087
rect 177674 272075 177680 272087
rect 178384 272075 178390 272087
rect 177674 272047 178390 272075
rect 177674 272035 177680 272047
rect 178384 272035 178390 272047
rect 178442 272035 178448 272087
rect 180016 272035 180022 272087
rect 180074 272075 180080 272087
rect 181360 272075 181366 272087
rect 180074 272047 181366 272075
rect 180074 272035 180080 272047
rect 181360 272035 181366 272047
rect 181418 272035 181424 272087
rect 181456 272035 181462 272087
rect 181514 272075 181520 272087
rect 390544 272075 390550 272087
rect 181514 272047 390550 272075
rect 181514 272035 181520 272047
rect 390544 272035 390550 272047
rect 390602 272035 390608 272087
rect 390658 272075 390686 272121
rect 400624 272109 400630 272121
rect 400682 272109 400688 272161
rect 401296 272075 401302 272087
rect 390658 272047 401302 272075
rect 401296 272035 401302 272047
rect 401354 272035 401360 272087
rect 401410 272075 401438 272269
rect 401506 272223 401534 272343
rect 401584 272331 401590 272383
rect 401642 272371 401648 272383
rect 547600 272371 547606 272383
rect 401642 272343 547606 272371
rect 401642 272331 401648 272343
rect 547600 272331 547606 272343
rect 547658 272331 547664 272383
rect 560080 272331 560086 272383
rect 560138 272371 560144 272383
rect 643888 272371 643894 272383
rect 560138 272343 643894 272371
rect 560138 272331 560144 272343
rect 643888 272331 643894 272343
rect 643946 272331 643952 272383
rect 406000 272257 406006 272309
rect 406058 272297 406064 272309
rect 418960 272297 418966 272309
rect 406058 272269 418966 272297
rect 406058 272257 406064 272269
rect 418960 272257 418966 272269
rect 419018 272257 419024 272309
rect 486736 272257 486742 272309
rect 486794 272297 486800 272309
rect 641488 272297 641494 272309
rect 486794 272269 641494 272297
rect 486794 272257 486800 272269
rect 641488 272257 641494 272269
rect 641546 272257 641552 272309
rect 407728 272223 407734 272235
rect 401506 272195 407734 272223
rect 407728 272183 407734 272195
rect 407786 272183 407792 272235
rect 480976 272183 480982 272235
rect 481034 272223 481040 272235
rect 634288 272223 634294 272235
rect 481034 272195 634294 272223
rect 481034 272183 481040 272195
rect 634288 272183 634294 272195
rect 634346 272183 634352 272235
rect 406096 272109 406102 272161
rect 406154 272149 406160 272161
rect 609424 272149 609430 272161
rect 406154 272121 609430 272149
rect 406154 272109 406160 272121
rect 609424 272109 609430 272121
rect 609482 272109 609488 272161
rect 406768 272075 406774 272087
rect 401410 272047 406774 272075
rect 406768 272035 406774 272047
rect 406826 272035 406832 272087
rect 409072 272035 409078 272087
rect 409130 272075 409136 272087
rect 486832 272075 486838 272087
rect 409130 272047 486838 272075
rect 409130 272035 409136 272047
rect 486832 272035 486838 272047
rect 486890 272035 486896 272087
rect 164560 271961 164566 272013
rect 164618 272001 164624 272013
rect 405520 272001 405526 272013
rect 164618 271973 405526 272001
rect 164618 271961 164624 271973
rect 405520 271961 405526 271973
rect 405578 271961 405584 272013
rect 411280 271961 411286 272013
rect 411338 272001 411344 272013
rect 468976 272001 468982 272013
rect 411338 271973 468982 272001
rect 411338 271961 411344 271973
rect 468976 271961 468982 271973
rect 469034 271961 469040 272013
rect 172912 271887 172918 271939
rect 172970 271927 172976 271939
rect 175600 271927 175606 271939
rect 172970 271899 175606 271927
rect 172970 271887 172976 271899
rect 175600 271887 175606 271899
rect 175658 271887 175664 271939
rect 176464 271887 176470 271939
rect 176522 271927 176528 271939
rect 178480 271927 178486 271939
rect 176522 271899 178486 271927
rect 176522 271887 176528 271899
rect 178480 271887 178486 271899
rect 178538 271887 178544 271939
rect 179440 271887 179446 271939
rect 179498 271927 179504 271939
rect 388816 271927 388822 271939
rect 179498 271899 388822 271927
rect 179498 271887 179504 271899
rect 388816 271887 388822 271899
rect 388874 271887 388880 271939
rect 388912 271887 388918 271939
rect 388970 271927 388976 271939
rect 408208 271927 408214 271939
rect 388970 271899 408214 271927
rect 388970 271887 388976 271899
rect 408208 271887 408214 271899
rect 408266 271887 408272 271939
rect 106288 271813 106294 271865
rect 106346 271853 106352 271865
rect 106346 271825 190718 271853
rect 106346 271813 106352 271825
rect 109840 271739 109846 271791
rect 109898 271779 109904 271791
rect 190576 271779 190582 271791
rect 109898 271751 190582 271779
rect 109898 271739 109904 271751
rect 190576 271739 190582 271751
rect 190634 271739 190640 271791
rect 190690 271779 190718 271825
rect 190768 271813 190774 271865
rect 190826 271853 190832 271865
rect 192880 271853 192886 271865
rect 190826 271825 192886 271853
rect 190826 271813 190832 271825
rect 192880 271813 192886 271825
rect 192938 271813 192944 271865
rect 209680 271813 209686 271865
rect 209738 271853 209744 271865
rect 213232 271853 213238 271865
rect 209738 271825 213238 271853
rect 209738 271813 209744 271825
rect 213232 271813 213238 271825
rect 213290 271813 213296 271865
rect 232432 271813 232438 271865
rect 232490 271853 232496 271865
rect 271216 271853 271222 271865
rect 232490 271825 271222 271853
rect 232490 271813 232496 271825
rect 271216 271813 271222 271825
rect 271274 271813 271280 271865
rect 271600 271813 271606 271865
rect 271658 271853 271664 271865
rect 279472 271853 279478 271865
rect 271658 271825 279478 271853
rect 271658 271813 271664 271825
rect 279472 271813 279478 271825
rect 279530 271813 279536 271865
rect 283792 271813 283798 271865
rect 283850 271853 283856 271865
rect 307312 271853 307318 271865
rect 283850 271825 307318 271853
rect 283850 271813 283856 271825
rect 307312 271813 307318 271825
rect 307370 271813 307376 271865
rect 312112 271813 312118 271865
rect 312170 271853 312176 271865
rect 321616 271853 321622 271865
rect 312170 271825 321622 271853
rect 312170 271813 312176 271825
rect 321616 271813 321622 271825
rect 321674 271813 321680 271865
rect 549904 271853 549910 271865
rect 321730 271825 549910 271853
rect 205840 271779 205846 271791
rect 190690 271751 205846 271779
rect 205840 271739 205846 271751
rect 205898 271739 205904 271791
rect 220816 271739 220822 271791
rect 220874 271779 220880 271791
rect 245488 271779 245494 271791
rect 220874 271751 245494 271779
rect 220874 271739 220880 271751
rect 245488 271739 245494 271751
rect 245546 271739 245552 271791
rect 250192 271739 250198 271791
rect 250250 271779 250256 271791
rect 267952 271779 267958 271791
rect 250250 271751 267958 271779
rect 250250 271739 250256 271751
rect 267952 271739 267958 271751
rect 268010 271739 268016 271791
rect 268048 271739 268054 271791
rect 268106 271779 268112 271791
rect 278992 271779 278998 271791
rect 268106 271751 278998 271779
rect 268106 271739 268112 271751
rect 278992 271739 278998 271751
rect 279050 271739 279056 271791
rect 283408 271739 283414 271791
rect 283466 271779 283472 271791
rect 303664 271779 303670 271791
rect 283466 271751 303670 271779
rect 283466 271739 283472 271751
rect 303664 271739 303670 271751
rect 303722 271739 303728 271791
rect 313648 271739 313654 271791
rect 313706 271779 313712 271791
rect 321730 271779 321758 271825
rect 549904 271813 549910 271825
rect 549962 271813 549968 271865
rect 313706 271751 321758 271779
rect 313706 271739 313712 271751
rect 321808 271739 321814 271791
rect 321866 271779 321872 271791
rect 329872 271779 329878 271791
rect 321866 271751 329878 271779
rect 321866 271739 321872 271751
rect 329872 271739 329878 271751
rect 329930 271739 329936 271791
rect 329968 271739 329974 271791
rect 330026 271779 330032 271791
rect 341776 271779 341782 271791
rect 330026 271751 341782 271779
rect 330026 271739 330032 271751
rect 341776 271739 341782 271751
rect 341834 271739 341840 271791
rect 347248 271739 347254 271791
rect 347306 271779 347312 271791
rect 358480 271779 358486 271791
rect 347306 271751 358486 271779
rect 347306 271739 347312 271751
rect 358480 271739 358486 271751
rect 358538 271739 358544 271791
rect 358576 271739 358582 271791
rect 358634 271779 358640 271791
rect 374416 271779 374422 271791
rect 358634 271751 374422 271779
rect 358634 271739 358640 271751
rect 374416 271739 374422 271751
rect 374474 271739 374480 271791
rect 375568 271739 375574 271791
rect 375626 271779 375632 271791
rect 378064 271779 378070 271791
rect 375626 271751 378070 271779
rect 375626 271739 375632 271751
rect 378064 271739 378070 271751
rect 378122 271739 378128 271791
rect 378160 271739 378166 271791
rect 378218 271779 378224 271791
rect 388624 271779 388630 271791
rect 378218 271751 388630 271779
rect 378218 271739 378224 271751
rect 388624 271739 388630 271751
rect 388682 271739 388688 271791
rect 388720 271739 388726 271791
rect 388778 271779 388784 271791
rect 608176 271779 608182 271791
rect 388778 271751 608182 271779
rect 388778 271739 388784 271751
rect 608176 271739 608182 271751
rect 608234 271739 608240 271791
rect 171664 271665 171670 271717
rect 171722 271705 171728 271717
rect 179440 271705 179446 271717
rect 171722 271677 179446 271705
rect 171722 271665 171728 271677
rect 179440 271665 179446 271677
rect 179498 271665 179504 271717
rect 388816 271705 388822 271717
rect 181090 271677 388822 271705
rect 175312 271591 175318 271643
rect 175370 271631 175376 271643
rect 181090 271631 181118 271677
rect 388816 271665 388822 271677
rect 388874 271665 388880 271717
rect 388912 271665 388918 271717
rect 388970 271705 388976 271717
rect 396208 271705 396214 271717
rect 388970 271677 396214 271705
rect 388970 271665 388976 271677
rect 396208 271665 396214 271677
rect 396266 271665 396272 271717
rect 397360 271665 397366 271717
rect 397418 271705 397424 271717
rect 405040 271705 405046 271717
rect 397418 271677 405046 271705
rect 397418 271665 397424 271677
rect 405040 271665 405046 271677
rect 405098 271665 405104 271717
rect 409264 271631 409270 271643
rect 175370 271603 181118 271631
rect 182338 271603 409270 271631
rect 175370 271591 175376 271603
rect 141136 271517 141142 271569
rect 141194 271557 141200 271569
rect 147184 271557 147190 271569
rect 141194 271529 147190 271557
rect 141194 271517 141200 271529
rect 147184 271517 147190 271529
rect 147242 271517 147248 271569
rect 178864 271517 178870 271569
rect 178922 271557 178928 271569
rect 182338 271557 182366 271603
rect 409264 271591 409270 271603
rect 409322 271591 409328 271643
rect 178922 271529 182366 271557
rect 178922 271517 178928 271529
rect 182416 271517 182422 271569
rect 182474 271557 182480 271569
rect 409936 271557 409942 271569
rect 182474 271529 409942 271557
rect 182474 271517 182480 271529
rect 409936 271517 409942 271529
rect 409994 271517 410000 271569
rect 124144 271443 124150 271495
rect 124202 271483 124208 271495
rect 212176 271483 212182 271495
rect 124202 271455 212182 271483
rect 124202 271443 124208 271455
rect 212176 271443 212182 271455
rect 212234 271443 212240 271495
rect 246640 271443 246646 271495
rect 246698 271483 246704 271495
rect 276112 271483 276118 271495
rect 246698 271455 276118 271483
rect 246698 271443 246704 271455
rect 276112 271443 276118 271455
rect 276170 271443 276176 271495
rect 282736 271443 282742 271495
rect 282794 271483 282800 271495
rect 296656 271483 296662 271495
rect 282794 271455 296662 271483
rect 282794 271443 282800 271455
rect 296656 271443 296662 271455
rect 296714 271443 296720 271495
rect 308464 271443 308470 271495
rect 308522 271483 308528 271495
rect 321808 271483 321814 271495
rect 308522 271455 321814 271483
rect 308522 271443 308528 271455
rect 321808 271443 321814 271455
rect 321866 271443 321872 271495
rect 323056 271443 323062 271495
rect 323114 271483 323120 271495
rect 325552 271483 325558 271495
rect 323114 271455 325558 271483
rect 323114 271443 323120 271455
rect 325552 271443 325558 271455
rect 325610 271443 325616 271495
rect 325648 271443 325654 271495
rect 325706 271483 325712 271495
rect 328048 271483 328054 271495
rect 325706 271455 328054 271483
rect 325706 271443 325712 271455
rect 328048 271443 328054 271455
rect 328106 271443 328112 271495
rect 328144 271443 328150 271495
rect 328202 271483 328208 271495
rect 329008 271483 329014 271495
rect 328202 271455 329014 271483
rect 328202 271443 328208 271455
rect 329008 271443 329014 271455
rect 329066 271443 329072 271495
rect 329872 271443 329878 271495
rect 329930 271483 329936 271495
rect 339376 271483 339382 271495
rect 329930 271455 339382 271483
rect 329930 271443 329936 271455
rect 339376 271443 339382 271455
rect 339434 271443 339440 271495
rect 346768 271443 346774 271495
rect 346826 271483 346832 271495
rect 349648 271483 349654 271495
rect 346826 271455 349654 271483
rect 346826 271443 346832 271455
rect 349648 271443 349654 271455
rect 349706 271443 349712 271495
rect 349744 271443 349750 271495
rect 349802 271483 349808 271495
rect 358576 271483 358582 271495
rect 349802 271455 358582 271483
rect 349802 271443 349808 271455
rect 358576 271443 358582 271455
rect 358634 271443 358640 271495
rect 362992 271443 362998 271495
rect 363050 271483 363056 271495
rect 365392 271483 365398 271495
rect 363050 271455 365398 271483
rect 363050 271443 363056 271455
rect 365392 271443 365398 271455
rect 365450 271443 365456 271495
rect 370000 271443 370006 271495
rect 370058 271483 370064 271495
rect 383248 271483 383254 271495
rect 370058 271455 383254 271483
rect 370058 271443 370064 271455
rect 383248 271443 383254 271455
rect 383306 271443 383312 271495
rect 383344 271443 383350 271495
rect 383402 271483 383408 271495
rect 601072 271483 601078 271495
rect 383402 271455 601078 271483
rect 383402 271443 383408 271455
rect 601072 271443 601078 271455
rect 601130 271443 601136 271495
rect 127696 271369 127702 271421
rect 127754 271409 127760 271421
rect 141136 271409 141142 271421
rect 127754 271381 141142 271409
rect 127754 271369 127760 271381
rect 141136 271369 141142 271381
rect 141194 271369 141200 271421
rect 151408 271369 151414 271421
rect 151466 271409 151472 271421
rect 152560 271409 152566 271421
rect 151466 271381 152566 271409
rect 151466 271369 151472 271381
rect 152560 271369 152566 271381
rect 152618 271369 152624 271421
rect 190576 271369 190582 271421
rect 190634 271409 190640 271421
rect 206992 271409 206998 271421
rect 190634 271381 206998 271409
rect 190634 271369 190640 271381
rect 206992 271369 206998 271381
rect 207050 271369 207056 271421
rect 207088 271369 207094 271421
rect 207146 271409 207152 271421
rect 411952 271409 411958 271421
rect 207146 271381 411958 271409
rect 207146 271369 207152 271381
rect 411952 271369 411958 271381
rect 412010 271369 412016 271421
rect 131248 271295 131254 271347
rect 131306 271335 131312 271347
rect 131306 271307 146750 271335
rect 131306 271295 131312 271307
rect 134800 270999 134806 271051
rect 134858 271039 134864 271051
rect 134858 271011 141182 271039
rect 134858 270999 134864 271011
rect 141154 270817 141182 271011
rect 146722 270965 146750 271307
rect 168112 271295 168118 271347
rect 168170 271335 168176 271347
rect 181456 271335 181462 271347
rect 168170 271307 181462 271335
rect 168170 271295 168176 271307
rect 181456 271295 181462 271307
rect 181514 271295 181520 271347
rect 185968 271295 185974 271347
rect 186026 271335 186032 271347
rect 410992 271335 410998 271347
rect 186026 271307 410998 271335
rect 186026 271295 186032 271307
rect 410992 271295 410998 271307
rect 411050 271295 411056 271347
rect 147184 271221 147190 271273
rect 147242 271261 147248 271273
rect 177040 271261 177046 271273
rect 147242 271233 177046 271261
rect 147242 271221 147248 271233
rect 177040 271221 177046 271233
rect 177098 271221 177104 271273
rect 184720 271221 184726 271273
rect 184778 271261 184784 271273
rect 187024 271261 187030 271273
rect 184778 271233 187030 271261
rect 184778 271221 184784 271233
rect 187024 271221 187030 271233
rect 187082 271221 187088 271273
rect 195184 271221 195190 271273
rect 195242 271261 195248 271273
rect 211888 271261 211894 271273
rect 195242 271233 211894 271261
rect 195242 271221 195248 271233
rect 211888 271221 211894 271233
rect 211946 271221 211952 271273
rect 220336 271221 220342 271273
rect 220394 271261 220400 271273
rect 241840 271261 241846 271273
rect 220394 271233 241846 271261
rect 220394 271221 220400 271233
rect 241840 271221 241846 271233
rect 241898 271221 241904 271273
rect 271216 271221 271222 271273
rect 271274 271261 271280 271273
rect 274672 271261 274678 271273
rect 271274 271233 274678 271261
rect 271274 271221 271280 271233
rect 274672 271221 274678 271233
rect 274730 271221 274736 271273
rect 282928 271221 282934 271273
rect 282986 271261 282992 271273
rect 300112 271261 300118 271273
rect 282986 271233 300118 271261
rect 282986 271221 282992 271233
rect 300112 271221 300118 271233
rect 300170 271221 300176 271273
rect 316336 271221 316342 271273
rect 316394 271261 316400 271273
rect 332272 271261 332278 271273
rect 316394 271233 332278 271261
rect 316394 271221 316400 271233
rect 332272 271221 332278 271233
rect 332330 271221 332336 271273
rect 334096 271221 334102 271273
rect 334154 271261 334160 271273
rect 339856 271261 339862 271273
rect 334154 271233 339862 271261
rect 334154 271221 334160 271233
rect 339856 271221 339862 271233
rect 339914 271221 339920 271273
rect 349552 271221 349558 271273
rect 349610 271261 349616 271273
rect 351184 271261 351190 271273
rect 349610 271233 351190 271261
rect 349610 271221 349616 271233
rect 351184 271221 351190 271233
rect 351242 271221 351248 271273
rect 351280 271221 351286 271273
rect 351338 271261 351344 271273
rect 351338 271233 370142 271261
rect 351338 271221 351344 271233
rect 211696 271187 211702 271199
rect 146914 271159 177086 271187
rect 146914 270965 146942 271159
rect 151120 271073 151126 271125
rect 151178 271113 151184 271125
rect 177058 271113 177086 271159
rect 189538 271159 211702 271187
rect 189538 271113 189566 271159
rect 211696 271147 211702 271159
rect 211754 271147 211760 271199
rect 219760 271147 219766 271199
rect 219818 271187 219824 271199
rect 238288 271187 238294 271199
rect 219818 271159 238294 271187
rect 219818 271147 219824 271159
rect 238288 271147 238294 271159
rect 238346 271147 238352 271199
rect 267952 271147 267958 271199
rect 268010 271187 268016 271199
rect 276784 271187 276790 271199
rect 268010 271159 276790 271187
rect 268010 271147 268016 271159
rect 276784 271147 276790 271159
rect 276842 271147 276848 271199
rect 281200 271147 281206 271199
rect 281258 271187 281264 271199
rect 285808 271187 285814 271199
rect 281258 271159 285814 271187
rect 281258 271147 281264 271159
rect 285808 271147 285814 271159
rect 285866 271147 285872 271199
rect 316816 271147 316822 271199
rect 316874 271187 316880 271199
rect 327184 271187 327190 271199
rect 316874 271159 327190 271187
rect 316874 271147 316880 271159
rect 327184 271147 327190 271159
rect 327242 271147 327248 271199
rect 328336 271147 328342 271199
rect 328394 271187 328400 271199
rect 331216 271187 331222 271199
rect 328394 271159 331222 271187
rect 328394 271147 328400 271159
rect 331216 271147 331222 271159
rect 331274 271147 331280 271199
rect 345712 271147 345718 271199
rect 345770 271187 345776 271199
rect 345770 271159 354974 271187
rect 345770 271147 345776 271159
rect 151178 271085 176990 271113
rect 177058 271085 189566 271113
rect 151178 271073 151184 271085
rect 146722 270937 146942 270965
rect 151120 270817 151126 270829
rect 141154 270789 151126 270817
rect 151120 270777 151126 270789
rect 151178 270777 151184 270829
rect 176962 270817 176990 271085
rect 189616 271073 189622 271125
rect 189674 271113 189680 271125
rect 212080 271113 212086 271125
rect 189674 271085 212086 271113
rect 189674 271073 189680 271085
rect 212080 271073 212086 271085
rect 212138 271073 212144 271125
rect 213040 271073 213046 271125
rect 213098 271113 213104 271125
rect 213098 271085 217406 271113
rect 213098 271073 213104 271085
rect 189520 270999 189526 271051
rect 189578 271039 189584 271051
rect 207088 271039 207094 271051
rect 189578 271011 207094 271039
rect 189578 270999 189584 271011
rect 207088 270999 207094 271011
rect 207146 270999 207152 271051
rect 207184 270999 207190 271051
rect 207242 271039 207248 271051
rect 213808 271039 213814 271051
rect 207242 271011 213814 271039
rect 207242 270999 207248 271011
rect 213808 270999 213814 271011
rect 213866 270999 213872 271051
rect 195472 270925 195478 270977
rect 195530 270965 195536 270977
rect 214480 270965 214486 270977
rect 195530 270937 214486 270965
rect 195530 270925 195536 270937
rect 214480 270925 214486 270937
rect 214538 270925 214544 270977
rect 177040 270851 177046 270903
rect 177098 270891 177104 270903
rect 195184 270891 195190 270903
rect 177098 270863 195190 270891
rect 177098 270851 177104 270863
rect 195184 270851 195190 270863
rect 195242 270851 195248 270903
rect 199120 270851 199126 270903
rect 199178 270891 199184 270903
rect 214960 270891 214966 270903
rect 199178 270863 214966 270891
rect 199178 270851 199184 270863
rect 214960 270851 214966 270863
rect 215018 270851 215024 270903
rect 189616 270817 189622 270829
rect 176962 270789 189622 270817
rect 189616 270777 189622 270789
rect 189674 270777 189680 270829
rect 202576 270777 202582 270829
rect 202634 270817 202640 270829
rect 215440 270817 215446 270829
rect 202634 270789 215446 270817
rect 202634 270777 202640 270789
rect 215440 270777 215446 270789
rect 215498 270777 215504 270829
rect 67600 270703 67606 270755
rect 67658 270743 67664 270755
rect 67658 270715 69182 270743
rect 67658 270703 67664 270715
rect 69154 270669 69182 270715
rect 191920 270703 191926 270755
rect 191978 270743 191984 270755
rect 191978 270715 206174 270743
rect 191978 270703 191984 270715
rect 81808 270669 81814 270681
rect 69154 270641 81814 270669
rect 81808 270629 81814 270641
rect 81866 270629 81872 270681
rect 206146 270669 206174 270715
rect 206224 270703 206230 270755
rect 206282 270743 206288 270755
rect 215536 270743 215542 270755
rect 206282 270715 215542 270743
rect 206282 270703 206288 270715
rect 215536 270703 215542 270715
rect 215594 270703 215600 270755
rect 217378 270743 217406 271085
rect 219280 271073 219286 271125
rect 219338 271113 219344 271125
rect 234640 271113 234646 271125
rect 219338 271085 234646 271113
rect 219338 271073 219344 271085
rect 234640 271073 234646 271085
rect 234698 271073 234704 271125
rect 264496 271073 264502 271125
rect 264554 271113 264560 271125
rect 278512 271113 278518 271125
rect 264554 271085 278518 271113
rect 264554 271073 264560 271085
rect 278512 271073 278518 271085
rect 278570 271073 278576 271125
rect 315664 271073 315670 271125
rect 315722 271113 315728 271125
rect 324592 271113 324598 271125
rect 315722 271085 324598 271113
rect 315722 271073 315728 271085
rect 324592 271073 324598 271085
rect 324650 271073 324656 271125
rect 324688 271073 324694 271125
rect 324746 271113 324752 271125
rect 325648 271113 325654 271125
rect 324746 271085 325654 271113
rect 324746 271073 324752 271085
rect 325648 271073 325654 271085
rect 325706 271073 325712 271125
rect 326320 271073 326326 271125
rect 326378 271113 326384 271125
rect 341488 271113 341494 271125
rect 326378 271085 341494 271113
rect 326378 271073 326384 271085
rect 341488 271073 341494 271085
rect 341546 271073 341552 271125
rect 345232 271073 345238 271125
rect 345290 271113 345296 271125
rect 354832 271113 354838 271125
rect 345290 271085 354838 271113
rect 345290 271073 345296 271085
rect 354832 271073 354838 271085
rect 354890 271073 354896 271125
rect 354946 271113 354974 271159
rect 355216 271147 355222 271199
rect 355274 271187 355280 271199
rect 370000 271187 370006 271199
rect 355274 271159 370006 271187
rect 355274 271147 355280 271159
rect 370000 271147 370006 271159
rect 370058 271147 370064 271199
rect 370114 271187 370142 271233
rect 370192 271221 370198 271273
rect 370250 271261 370256 271273
rect 389392 271261 389398 271273
rect 370250 271233 389398 271261
rect 370250 271221 370256 271233
rect 389392 271221 389398 271233
rect 389450 271221 389456 271273
rect 390448 271221 390454 271273
rect 390506 271261 390512 271273
rect 394384 271261 394390 271273
rect 390506 271233 394390 271261
rect 390506 271221 390512 271233
rect 394384 271221 394390 271233
rect 394442 271221 394448 271273
rect 394480 271221 394486 271273
rect 394538 271261 394544 271273
rect 511888 271261 511894 271273
rect 394538 271233 511894 271261
rect 394538 271221 394544 271233
rect 511888 271221 511894 271233
rect 511946 271221 511952 271273
rect 383152 271187 383158 271199
rect 370114 271159 383158 271187
rect 383152 271147 383158 271159
rect 383210 271147 383216 271199
rect 385456 271147 385462 271199
rect 385514 271187 385520 271199
rect 389296 271187 389302 271199
rect 385514 271159 389302 271187
rect 385514 271147 385520 271159
rect 389296 271147 389302 271159
rect 389354 271147 389360 271199
rect 398032 271187 398038 271199
rect 390274 271159 398038 271187
rect 358384 271113 358390 271125
rect 354946 271085 358390 271113
rect 358384 271073 358390 271085
rect 358442 271073 358448 271125
rect 358480 271073 358486 271125
rect 358538 271113 358544 271125
rect 365008 271113 365014 271125
rect 358538 271085 365014 271113
rect 358538 271073 358544 271085
rect 365008 271073 365014 271085
rect 365066 271073 365072 271125
rect 367024 271073 367030 271125
rect 367082 271113 367088 271125
rect 371920 271113 371926 271125
rect 367082 271085 371926 271113
rect 367082 271073 367088 271085
rect 371920 271073 371926 271085
rect 371978 271073 371984 271125
rect 372880 271073 372886 271125
rect 372938 271113 372944 271125
rect 390274 271113 390302 271159
rect 398032 271147 398038 271159
rect 398090 271147 398096 271199
rect 398224 271147 398230 271199
rect 398282 271187 398288 271199
rect 483280 271187 483286 271199
rect 398282 271159 483286 271187
rect 398282 271147 398288 271159
rect 483280 271147 483286 271159
rect 483338 271147 483344 271199
rect 372938 271085 390302 271113
rect 390370 271085 390590 271113
rect 372938 271073 372944 271085
rect 218896 270999 218902 271051
rect 218954 271039 218960 271051
rect 231184 271039 231190 271051
rect 218954 271011 231190 271039
rect 218954 270999 218960 271011
rect 231184 270999 231190 271011
rect 231242 270999 231248 271051
rect 253744 270999 253750 271051
rect 253802 271039 253808 271051
rect 277264 271039 277270 271051
rect 253802 271011 277270 271039
rect 253802 270999 253808 271011
rect 277264 270999 277270 271011
rect 277322 270999 277328 271051
rect 282160 270999 282166 271051
rect 282218 271039 282224 271051
rect 293008 271039 293014 271051
rect 282218 271011 293014 271039
rect 282218 270999 282224 271011
rect 293008 270999 293014 271011
rect 293066 270999 293072 271051
rect 300208 270999 300214 271051
rect 300266 271039 300272 271051
rect 317968 271039 317974 271051
rect 300266 271011 317974 271039
rect 300266 270999 300272 271011
rect 317968 270999 317974 271011
rect 318026 270999 318032 271051
rect 320368 270999 320374 271051
rect 320426 271039 320432 271051
rect 325360 271039 325366 271051
rect 320426 271011 325366 271039
rect 320426 270999 320432 271011
rect 325360 270999 325366 271011
rect 325418 270999 325424 271051
rect 325552 270999 325558 271051
rect 325610 271039 325616 271051
rect 341296 271039 341302 271051
rect 325610 271011 341302 271039
rect 325610 270999 325616 271011
rect 341296 270999 341302 271011
rect 341354 270999 341360 271051
rect 344752 270999 344758 271051
rect 344810 271039 344816 271051
rect 350992 271039 350998 271051
rect 344810 271011 350998 271039
rect 344810 270999 344816 271011
rect 350992 270999 350998 271011
rect 351050 270999 351056 271051
rect 362992 271039 362998 271051
rect 351106 271011 362998 271039
rect 218704 270925 218710 270977
rect 218762 270965 218768 270977
rect 227632 270965 227638 270977
rect 218762 270937 227638 270965
rect 218762 270925 218768 270937
rect 227632 270925 227638 270937
rect 227690 270925 227696 270977
rect 268720 270925 268726 270977
rect 268778 270965 268784 270977
rect 270544 270965 270550 270977
rect 268778 270937 270550 270965
rect 268778 270925 268784 270937
rect 270544 270925 270550 270937
rect 270602 270925 270608 270977
rect 281680 270925 281686 270977
rect 281738 270965 281744 270977
rect 289456 270965 289462 270977
rect 281738 270937 289462 270965
rect 281738 270925 281744 270937
rect 289456 270925 289462 270937
rect 289514 270925 289520 270977
rect 313840 270925 313846 270977
rect 313898 270965 313904 270977
rect 320464 270965 320470 270977
rect 313898 270937 320470 270965
rect 313898 270925 313904 270937
rect 320464 270925 320470 270937
rect 320522 270925 320528 270977
rect 320560 270925 320566 270977
rect 320618 270965 320624 270977
rect 327952 270965 327958 270977
rect 320618 270937 327958 270965
rect 320618 270925 320624 270937
rect 327952 270925 327958 270937
rect 328010 270925 328016 270977
rect 328048 270925 328054 270977
rect 328106 270965 328112 270977
rect 340432 270965 340438 270977
rect 328106 270937 340438 270965
rect 328106 270925 328112 270937
rect 340432 270925 340438 270937
rect 340490 270925 340496 270977
rect 346384 270925 346390 270977
rect 346442 270965 346448 270977
rect 349552 270965 349558 270977
rect 346442 270937 349558 270965
rect 346442 270925 346448 270937
rect 349552 270925 349558 270937
rect 349610 270925 349616 270977
rect 349648 270925 349654 270977
rect 349706 270965 349712 270977
rect 351106 270965 351134 271011
rect 362992 270999 362998 271011
rect 363050 270999 363056 271051
rect 363088 270999 363094 271051
rect 363146 271039 363152 271051
rect 377968 271039 377974 271051
rect 363146 271011 377974 271039
rect 363146 270999 363152 271011
rect 377968 270999 377974 271011
rect 378026 270999 378032 271051
rect 378064 270999 378070 271051
rect 378122 271039 378128 271051
rect 378122 271011 378878 271039
rect 378122 270999 378128 271011
rect 349706 270937 351134 270965
rect 349706 270925 349712 270937
rect 358480 270925 358486 270977
rect 358538 270965 358544 270977
rect 378850 270965 378878 271011
rect 378928 270999 378934 271051
rect 378986 271039 378992 271051
rect 379408 271039 379414 271051
rect 378986 271011 379414 271039
rect 378986 270999 378992 271011
rect 379408 270999 379414 271011
rect 379466 270999 379472 271051
rect 379504 270999 379510 271051
rect 379562 271039 379568 271051
rect 379792 271039 379798 271051
rect 379562 271011 379798 271039
rect 379562 270999 379568 271011
rect 379792 270999 379798 271011
rect 379850 270999 379856 271051
rect 379888 270999 379894 271051
rect 379946 271039 379952 271051
rect 380080 271039 380086 271051
rect 379946 271011 380086 271039
rect 379946 270999 379952 271011
rect 380080 270999 380086 271011
rect 380138 270999 380144 271051
rect 380272 270999 380278 271051
rect 380330 271039 380336 271051
rect 380944 271039 380950 271051
rect 380330 271011 380950 271039
rect 380330 270999 380336 271011
rect 380944 270999 380950 271011
rect 381002 270999 381008 271051
rect 381424 270999 381430 271051
rect 381482 271039 381488 271051
rect 388912 271039 388918 271051
rect 381482 271011 388918 271039
rect 381482 270999 381488 271011
rect 388912 270999 388918 271011
rect 388970 270999 388976 271051
rect 381136 270965 381142 270977
rect 358538 270937 378782 270965
rect 378850 270937 381142 270965
rect 358538 270925 358544 270937
rect 221008 270851 221014 270903
rect 221066 270891 221072 270903
rect 249040 270891 249046 270903
rect 221066 270863 249046 270891
rect 221066 270851 221072 270863
rect 249040 270851 249046 270863
rect 249098 270851 249104 270903
rect 253456 270851 253462 270903
rect 253514 270891 253520 270903
rect 259696 270891 259702 270903
rect 253514 270863 259702 270891
rect 253514 270851 253520 270863
rect 259696 270851 259702 270863
rect 259754 270851 259760 270903
rect 260944 270851 260950 270903
rect 261002 270891 261008 270903
rect 277936 270891 277942 270903
rect 261002 270863 277942 270891
rect 261002 270851 261008 270863
rect 277936 270851 277942 270863
rect 277994 270851 278000 270903
rect 279952 270851 279958 270903
rect 280010 270891 280016 270903
rect 284848 270891 284854 270903
rect 280010 270863 284854 270891
rect 280010 270851 280016 270863
rect 284848 270851 284854 270863
rect 284906 270851 284912 270903
rect 296752 270851 296758 270903
rect 296810 270891 296816 270903
rect 378754 270891 378782 270937
rect 381136 270925 381142 270937
rect 381194 270925 381200 270977
rect 381232 270925 381238 270977
rect 381290 270965 381296 270977
rect 390370 270965 390398 271085
rect 381290 270937 390398 270965
rect 390562 270965 390590 271085
rect 390640 271073 390646 271125
rect 390698 271113 390704 271125
rect 409552 271113 409558 271125
rect 390698 271085 409558 271113
rect 390698 271073 390704 271085
rect 409552 271073 409558 271085
rect 409610 271073 409616 271125
rect 410416 271073 410422 271125
rect 410474 271113 410480 271125
rect 416656 271113 416662 271125
rect 410474 271085 416662 271113
rect 410474 271073 410480 271085
rect 416656 271073 416662 271085
rect 416714 271073 416720 271125
rect 398800 270999 398806 271051
rect 398858 271039 398864 271051
rect 516592 271039 516598 271051
rect 398858 271011 516598 271039
rect 398858 270999 398864 271011
rect 516592 270999 516598 271011
rect 516650 270999 516656 271051
rect 527344 270965 527350 270977
rect 390562 270937 527350 270965
rect 381290 270925 381296 270937
rect 527344 270925 527350 270937
rect 527402 270925 527408 270977
rect 382000 270891 382006 270903
rect 296810 270863 378686 270891
rect 378754 270863 382006 270891
rect 296810 270851 296816 270863
rect 257296 270777 257302 270829
rect 257354 270817 257360 270829
rect 277456 270817 277462 270829
rect 257354 270789 277462 270817
rect 257354 270777 257360 270789
rect 277456 270777 277462 270789
rect 277514 270777 277520 270829
rect 317200 270777 317206 270829
rect 317258 270817 317264 270829
rect 327088 270817 327094 270829
rect 317258 270789 327094 270817
rect 317258 270777 317264 270789
rect 327088 270777 327094 270789
rect 327146 270777 327152 270829
rect 327184 270777 327190 270829
rect 327242 270817 327248 270829
rect 372880 270817 372886 270829
rect 327242 270789 372886 270817
rect 327242 270777 327248 270789
rect 372880 270777 372886 270789
rect 372938 270777 372944 270829
rect 372976 270777 372982 270829
rect 373034 270817 373040 270829
rect 377776 270817 377782 270829
rect 373034 270789 377782 270817
rect 373034 270777 373040 270789
rect 377776 270777 377782 270789
rect 377834 270777 377840 270829
rect 378658 270817 378686 270863
rect 382000 270851 382006 270863
rect 382058 270851 382064 270903
rect 383152 270851 383158 270903
rect 383210 270891 383216 270903
rect 383632 270891 383638 270903
rect 383210 270863 383638 270891
rect 383210 270851 383216 270863
rect 383632 270851 383638 270863
rect 383690 270851 383696 270903
rect 385936 270851 385942 270903
rect 385994 270891 386000 270903
rect 390448 270891 390454 270903
rect 385994 270863 390454 270891
rect 385994 270851 386000 270863
rect 390448 270851 390454 270863
rect 390506 270851 390512 270903
rect 390544 270851 390550 270903
rect 390602 270891 390608 270903
rect 406672 270891 406678 270903
rect 390602 270863 406678 270891
rect 390602 270851 390608 270863
rect 406672 270851 406678 270863
rect 406730 270851 406736 270903
rect 406768 270851 406774 270903
rect 406826 270891 406832 270903
rect 543952 270891 543958 270903
rect 406826 270863 543958 270891
rect 406826 270851 406832 270863
rect 543952 270851 543958 270863
rect 544010 270851 544016 270903
rect 392080 270817 392086 270829
rect 378658 270789 392086 270817
rect 392080 270777 392086 270789
rect 392138 270777 392144 270829
rect 394384 270777 394390 270829
rect 394442 270817 394448 270829
rect 402448 270817 402454 270829
rect 394442 270789 402454 270817
rect 394442 270777 394448 270789
rect 402448 270777 402454 270789
rect 402506 270777 402512 270829
rect 402544 270777 402550 270829
rect 402602 270817 402608 270829
rect 536848 270817 536854 270829
rect 402602 270789 536854 270817
rect 402602 270777 402608 270789
rect 536848 270777 536854 270789
rect 536906 270777 536912 270829
rect 358480 270743 358486 270755
rect 217378 270715 358486 270743
rect 358480 270703 358486 270715
rect 358538 270703 358544 270755
rect 364144 270703 364150 270755
rect 364202 270743 364208 270755
rect 369040 270743 369046 270755
rect 364202 270715 369046 270743
rect 364202 270703 364208 270715
rect 369040 270703 369046 270715
rect 369098 270703 369104 270755
rect 373456 270743 373462 270755
rect 369154 270715 373462 270743
rect 207184 270669 207190 270681
rect 206146 270641 207190 270669
rect 207184 270629 207190 270641
rect 207242 270629 207248 270681
rect 231280 270629 231286 270681
rect 231338 270669 231344 270681
rect 328144 270669 328150 270681
rect 231338 270641 328150 270669
rect 231338 270629 231344 270641
rect 328144 270629 328150 270641
rect 328202 270629 328208 270681
rect 328240 270629 328246 270681
rect 328298 270669 328304 270681
rect 338896 270669 338902 270681
rect 328298 270641 338902 270669
rect 328298 270629 328304 270641
rect 338896 270629 338902 270641
rect 338954 270629 338960 270681
rect 341968 270629 341974 270681
rect 342026 270669 342032 270681
rect 369154 270669 369182 270715
rect 373456 270703 373462 270715
rect 373514 270703 373520 270755
rect 374992 270703 374998 270755
rect 375050 270743 375056 270755
rect 375050 270715 381182 270743
rect 375050 270703 375056 270715
rect 342026 270641 369182 270669
rect 342026 270629 342032 270641
rect 369232 270629 369238 270681
rect 369290 270669 369296 270681
rect 380368 270669 380374 270681
rect 369290 270641 380374 270669
rect 369290 270629 369296 270641
rect 380368 270629 380374 270641
rect 380426 270629 380432 270681
rect 381154 270669 381182 270715
rect 381232 270703 381238 270755
rect 381290 270743 381296 270755
rect 383344 270743 383350 270755
rect 381290 270715 383350 270743
rect 381290 270703 381296 270715
rect 383344 270703 383350 270715
rect 383402 270703 383408 270755
rect 383632 270703 383638 270755
rect 383690 270743 383696 270755
rect 387760 270743 387766 270755
rect 383690 270715 387766 270743
rect 383690 270703 383696 270715
rect 387760 270703 387766 270715
rect 387818 270703 387824 270755
rect 389008 270703 389014 270755
rect 389066 270743 389072 270755
rect 411472 270743 411478 270755
rect 389066 270715 411478 270743
rect 389066 270703 389072 270715
rect 411472 270703 411478 270715
rect 411530 270703 411536 270755
rect 414832 270703 414838 270755
rect 414890 270743 414896 270755
rect 434800 270743 434806 270755
rect 414890 270715 434806 270743
rect 414890 270703 414896 270715
rect 434800 270703 434806 270715
rect 434858 270703 434864 270755
rect 385936 270669 385942 270681
rect 381154 270641 385942 270669
rect 385936 270629 385942 270641
rect 385994 270629 386000 270681
rect 386032 270629 386038 270681
rect 386090 270669 386096 270681
rect 565456 270669 565462 270681
rect 386090 270641 565462 270669
rect 386090 270629 386096 270641
rect 565456 270629 565462 270641
rect 565514 270629 565520 270681
rect 245296 270555 245302 270607
rect 245354 270595 245360 270607
rect 445264 270595 445270 270607
rect 245354 270567 445270 270595
rect 245354 270555 245360 270567
rect 445264 270555 445270 270567
rect 445322 270555 445328 270607
rect 231952 270481 231958 270533
rect 232010 270521 232016 270533
rect 328336 270521 328342 270533
rect 232010 270493 328342 270521
rect 232010 270481 232016 270493
rect 328336 270481 328342 270493
rect 328394 270481 328400 270533
rect 331216 270481 331222 270533
rect 331274 270521 331280 270533
rect 338224 270521 338230 270533
rect 331274 270493 338230 270521
rect 331274 270481 331280 270493
rect 338224 270481 338230 270493
rect 338282 270481 338288 270533
rect 338320 270481 338326 270533
rect 338378 270521 338384 270533
rect 348208 270521 348214 270533
rect 338378 270493 348214 270521
rect 338378 270481 338384 270493
rect 348208 270481 348214 270493
rect 348266 270481 348272 270533
rect 348400 270481 348406 270533
rect 348458 270521 348464 270533
rect 362704 270521 362710 270533
rect 348458 270493 362710 270521
rect 348458 270481 348464 270493
rect 362704 270481 362710 270493
rect 362762 270481 362768 270533
rect 365200 270481 365206 270533
rect 365258 270521 365264 270533
rect 368464 270521 368470 270533
rect 365258 270493 368470 270521
rect 365258 270481 365264 270493
rect 368464 270481 368470 270493
rect 368522 270481 368528 270533
rect 378544 270521 378550 270533
rect 368674 270493 378550 270521
rect 245872 270407 245878 270459
rect 245930 270447 245936 270459
rect 368560 270447 368566 270459
rect 245930 270419 368566 270447
rect 245930 270407 245936 270419
rect 368560 270407 368566 270419
rect 368618 270407 368624 270459
rect 232816 270333 232822 270385
rect 232874 270373 232880 270385
rect 328336 270373 328342 270385
rect 232874 270345 328342 270373
rect 232874 270333 232880 270345
rect 328336 270333 328342 270345
rect 328394 270333 328400 270385
rect 328432 270333 328438 270385
rect 328490 270373 328496 270385
rect 334096 270373 334102 270385
rect 328490 270345 334102 270373
rect 328490 270333 328496 270345
rect 334096 270333 334102 270345
rect 334154 270333 334160 270385
rect 352432 270373 352438 270385
rect 336514 270345 352438 270373
rect 233968 270259 233974 270311
rect 234026 270299 234032 270311
rect 336514 270299 336542 270345
rect 352432 270333 352438 270345
rect 352490 270333 352496 270385
rect 353296 270333 353302 270385
rect 353354 270373 353360 270385
rect 368674 270373 368702 270493
rect 378544 270481 378550 270493
rect 378602 270481 378608 270533
rect 378640 270481 378646 270533
rect 378698 270521 378704 270533
rect 394480 270521 394486 270533
rect 378698 270493 394486 270521
rect 378698 270481 378704 270493
rect 394480 270481 394486 270493
rect 394538 270481 394544 270533
rect 394576 270481 394582 270533
rect 394634 270521 394640 270533
rect 403120 270521 403126 270533
rect 394634 270493 403126 270521
rect 394634 270481 394640 270493
rect 403120 270481 403126 270493
rect 403178 270481 403184 270533
rect 427600 270481 427606 270533
rect 427658 270521 427664 270533
rect 437680 270521 437686 270533
rect 427658 270493 437686 270521
rect 427658 270481 427664 270493
rect 437680 270481 437686 270493
rect 437738 270481 437744 270533
rect 368848 270407 368854 270459
rect 368906 270447 368912 270459
rect 452368 270447 452374 270459
rect 368906 270419 452374 270447
rect 368906 270407 368912 270419
rect 452368 270407 452374 270419
rect 452426 270407 452432 270459
rect 552976 270407 552982 270459
rect 553034 270447 553040 270459
rect 573040 270447 573046 270459
rect 553034 270419 573046 270447
rect 553034 270407 553040 270419
rect 573040 270407 573046 270419
rect 573098 270407 573104 270459
rect 590416 270407 590422 270459
rect 590474 270447 590480 270459
rect 600496 270447 600502 270459
rect 590474 270419 600502 270447
rect 590474 270407 590480 270419
rect 600496 270407 600502 270419
rect 600554 270407 600560 270459
rect 388432 270373 388438 270385
rect 353354 270345 368702 270373
rect 368962 270345 388438 270373
rect 353354 270333 353360 270345
rect 234026 270271 336542 270299
rect 234026 270259 234032 270271
rect 336592 270259 336598 270311
rect 336650 270299 336656 270311
rect 343120 270299 343126 270311
rect 336650 270271 343126 270299
rect 336650 270259 336656 270271
rect 343120 270259 343126 270271
rect 343178 270259 343184 270311
rect 359440 270259 359446 270311
rect 359498 270299 359504 270311
rect 368962 270299 368990 270345
rect 388432 270333 388438 270345
rect 388490 270333 388496 270385
rect 388528 270333 388534 270385
rect 388586 270373 388592 270385
rect 579664 270373 579670 270385
rect 388586 270345 579670 270373
rect 388586 270333 388592 270345
rect 579664 270333 579670 270345
rect 579722 270333 579728 270385
rect 359498 270271 368990 270299
rect 359498 270259 359504 270271
rect 369040 270259 369046 270311
rect 369098 270299 369104 270311
rect 383632 270299 383638 270311
rect 369098 270271 383638 270299
rect 369098 270259 369104 270271
rect 383632 270259 383638 270271
rect 383690 270259 383696 270311
rect 383920 270259 383926 270311
rect 383978 270299 383984 270311
rect 586768 270299 586774 270311
rect 383978 270271 586774 270299
rect 383978 270259 383984 270271
rect 586768 270259 586774 270271
rect 586826 270259 586832 270311
rect 247024 270185 247030 270237
rect 247082 270225 247088 270237
rect 348304 270225 348310 270237
rect 247082 270197 348310 270225
rect 247082 270185 247088 270197
rect 348304 270185 348310 270197
rect 348362 270185 348368 270237
rect 459568 270225 459574 270237
rect 349954 270197 459574 270225
rect 234544 270111 234550 270163
rect 234602 270151 234608 270163
rect 323152 270151 323158 270163
rect 234602 270123 323158 270151
rect 234602 270111 234608 270123
rect 323152 270111 323158 270123
rect 323210 270111 323216 270163
rect 323344 270111 323350 270163
rect 323402 270151 323408 270163
rect 336880 270151 336886 270163
rect 323402 270123 336886 270151
rect 323402 270111 323408 270123
rect 336880 270111 336886 270123
rect 336938 270111 336944 270163
rect 342160 270151 342166 270163
rect 336994 270123 342166 270151
rect 235696 270037 235702 270089
rect 235754 270077 235760 270089
rect 336994 270077 337022 270123
rect 342160 270111 342166 270123
rect 342218 270111 342224 270163
rect 235754 270049 337022 270077
rect 235754 270037 235760 270049
rect 341872 270037 341878 270089
rect 341930 270077 341936 270089
rect 348112 270077 348118 270089
rect 341930 270049 348118 270077
rect 341930 270037 341936 270049
rect 348112 270037 348118 270049
rect 348170 270037 348176 270089
rect 348304 270037 348310 270089
rect 348362 270077 348368 270089
rect 349954 270077 349982 270197
rect 459568 270185 459574 270197
rect 459626 270185 459632 270237
rect 355408 270111 355414 270163
rect 355466 270151 355472 270163
rect 364144 270151 364150 270163
rect 355466 270123 364150 270151
rect 355466 270111 355472 270123
rect 364144 270111 364150 270123
rect 364202 270111 364208 270163
rect 364336 270111 364342 270163
rect 364394 270151 364400 270163
rect 378160 270151 378166 270163
rect 364394 270123 378166 270151
rect 364394 270111 364400 270123
rect 378160 270111 378166 270123
rect 378218 270111 378224 270163
rect 380272 270151 380278 270163
rect 378274 270123 380278 270151
rect 348362 270049 349982 270077
rect 348362 270037 348368 270049
rect 355600 270037 355606 270089
rect 355658 270077 355664 270089
rect 370000 270077 370006 270089
rect 355658 270049 370006 270077
rect 355658 270037 355664 270049
rect 370000 270037 370006 270049
rect 370058 270037 370064 270089
rect 370192 270037 370198 270089
rect 370250 270077 370256 270089
rect 374992 270077 374998 270089
rect 370250 270049 374998 270077
rect 370250 270037 370256 270049
rect 374992 270037 374998 270049
rect 375050 270037 375056 270089
rect 375088 270037 375094 270089
rect 375146 270077 375152 270089
rect 378274 270077 378302 270123
rect 380272 270111 380278 270123
rect 380330 270111 380336 270163
rect 380368 270111 380374 270163
rect 380426 270151 380432 270163
rect 381040 270151 381046 270163
rect 380426 270123 381046 270151
rect 380426 270111 380432 270123
rect 381040 270111 381046 270123
rect 381098 270111 381104 270163
rect 381136 270111 381142 270163
rect 381194 270151 381200 270163
rect 593968 270151 593974 270163
rect 381194 270123 593974 270151
rect 381194 270111 381200 270123
rect 593968 270111 593974 270123
rect 594026 270111 594032 270163
rect 375146 270049 378302 270077
rect 375146 270037 375152 270049
rect 378544 270037 378550 270089
rect 378602 270077 378608 270089
rect 380080 270077 380086 270089
rect 378602 270049 380086 270077
rect 378602 270037 378608 270049
rect 380080 270037 380086 270049
rect 380138 270037 380144 270089
rect 380464 270037 380470 270089
rect 380522 270077 380528 270089
rect 380848 270077 380854 270089
rect 380522 270049 380854 270077
rect 380522 270037 380528 270049
rect 380848 270037 380854 270049
rect 380906 270037 380912 270089
rect 380944 270037 380950 270089
rect 381002 270077 381008 270089
rect 427600 270077 427606 270089
rect 381002 270049 427606 270077
rect 381002 270037 381008 270049
rect 427600 270037 427606 270049
rect 427658 270037 427664 270089
rect 437314 270049 437630 270077
rect 159856 269963 159862 270015
rect 159914 270003 159920 270015
rect 161104 270003 161110 270015
rect 159914 269975 161110 270003
rect 159914 269963 159920 269975
rect 161104 269963 161110 269975
rect 161162 269963 161168 270015
rect 247600 269963 247606 270015
rect 247658 270003 247664 270015
rect 437314 270003 437342 270049
rect 247658 269975 437342 270003
rect 437602 270003 437630 270049
rect 437680 270037 437686 270089
rect 437738 270077 437744 270089
rect 597520 270077 597526 270089
rect 437738 270049 597526 270077
rect 437738 270037 437744 270049
rect 597520 270037 597526 270049
rect 597578 270037 597584 270089
rect 466576 270003 466582 270015
rect 437602 269975 466582 270003
rect 247658 269963 247664 269975
rect 466576 269963 466582 269975
rect 466634 269963 466640 270015
rect 573136 269963 573142 270015
rect 573194 270003 573200 270015
rect 589168 270003 589174 270015
rect 573194 269975 589174 270003
rect 573194 269963 573200 269975
rect 589168 269963 589174 269975
rect 589226 269963 589232 270015
rect 216016 269889 216022 269941
rect 216074 269929 216080 269941
rect 243280 269929 243286 269941
rect 216074 269901 243286 269929
rect 216074 269889 216080 269901
rect 243280 269889 243286 269901
rect 243338 269889 243344 269941
rect 248560 269889 248566 269941
rect 248618 269929 248624 269941
rect 427600 269929 427606 269941
rect 248618 269901 342302 269929
rect 248618 269889 248624 269901
rect 226960 269815 226966 269867
rect 227018 269855 227024 269867
rect 295408 269855 295414 269867
rect 227018 269827 295414 269855
rect 227018 269815 227024 269827
rect 295408 269815 295414 269827
rect 295466 269815 295472 269867
rect 295504 269815 295510 269867
rect 295562 269855 295568 269867
rect 302512 269855 302518 269867
rect 295562 269827 302518 269855
rect 295562 269815 295568 269827
rect 302512 269815 302518 269827
rect 302570 269815 302576 269867
rect 308176 269815 308182 269867
rect 308234 269855 308240 269867
rect 311920 269855 311926 269867
rect 308234 269827 311926 269855
rect 308234 269815 308240 269827
rect 311920 269815 311926 269827
rect 311978 269815 311984 269867
rect 312016 269815 312022 269867
rect 312074 269855 312080 269867
rect 316336 269855 316342 269867
rect 312074 269827 316342 269855
rect 312074 269815 312080 269827
rect 316336 269815 316342 269827
rect 316394 269815 316400 269867
rect 316432 269815 316438 269867
rect 316490 269855 316496 269867
rect 327856 269855 327862 269867
rect 316490 269827 327862 269855
rect 316490 269815 316496 269827
rect 327856 269815 327862 269827
rect 327914 269815 327920 269867
rect 327952 269815 327958 269867
rect 328010 269855 328016 269867
rect 338320 269855 338326 269867
rect 328010 269827 338326 269855
rect 328010 269815 328016 269827
rect 338320 269815 338326 269827
rect 338378 269815 338384 269867
rect 342160 269815 342166 269867
rect 342218 269815 342224 269867
rect 342274 269855 342302 269901
rect 342562 269901 427606 269929
rect 342562 269855 342590 269901
rect 427600 269889 427606 269901
rect 427658 269889 427664 269941
rect 437584 269889 437590 269941
rect 437642 269929 437648 269941
rect 473776 269929 473782 269941
rect 437642 269901 473782 269929
rect 437642 269889 437648 269901
rect 473776 269889 473782 269901
rect 473834 269889 473840 269941
rect 342274 269827 342590 269855
rect 348208 269815 348214 269867
rect 348266 269855 348272 269867
rect 437104 269855 437110 269867
rect 348266 269827 437110 269855
rect 348266 269815 348272 269827
rect 437104 269815 437110 269827
rect 437162 269815 437168 269867
rect 437488 269815 437494 269867
rect 437546 269855 437552 269867
rect 539248 269855 539254 269867
rect 437546 269827 539254 269855
rect 437546 269815 437552 269827
rect 539248 269815 539254 269827
rect 539306 269815 539312 269867
rect 249616 269741 249622 269793
rect 249674 269781 249680 269793
rect 342178 269781 342206 269815
rect 342544 269781 342550 269793
rect 249674 269753 342110 269781
rect 342178 269753 342550 269781
rect 249674 269741 249680 269753
rect 250288 269667 250294 269719
rect 250346 269707 250352 269719
rect 341872 269707 341878 269719
rect 250346 269679 341878 269707
rect 250346 269667 250352 269679
rect 341872 269667 341878 269679
rect 341930 269667 341936 269719
rect 342082 269707 342110 269753
rect 342544 269741 342550 269753
rect 342602 269741 342608 269793
rect 481072 269781 481078 269793
rect 342658 269753 481078 269781
rect 342658 269707 342686 269753
rect 481072 269741 481078 269753
rect 481130 269741 481136 269793
rect 483952 269741 483958 269793
rect 484010 269781 484016 269793
rect 518320 269781 518326 269793
rect 484010 269753 518326 269781
rect 484010 269741 484016 269753
rect 518320 269741 518326 269753
rect 518378 269741 518384 269793
rect 342082 269679 342686 269707
rect 348112 269667 348118 269719
rect 348170 269707 348176 269719
rect 365200 269707 365206 269719
rect 348170 269679 365206 269707
rect 348170 269667 348176 269679
rect 365200 269667 365206 269679
rect 365258 269667 365264 269719
rect 365296 269667 365302 269719
rect 365354 269707 365360 269719
rect 379696 269707 379702 269719
rect 365354 269679 379702 269707
rect 365354 269667 365360 269679
rect 379696 269667 379702 269679
rect 379754 269667 379760 269719
rect 379792 269667 379798 269719
rect 379850 269707 379856 269719
rect 437968 269707 437974 269719
rect 379850 269679 437974 269707
rect 379850 269667 379856 269679
rect 437968 269667 437974 269679
rect 438026 269667 438032 269719
rect 438160 269667 438166 269719
rect 438218 269707 438224 269719
rect 488080 269707 488086 269719
rect 438218 269679 488086 269707
rect 438218 269667 438224 269679
rect 488080 269667 488086 269679
rect 488138 269667 488144 269719
rect 251344 269593 251350 269645
rect 251402 269633 251408 269645
rect 336208 269633 336214 269645
rect 251402 269605 336214 269633
rect 251402 269593 251408 269605
rect 336208 269593 336214 269605
rect 336266 269593 336272 269645
rect 342832 269593 342838 269645
rect 342890 269633 342896 269645
rect 437392 269633 437398 269645
rect 342890 269605 437398 269633
rect 342890 269593 342896 269605
rect 437392 269593 437398 269605
rect 437450 269593 437456 269645
rect 437584 269593 437590 269645
rect 437642 269633 437648 269645
rect 437776 269633 437782 269645
rect 437642 269605 437782 269633
rect 437642 269593 437648 269605
rect 437776 269593 437782 269605
rect 437834 269593 437840 269645
rect 437872 269593 437878 269645
rect 437930 269633 437936 269645
rect 495184 269633 495190 269645
rect 437930 269605 495190 269633
rect 437930 269593 437936 269605
rect 495184 269593 495190 269605
rect 495242 269593 495248 269645
rect 509872 269633 509878 269645
rect 502402 269605 509878 269633
rect 85264 269519 85270 269571
rect 85322 269559 85328 269571
rect 86512 269559 86518 269571
rect 85322 269531 86518 269559
rect 85322 269519 85328 269531
rect 86512 269519 86518 269531
rect 86570 269519 86576 269571
rect 227536 269519 227542 269571
rect 227594 269559 227600 269571
rect 295504 269559 295510 269571
rect 227594 269531 295510 269559
rect 227594 269519 227600 269531
rect 295504 269519 295510 269531
rect 295562 269519 295568 269571
rect 297904 269519 297910 269571
rect 297962 269559 297968 269571
rect 308176 269559 308182 269571
rect 297962 269531 308182 269559
rect 297962 269519 297968 269531
rect 308176 269519 308182 269531
rect 308234 269519 308240 269571
rect 308272 269519 308278 269571
rect 308330 269559 308336 269571
rect 316816 269559 316822 269571
rect 308330 269531 316822 269559
rect 308330 269519 308336 269531
rect 316816 269519 316822 269531
rect 316874 269519 316880 269571
rect 318160 269519 318166 269571
rect 318218 269559 318224 269571
rect 326800 269559 326806 269571
rect 318218 269531 326806 269559
rect 318218 269519 318224 269531
rect 326800 269519 326806 269531
rect 326858 269519 326864 269571
rect 328048 269519 328054 269571
rect 328106 269559 328112 269571
rect 417712 269559 417718 269571
rect 328106 269531 342110 269559
rect 328106 269519 328112 269531
rect 236272 269445 236278 269497
rect 236330 269485 236336 269497
rect 341968 269485 341974 269497
rect 236330 269457 341974 269485
rect 236330 269445 236336 269457
rect 341968 269445 341974 269457
rect 342026 269445 342032 269497
rect 342082 269485 342110 269531
rect 342754 269531 417718 269559
rect 342754 269485 342782 269531
rect 417712 269519 417718 269531
rect 417770 269519 417776 269571
rect 437680 269519 437686 269571
rect 437738 269559 437744 269571
rect 458224 269559 458230 269571
rect 437738 269531 458230 269559
rect 437738 269519 437744 269531
rect 458224 269519 458230 269531
rect 458282 269519 458288 269571
rect 478000 269519 478006 269571
rect 478058 269559 478064 269571
rect 501040 269559 501046 269571
rect 478058 269531 501046 269559
rect 478058 269519 478064 269531
rect 501040 269519 501046 269531
rect 501098 269519 501104 269571
rect 501136 269519 501142 269571
rect 501194 269559 501200 269571
rect 502402 269559 502430 269605
rect 509872 269593 509878 269605
rect 509930 269593 509936 269645
rect 532834 269605 555806 269633
rect 501194 269531 502430 269559
rect 501194 269519 501200 269531
rect 529840 269519 529846 269571
rect 529898 269559 529904 269571
rect 532834 269559 532862 269605
rect 529898 269531 532862 269559
rect 555778 269559 555806 269605
rect 560656 269559 560662 269571
rect 555778 269531 560662 269559
rect 529898 269519 529904 269531
rect 560656 269519 560662 269531
rect 560714 269519 560720 269571
rect 573136 269519 573142 269571
rect 573194 269559 573200 269571
rect 593200 269559 593206 269571
rect 573194 269531 593206 269559
rect 573194 269519 573200 269531
rect 593200 269519 593206 269531
rect 593258 269519 593264 269571
rect 342082 269457 342782 269485
rect 360976 269445 360982 269497
rect 361034 269485 361040 269497
rect 378544 269485 378550 269497
rect 361034 269457 378550 269485
rect 361034 269445 361040 269457
rect 378544 269445 378550 269457
rect 378602 269445 378608 269497
rect 378640 269445 378646 269497
rect 378698 269485 378704 269497
rect 393136 269485 393142 269497
rect 378698 269457 393142 269485
rect 378698 269445 378704 269457
rect 393136 269445 393142 269457
rect 393194 269445 393200 269497
rect 398800 269445 398806 269497
rect 398858 269485 398864 269497
rect 437488 269485 437494 269497
rect 398858 269457 437494 269485
rect 398858 269445 398864 269457
rect 437488 269445 437494 269457
rect 437546 269445 437552 269497
rect 437584 269445 437590 269497
rect 437642 269485 437648 269497
rect 457936 269485 457942 269497
rect 437642 269457 457942 269485
rect 437642 269445 437648 269457
rect 457936 269445 457942 269457
rect 457994 269445 458000 269497
rect 458608 269445 458614 269497
rect 458666 269485 458672 269497
rect 532816 269485 532822 269497
rect 458666 269457 532822 269485
rect 458666 269445 458672 269457
rect 532816 269445 532822 269457
rect 532874 269445 532880 269497
rect 533104 269445 533110 269497
rect 533162 269485 533168 269497
rect 626032 269485 626038 269497
rect 533162 269457 626038 269485
rect 533162 269445 533168 269457
rect 626032 269445 626038 269457
rect 626090 269445 626096 269497
rect 228496 269371 228502 269423
rect 228554 269411 228560 269423
rect 228554 269383 298046 269411
rect 228554 269371 228560 269383
rect 229552 269297 229558 269349
rect 229610 269337 229616 269349
rect 297904 269337 297910 269349
rect 229610 269309 297910 269337
rect 229610 269297 229616 269309
rect 297904 269297 297910 269309
rect 297962 269297 297968 269349
rect 298018 269337 298046 269383
rect 304912 269371 304918 269423
rect 304970 269411 304976 269423
rect 327952 269411 327958 269423
rect 304970 269383 327958 269411
rect 304970 269371 304976 269383
rect 327952 269371 327958 269383
rect 328010 269371 328016 269423
rect 328432 269371 328438 269423
rect 328490 269411 328496 269423
rect 437296 269411 437302 269423
rect 328490 269383 437302 269411
rect 328490 269371 328496 269383
rect 437296 269371 437302 269383
rect 437354 269371 437360 269423
rect 437392 269371 437398 269423
rect 437450 269411 437456 269423
rect 437776 269411 437782 269423
rect 437450 269383 437782 269411
rect 437450 269371 437456 269383
rect 437776 269371 437782 269383
rect 437834 269371 437840 269423
rect 437986 269383 438206 269411
rect 309712 269337 309718 269349
rect 298018 269309 309718 269337
rect 309712 269297 309718 269309
rect 309770 269297 309776 269349
rect 311920 269297 311926 269349
rect 311978 269337 311984 269349
rect 316048 269337 316054 269349
rect 311978 269309 316054 269337
rect 311978 269297 311984 269309
rect 316048 269297 316054 269309
rect 316106 269297 316112 269349
rect 316144 269297 316150 269349
rect 316202 269337 316208 269349
rect 327568 269337 327574 269349
rect 316202 269309 327574 269337
rect 316202 269297 316208 269309
rect 327568 269297 327574 269309
rect 327626 269297 327632 269349
rect 327856 269297 327862 269349
rect 327914 269337 327920 269349
rect 437986 269337 438014 269383
rect 327914 269309 438014 269337
rect 438178 269337 438206 269383
rect 438256 269371 438262 269423
rect 438314 269411 438320 269423
rect 567760 269411 567766 269423
rect 438314 269383 567766 269411
rect 438314 269371 438320 269383
rect 567760 269371 567766 269383
rect 567818 269371 567824 269423
rect 574864 269337 574870 269349
rect 438178 269309 458174 269337
rect 327914 269297 327920 269309
rect 53872 269223 53878 269275
rect 53930 269263 53936 269275
rect 205936 269263 205942 269275
rect 53930 269235 205942 269263
rect 53930 269223 53936 269235
rect 205936 269223 205942 269235
rect 205994 269223 206000 269275
rect 221488 269223 221494 269275
rect 221546 269263 221552 269275
rect 252496 269263 252502 269275
rect 221546 269235 252502 269263
rect 221546 269223 221552 269235
rect 252496 269223 252502 269235
rect 252554 269223 252560 269275
rect 254128 269223 254134 269275
rect 254186 269263 254192 269275
rect 342064 269263 342070 269275
rect 254186 269235 342070 269263
rect 254186 269223 254192 269235
rect 342064 269223 342070 269235
rect 342122 269223 342128 269275
rect 342448 269223 342454 269275
rect 342506 269263 342512 269275
rect 380176 269263 380182 269275
rect 342506 269235 380182 269263
rect 342506 269223 342512 269235
rect 380176 269223 380182 269235
rect 380234 269223 380240 269275
rect 380290 269235 381470 269263
rect 244144 269149 244150 269201
rect 244202 269189 244208 269201
rect 341968 269189 341974 269201
rect 244202 269161 341974 269189
rect 244202 269149 244208 269161
rect 341968 269149 341974 269161
rect 342026 269149 342032 269201
rect 342544 269149 342550 269201
rect 342602 269189 342608 269201
rect 380290 269189 380318 269235
rect 381442 269189 381470 269235
rect 381616 269223 381622 269275
rect 381674 269263 381680 269275
rect 458146 269263 458174 269309
rect 458530 269309 574870 269337
rect 458530 269263 458558 269309
rect 574864 269297 574870 269309
rect 574922 269297 574928 269349
rect 381674 269235 457982 269263
rect 458146 269235 458558 269263
rect 381674 269223 381680 269235
rect 457954 269201 457982 269235
rect 467920 269223 467926 269275
rect 467978 269263 467984 269275
rect 520144 269263 520150 269275
rect 467978 269235 520150 269263
rect 467978 269223 467984 269235
rect 520144 269223 520150 269235
rect 520202 269223 520208 269275
rect 632080 269223 632086 269275
rect 632138 269263 632144 269275
rect 649360 269263 649366 269275
rect 632138 269235 649366 269263
rect 632138 269223 632144 269235
rect 649360 269223 649366 269235
rect 649418 269223 649424 269275
rect 438352 269189 438358 269201
rect 342602 269161 380318 269189
rect 380386 269161 381374 269189
rect 381442 269161 438358 269189
rect 342602 269149 342608 269161
rect 203824 269075 203830 269127
rect 203882 269115 203888 269127
rect 270928 269115 270934 269127
rect 203882 269087 270934 269115
rect 203882 269075 203888 269087
rect 270928 269075 270934 269087
rect 270986 269075 270992 269127
rect 272752 269075 272758 269127
rect 272810 269115 272816 269127
rect 316144 269115 316150 269127
rect 272810 269087 316150 269115
rect 272810 269075 272816 269087
rect 316144 269075 316150 269087
rect 316202 269075 316208 269127
rect 316240 269075 316246 269127
rect 316298 269115 316304 269127
rect 336112 269115 336118 269127
rect 316298 269087 336118 269115
rect 316298 269075 316304 269087
rect 336112 269075 336118 269087
rect 336170 269075 336176 269127
rect 336208 269075 336214 269127
rect 336266 269115 336272 269127
rect 342640 269115 342646 269127
rect 336266 269087 342646 269115
rect 336266 269075 336272 269087
rect 342640 269075 342646 269087
rect 342698 269075 342704 269127
rect 342736 269075 342742 269127
rect 342794 269115 342800 269127
rect 366736 269115 366742 269127
rect 342794 269087 366742 269115
rect 342794 269075 342800 269087
rect 366736 269075 366742 269087
rect 366794 269075 366800 269127
rect 367312 269075 367318 269127
rect 367370 269115 367376 269127
rect 378640 269115 378646 269127
rect 367370 269087 378646 269115
rect 367370 269075 367376 269087
rect 378640 269075 378646 269087
rect 378698 269075 378704 269127
rect 378736 269075 378742 269127
rect 378794 269115 378800 269127
rect 380386 269115 380414 269161
rect 381346 269115 381374 269161
rect 438352 269149 438358 269161
rect 438410 269149 438416 269201
rect 457936 269149 457942 269201
rect 457994 269149 458000 269201
rect 509872 269149 509878 269201
rect 509930 269189 509936 269201
rect 529840 269189 529846 269201
rect 509930 269161 529846 269189
rect 509930 269149 509936 269161
rect 529840 269149 529846 269161
rect 529898 269149 529904 269201
rect 558256 269115 558262 269127
rect 378794 269087 380414 269115
rect 380482 269087 381278 269115
rect 381346 269087 558262 269115
rect 378794 269075 378800 269087
rect 243280 269001 243286 269053
rect 243338 269041 243344 269053
rect 380482 269041 380510 269087
rect 381250 269041 381278 269087
rect 558256 269075 558262 269087
rect 558314 269075 558320 269127
rect 431056 269041 431062 269053
rect 243338 269013 380510 269041
rect 380578 269013 381182 269041
rect 381250 269013 431062 269041
rect 243338 269001 243344 269013
rect 242608 268927 242614 268979
rect 242666 268967 242672 268979
rect 380578 268967 380606 269013
rect 381154 268967 381182 269013
rect 431056 269001 431062 269013
rect 431114 269001 431120 269053
rect 458032 269001 458038 269053
rect 458090 269041 458096 269053
rect 467920 269041 467926 269053
rect 458090 269013 467926 269041
rect 458090 269001 458096 269013
rect 467920 269001 467926 269013
rect 467978 269001 467984 269053
rect 423856 268967 423862 268979
rect 242666 268939 380606 268967
rect 380674 268939 381086 268967
rect 381154 268939 423862 268967
rect 242666 268927 242672 268939
rect 237136 268853 237142 268905
rect 237194 268893 237200 268905
rect 355408 268893 355414 268905
rect 237194 268865 355414 268893
rect 237194 268853 237200 268865
rect 355408 268853 355414 268865
rect 355466 268853 355472 268905
rect 355504 268853 355510 268905
rect 355562 268893 355568 268905
rect 360880 268893 360886 268905
rect 355562 268865 360886 268893
rect 355562 268853 355568 268865
rect 360880 268853 360886 268865
rect 360938 268853 360944 268905
rect 362704 268853 362710 268905
rect 362762 268893 362768 268905
rect 377584 268893 377590 268905
rect 362762 268865 377590 268893
rect 362762 268853 362768 268865
rect 377584 268853 377590 268865
rect 377642 268853 377648 268905
rect 378352 268853 378358 268905
rect 378410 268893 378416 268905
rect 380674 268893 380702 268939
rect 378410 268865 380702 268893
rect 381058 268893 381086 268939
rect 423856 268927 423862 268939
rect 423914 268927 423920 268979
rect 458512 268927 458518 268979
rect 458570 268967 458576 268979
rect 478000 268967 478006 268979
rect 458570 268939 478006 268967
rect 458570 268927 458576 268939
rect 478000 268927 478006 268939
rect 478058 268927 478064 268979
rect 541378 268939 550142 268967
rect 398800 268893 398806 268905
rect 381058 268865 398806 268893
rect 378410 268853 378416 268865
rect 398800 268853 398806 268865
rect 398858 268853 398864 268905
rect 417712 268853 417718 268905
rect 417770 268893 417776 268905
rect 437680 268893 437686 268905
rect 417770 268865 437686 268893
rect 417770 268853 417776 268865
rect 437680 268853 437686 268865
rect 437738 268853 437744 268905
rect 442594 268865 467966 268893
rect 241552 268779 241558 268831
rect 241610 268819 241616 268831
rect 380176 268819 380182 268831
rect 241610 268791 380182 268819
rect 241610 268779 241616 268791
rect 380176 268779 380182 268791
rect 380234 268779 380240 268831
rect 380848 268819 380854 268831
rect 380578 268791 380854 268819
rect 240880 268705 240886 268757
rect 240938 268745 240944 268757
rect 380578 268745 380606 268791
rect 380848 268779 380854 268791
rect 380906 268779 380912 268831
rect 410416 268819 410422 268831
rect 381058 268791 398846 268819
rect 381058 268745 381086 268791
rect 390640 268745 390646 268757
rect 240938 268717 380606 268745
rect 380674 268717 381086 268745
rect 381154 268717 390646 268745
rect 240938 268705 240944 268717
rect 238288 268631 238294 268683
rect 238346 268671 238352 268683
rect 379888 268671 379894 268683
rect 238346 268643 379894 268671
rect 238346 268631 238352 268643
rect 379888 268631 379894 268643
rect 379946 268631 379952 268683
rect 380176 268631 380182 268683
rect 380234 268671 380240 268683
rect 380674 268671 380702 268717
rect 380234 268643 380702 268671
rect 380234 268631 380240 268643
rect 380848 268631 380854 268683
rect 380906 268671 380912 268683
rect 381154 268671 381182 268717
rect 390640 268705 390646 268717
rect 390698 268705 390704 268757
rect 398818 268745 398846 268791
rect 399010 268791 410422 268819
rect 399010 268745 399038 268791
rect 410416 268779 410422 268791
rect 410474 268779 410480 268831
rect 442594 268819 442622 268865
rect 427714 268791 442622 268819
rect 398818 268717 399038 268745
rect 413218 268717 423230 268745
rect 380906 268643 381182 268671
rect 380906 268631 380912 268643
rect 381232 268631 381238 268683
rect 381290 268671 381296 268683
rect 413218 268671 413246 268717
rect 381290 268643 413246 268671
rect 423202 268671 423230 268717
rect 427714 268671 427742 268791
rect 467938 268745 467966 268865
rect 483952 268853 483958 268905
rect 484010 268893 484016 268905
rect 484010 268865 511166 268893
rect 484010 268853 484016 268865
rect 483856 268819 483862 268831
rect 469570 268791 483862 268819
rect 469570 268745 469598 268791
rect 483856 268779 483862 268791
rect 483914 268779 483920 268831
rect 511138 268819 511166 268865
rect 541378 268819 541406 268939
rect 511138 268791 541406 268819
rect 550114 268819 550142 268939
rect 560080 268819 560086 268831
rect 550114 268791 560086 268819
rect 560080 268779 560086 268791
rect 560138 268779 560144 268831
rect 467938 268717 469598 268745
rect 423202 268643 427742 268671
rect 381290 268631 381296 268643
rect 238864 268557 238870 268609
rect 238922 268597 238928 268609
rect 368656 268597 368662 268609
rect 238922 268569 368662 268597
rect 238922 268557 238928 268569
rect 368656 268557 368662 268569
rect 368714 268557 368720 268609
rect 370192 268597 370198 268609
rect 368770 268569 370198 268597
rect 240016 268483 240022 268535
rect 240074 268523 240080 268535
rect 368770 268523 368798 268569
rect 370192 268557 370198 268569
rect 370250 268557 370256 268609
rect 370288 268557 370294 268609
rect 370346 268597 370352 268609
rect 378736 268597 378742 268609
rect 370346 268569 378742 268597
rect 370346 268557 370352 268569
rect 378736 268557 378742 268569
rect 378794 268557 378800 268609
rect 378832 268557 378838 268609
rect 378890 268597 378896 268609
rect 380272 268597 380278 268609
rect 378890 268569 380278 268597
rect 378890 268557 378896 268569
rect 380272 268557 380278 268569
rect 380330 268557 380336 268609
rect 380560 268557 380566 268609
rect 380618 268597 380624 268609
rect 388528 268597 388534 268609
rect 380618 268569 388534 268597
rect 380618 268557 380624 268569
rect 388528 268557 388534 268569
rect 388586 268557 388592 268609
rect 388816 268557 388822 268609
rect 388874 268597 388880 268609
rect 389392 268597 389398 268609
rect 388874 268569 389398 268597
rect 388874 268557 388880 268569
rect 389392 268557 389398 268569
rect 389450 268557 389456 268609
rect 389488 268557 389494 268609
rect 389546 268597 389552 268609
rect 400720 268597 400726 268609
rect 389546 268569 400726 268597
rect 389546 268557 389552 268569
rect 400720 268557 400726 268569
rect 400778 268557 400784 268609
rect 240074 268495 368798 268523
rect 240074 268483 240080 268495
rect 368848 268483 368854 268535
rect 368906 268523 368912 268535
rect 387664 268523 387670 268535
rect 368906 268495 387670 268523
rect 368906 268483 368912 268495
rect 387664 268483 387670 268495
rect 387722 268483 387728 268535
rect 387760 268483 387766 268535
rect 387818 268523 387824 268535
rect 397360 268523 397366 268535
rect 387818 268495 397366 268523
rect 387818 268483 387824 268495
rect 397360 268483 397366 268495
rect 397418 268483 397424 268535
rect 225808 268409 225814 268461
rect 225866 268449 225872 268461
rect 288208 268449 288214 268461
rect 225866 268421 288214 268449
rect 225866 268409 225872 268421
rect 288208 268409 288214 268421
rect 288266 268409 288272 268461
rect 294256 268409 294262 268461
rect 294314 268449 294320 268461
rect 294314 268421 316766 268449
rect 294314 268409 294320 268421
rect 210928 268335 210934 268387
rect 210986 268375 210992 268387
rect 271984 268375 271990 268387
rect 210986 268347 271990 268375
rect 210986 268335 210992 268347
rect 271984 268335 271990 268347
rect 272042 268335 272048 268387
rect 284848 268335 284854 268387
rect 284906 268375 284912 268387
rect 316240 268375 316246 268387
rect 284906 268347 316246 268375
rect 284906 268335 284912 268347
rect 316240 268335 316246 268347
rect 316298 268335 316304 268387
rect 316738 268375 316766 268421
rect 321904 268409 321910 268461
rect 321962 268449 321968 268461
rect 324592 268449 324598 268461
rect 321962 268421 324598 268449
rect 321962 268409 321968 268421
rect 324592 268409 324598 268421
rect 324650 268409 324656 268461
rect 324688 268409 324694 268461
rect 324746 268449 324752 268461
rect 338032 268449 338038 268461
rect 324746 268421 338038 268449
rect 324746 268409 324752 268421
rect 338032 268409 338038 268421
rect 338090 268409 338096 268461
rect 357040 268409 357046 268461
rect 357098 268449 357104 268461
rect 451120 268449 451126 268461
rect 357098 268421 451126 268449
rect 357098 268409 357104 268421
rect 451120 268409 451126 268421
rect 451178 268409 451184 268461
rect 337840 268375 337846 268387
rect 316738 268347 337846 268375
rect 337840 268335 337846 268347
rect 337898 268335 337904 268387
rect 357616 268335 357622 268387
rect 357674 268375 357680 268387
rect 357674 268347 360350 268375
rect 357674 268335 357680 268347
rect 218032 268261 218038 268313
rect 218090 268301 218096 268313
rect 272656 268301 272662 268313
rect 218090 268273 272662 268301
rect 218090 268261 218096 268273
rect 272656 268261 272662 268273
rect 272714 268261 272720 268313
rect 287056 268261 287062 268313
rect 287114 268301 287120 268313
rect 312016 268301 312022 268313
rect 287114 268273 312022 268301
rect 287114 268261 287120 268273
rect 312016 268261 312022 268273
rect 312074 268261 312080 268313
rect 312208 268261 312214 268313
rect 312266 268301 312272 268313
rect 330064 268301 330070 268313
rect 312266 268273 330070 268301
rect 312266 268261 312272 268273
rect 330064 268261 330070 268273
rect 330122 268261 330128 268313
rect 333424 268261 333430 268313
rect 333482 268301 333488 268313
rect 342640 268301 342646 268313
rect 333482 268273 342646 268301
rect 333482 268261 333488 268273
rect 342640 268261 342646 268273
rect 342698 268261 342704 268313
rect 355408 268261 355414 268313
rect 355466 268301 355472 268313
rect 360112 268301 360118 268313
rect 355466 268273 360118 268301
rect 355466 268261 355472 268273
rect 360112 268261 360118 268273
rect 360170 268261 360176 268313
rect 223696 268187 223702 268239
rect 223754 268227 223760 268239
rect 270352 268227 270358 268239
rect 223754 268199 270358 268227
rect 223754 268187 223760 268199
rect 270352 268187 270358 268199
rect 270410 268187 270416 268239
rect 285040 268187 285046 268239
rect 285098 268227 285104 268239
rect 312880 268227 312886 268239
rect 285098 268199 312886 268227
rect 285098 268187 285104 268199
rect 312880 268187 312886 268199
rect 312938 268187 312944 268239
rect 314800 268187 314806 268239
rect 314858 268227 314864 268239
rect 322480 268227 322486 268239
rect 314858 268199 322486 268227
rect 314858 268187 314864 268199
rect 322480 268187 322486 268199
rect 322538 268187 322544 268239
rect 322768 268187 322774 268239
rect 322826 268227 322832 268239
rect 326704 268227 326710 268239
rect 322826 268199 326710 268227
rect 322826 268187 322832 268199
rect 326704 268187 326710 268199
rect 326762 268187 326768 268239
rect 326800 268187 326806 268239
rect 326858 268227 326864 268239
rect 355600 268227 355606 268239
rect 326858 268199 355606 268227
rect 326858 268187 326864 268199
rect 355600 268187 355606 268199
rect 355658 268187 355664 268239
rect 355888 268187 355894 268239
rect 355946 268227 355952 268239
rect 360208 268227 360214 268239
rect 355946 268199 360214 268227
rect 355946 268187 355952 268199
rect 360208 268187 360214 268199
rect 360266 268187 360272 268239
rect 360322 268227 360350 268347
rect 360880 268335 360886 268387
rect 360938 268375 360944 268387
rect 436912 268375 436918 268387
rect 360938 268347 436918 268375
rect 360938 268335 360944 268347
rect 436912 268335 436918 268347
rect 436970 268335 436976 268387
rect 360400 268261 360406 268313
rect 360458 268301 360464 268313
rect 380368 268301 380374 268313
rect 360458 268273 380374 268301
rect 360458 268261 360464 268273
rect 380368 268261 380374 268273
rect 380426 268261 380432 268313
rect 380464 268261 380470 268313
rect 380522 268301 380528 268313
rect 419056 268301 419062 268313
rect 380522 268273 419062 268301
rect 380522 268261 380528 268273
rect 419056 268261 419062 268273
rect 419114 268261 419120 268313
rect 377104 268227 377110 268239
rect 360322 268199 377110 268227
rect 377104 268187 377110 268199
rect 377162 268187 377168 268239
rect 378640 268187 378646 268239
rect 378698 268227 378704 268239
rect 378698 268199 388382 268227
rect 378698 268187 378704 268199
rect 223216 268113 223222 268165
rect 223274 268153 223280 268165
rect 266512 268153 266518 268165
rect 223274 268125 266518 268153
rect 223274 268113 223280 268125
rect 266512 268113 266518 268125
rect 266570 268113 266576 268165
rect 286000 268113 286006 268165
rect 286058 268153 286064 268165
rect 315760 268153 315766 268165
rect 286058 268125 315766 268153
rect 286058 268113 286064 268125
rect 315760 268113 315766 268125
rect 315818 268113 315824 268165
rect 315856 268113 315862 268165
rect 315914 268153 315920 268165
rect 317872 268153 317878 268165
rect 315914 268125 317878 268153
rect 315914 268113 315920 268125
rect 317872 268113 317878 268125
rect 317930 268113 317936 268165
rect 322192 268153 322198 268165
rect 317986 268125 322198 268153
rect 235888 268039 235894 268091
rect 235946 268079 235952 268091
rect 274864 268079 274870 268091
rect 235946 268051 253598 268079
rect 235946 268039 235952 268051
rect 222544 267965 222550 268017
rect 222602 268005 222608 268017
rect 253456 268005 253462 268017
rect 222602 267977 253462 268005
rect 222602 267965 222608 267977
rect 253456 267965 253462 267977
rect 253514 267965 253520 268017
rect 253570 268005 253598 268051
rect 253762 268051 274870 268079
rect 253762 268005 253790 268051
rect 274864 268039 274870 268051
rect 274922 268039 274928 268091
rect 310960 268039 310966 268091
rect 311018 268079 311024 268091
rect 317680 268079 317686 268091
rect 311018 268051 317686 268079
rect 311018 268039 311024 268051
rect 317680 268039 317686 268051
rect 317738 268039 317744 268091
rect 317986 268079 318014 268125
rect 322192 268113 322198 268125
rect 322250 268113 322256 268165
rect 322288 268113 322294 268165
rect 322346 268153 322352 268165
rect 328048 268153 328054 268165
rect 322346 268125 328054 268153
rect 322346 268113 322352 268125
rect 328048 268113 328054 268125
rect 328106 268113 328112 268165
rect 328240 268113 328246 268165
rect 328298 268153 328304 268165
rect 334960 268153 334966 268165
rect 328298 268125 334966 268153
rect 328298 268113 328304 268125
rect 334960 268113 334966 268125
rect 335018 268113 335024 268165
rect 335074 268125 356030 268153
rect 317794 268051 318014 268079
rect 275728 268005 275734 268017
rect 253570 267977 253790 268005
rect 255874 267977 275734 268005
rect 243088 267891 243094 267943
rect 243146 267931 243152 267943
rect 255874 267931 255902 267977
rect 275728 267965 275734 267977
rect 275786 267965 275792 268017
rect 296656 267965 296662 268017
rect 296714 268005 296720 268017
rect 308272 268005 308278 268017
rect 296714 267977 308278 268005
rect 296714 267965 296720 267977
rect 308272 267965 308278 267977
rect 308330 267965 308336 268017
rect 312592 267965 312598 268017
rect 312650 268005 312656 268017
rect 317794 268005 317822 268051
rect 321424 268039 321430 268091
rect 321482 268079 321488 268091
rect 326608 268079 326614 268091
rect 321482 268051 326614 268079
rect 321482 268039 321488 268051
rect 326608 268039 326614 268051
rect 326666 268039 326672 268091
rect 326704 268039 326710 268091
rect 326762 268079 326768 268091
rect 335074 268079 335102 268125
rect 326762 268051 335102 268079
rect 326762 268039 326768 268051
rect 347152 268039 347158 268091
rect 347210 268079 347216 268091
rect 355888 268079 355894 268091
rect 347210 268051 355894 268079
rect 347210 268039 347216 268051
rect 355888 268039 355894 268051
rect 355946 268039 355952 268091
rect 356002 268079 356030 268125
rect 357424 268113 357430 268165
rect 357482 268153 357488 268165
rect 369232 268153 369238 268165
rect 357482 268125 369238 268153
rect 357482 268113 357488 268125
rect 369232 268113 369238 268125
rect 369290 268113 369296 268165
rect 371824 268113 371830 268165
rect 371882 268153 371888 268165
rect 388240 268153 388246 268165
rect 371882 268125 388246 268153
rect 371882 268113 371888 268125
rect 388240 268113 388246 268125
rect 388298 268113 388304 268165
rect 388354 268153 388382 268199
rect 388432 268187 388438 268239
rect 388490 268227 388496 268239
rect 411280 268227 411286 268239
rect 388490 268199 411286 268227
rect 388490 268187 388496 268199
rect 411280 268187 411286 268199
rect 411338 268187 411344 268239
rect 398224 268153 398230 268165
rect 388354 268125 398230 268153
rect 398224 268113 398230 268125
rect 398282 268113 398288 268165
rect 371440 268079 371446 268091
rect 356002 268051 371446 268079
rect 371440 268039 371446 268051
rect 371498 268039 371504 268091
rect 372688 268039 372694 268091
rect 372746 268079 372752 268091
rect 372746 268051 388286 268079
rect 372746 268039 372752 268051
rect 312650 267977 317822 268005
rect 312650 267965 312656 267977
rect 317872 267965 317878 268017
rect 317930 268005 317936 268017
rect 328432 268005 328438 268017
rect 317930 267977 328438 268005
rect 317930 267965 317936 267977
rect 328432 267965 328438 267977
rect 328490 267965 328496 268017
rect 328528 267965 328534 268017
rect 328586 268005 328592 268017
rect 345328 268005 345334 268017
rect 328586 267977 345334 268005
rect 328586 267965 328592 267977
rect 345328 267965 345334 267977
rect 345386 267965 345392 268017
rect 349840 267965 349846 268017
rect 349898 268005 349904 268017
rect 349898 267977 357662 268005
rect 349898 267965 349904 267977
rect 243146 267903 255902 267931
rect 243146 267891 243152 267903
rect 266608 267891 266614 267943
rect 266666 267931 266672 267943
rect 355408 267931 355414 267943
rect 266666 267903 355414 267931
rect 266666 267891 266672 267903
rect 355408 267891 355414 267903
rect 355466 267891 355472 267943
rect 357634 267931 357662 267977
rect 358672 267965 358678 268017
rect 358730 268005 358736 268017
rect 368848 268005 368854 268017
rect 358730 267977 368854 268005
rect 358730 267965 358736 267977
rect 368848 267965 368854 267977
rect 368906 267965 368912 268017
rect 368944 267965 368950 268017
rect 369002 268005 369008 268017
rect 374224 268005 374230 268017
rect 369002 267977 374230 268005
rect 369002 267965 369008 267977
rect 374224 267965 374230 267977
rect 374282 267965 374288 268017
rect 374704 267965 374710 268017
rect 374762 268005 374768 268017
rect 378832 268005 378838 268017
rect 374762 267977 378838 268005
rect 374762 267965 374768 267977
rect 378832 267965 378838 267977
rect 378890 267965 378896 268017
rect 379216 267965 379222 268017
rect 379274 268005 379280 268017
rect 385360 268005 385366 268017
rect 379274 267977 385366 268005
rect 379274 267965 379280 267977
rect 385360 267965 385366 267977
rect 385418 267965 385424 268017
rect 368752 267931 368758 267943
rect 357634 267903 368758 267931
rect 368752 267891 368758 267903
rect 368810 267891 368816 267943
rect 370960 267891 370966 267943
rect 371018 267931 371024 267943
rect 376624 267931 376630 267943
rect 371018 267903 376630 267931
rect 371018 267891 371024 267903
rect 376624 267891 376630 267903
rect 376682 267891 376688 267943
rect 377200 267891 377206 267943
rect 377258 267931 377264 267943
rect 380272 267931 380278 267943
rect 377258 267903 380278 267931
rect 377258 267891 377264 267903
rect 380272 267891 380278 267903
rect 380330 267891 380336 267943
rect 380368 267891 380374 267943
rect 380426 267931 380432 267943
rect 382960 267931 382966 267943
rect 380426 267903 382966 267931
rect 380426 267891 380432 267903
rect 382960 267891 382966 267903
rect 383018 267891 383024 267943
rect 383056 267891 383062 267943
rect 383114 267931 383120 267943
rect 388144 267931 388150 267943
rect 383114 267903 388150 267931
rect 383114 267891 383120 267903
rect 388144 267891 388150 267903
rect 388202 267891 388208 267943
rect 388258 267931 388286 268051
rect 388912 268039 388918 268091
rect 388970 268079 388976 268091
rect 572464 268079 572470 268091
rect 388970 268051 572470 268079
rect 388970 268039 388976 268051
rect 572464 268039 572470 268051
rect 572522 268039 572528 268091
rect 389008 267965 389014 268017
rect 389066 268005 389072 268017
rect 397552 268005 397558 268017
rect 389066 267977 397558 268005
rect 389066 267965 389072 267977
rect 397552 267965 397558 267977
rect 397610 267965 397616 268017
rect 393808 267931 393814 267943
rect 388258 267903 393814 267931
rect 393808 267891 393814 267903
rect 393866 267891 393872 267943
rect 393904 267891 393910 267943
rect 393962 267931 393968 267943
rect 399376 267931 399382 267943
rect 393962 267903 399382 267931
rect 393962 267891 393968 267903
rect 399376 267891 399382 267903
rect 399434 267891 399440 267943
rect 65008 267817 65014 267869
rect 65066 267857 65072 267869
rect 65066 267829 74942 267857
rect 65066 267817 65072 267829
rect 74914 267783 74942 267829
rect 221968 267817 221974 267869
rect 222026 267857 222032 267869
rect 256144 267857 256150 267869
rect 222026 267829 256150 267857
rect 222026 267817 222032 267829
rect 256144 267817 256150 267829
rect 256202 267817 256208 267869
rect 267664 267817 267670 267869
rect 267722 267857 267728 267869
rect 357328 267857 357334 267869
rect 267722 267829 357334 267857
rect 267722 267817 267728 267829
rect 357328 267817 357334 267829
rect 357386 267817 357392 267869
rect 359056 267817 359062 267869
rect 359114 267857 359120 267869
rect 388816 267857 388822 267869
rect 359114 267829 388822 267857
rect 359114 267817 359120 267829
rect 388816 267817 388822 267829
rect 388874 267817 388880 267869
rect 389104 267817 389110 267869
rect 389162 267857 389168 267869
rect 401104 267857 401110 267869
rect 389162 267829 401110 267857
rect 389162 267817 389168 267829
rect 401104 267817 401110 267829
rect 401162 267817 401168 267869
rect 77776 267783 77782 267795
rect 74914 267755 77782 267783
rect 77776 267743 77782 267755
rect 77834 267743 77840 267795
rect 290608 267743 290614 267795
rect 290666 267783 290672 267795
rect 315088 267783 315094 267795
rect 290666 267755 315094 267783
rect 290666 267743 290672 267755
rect 315088 267743 315094 267755
rect 315146 267743 315152 267795
rect 315184 267743 315190 267795
rect 315242 267783 315248 267795
rect 322288 267783 322294 267795
rect 315242 267755 322294 267783
rect 315242 267743 315248 267755
rect 322288 267743 322294 267755
rect 322346 267743 322352 267795
rect 322384 267743 322390 267795
rect 322442 267783 322448 267795
rect 326320 267783 326326 267795
rect 322442 267755 326326 267783
rect 322442 267743 322448 267755
rect 326320 267743 326326 267755
rect 326378 267743 326384 267795
rect 326416 267743 326422 267795
rect 326474 267783 326480 267795
rect 327568 267783 327574 267795
rect 326474 267755 327574 267783
rect 326474 267743 326480 267755
rect 327568 267743 327574 267755
rect 327626 267743 327632 267795
rect 328048 267743 328054 267795
rect 328106 267783 328112 267795
rect 329296 267783 329302 267795
rect 328106 267755 329302 267783
rect 328106 267743 328112 267755
rect 329296 267743 329302 267755
rect 329354 267743 329360 267795
rect 329392 267743 329398 267795
rect 329450 267783 329456 267795
rect 332560 267783 332566 267795
rect 329450 267755 332566 267783
rect 329450 267743 329456 267755
rect 332560 267743 332566 267755
rect 332618 267743 332624 267795
rect 336880 267743 336886 267795
rect 336938 267783 336944 267795
rect 628432 267783 628438 267795
rect 336938 267755 628438 267783
rect 336938 267743 336944 267755
rect 628432 267743 628438 267755
rect 628490 267743 628496 267795
rect 255664 267669 255670 267721
rect 255722 267709 255728 267721
rect 267760 267709 267766 267721
rect 255722 267681 267766 267709
rect 255722 267669 255728 267681
rect 267760 267669 267766 267681
rect 267818 267669 267824 267721
rect 298096 267669 298102 267721
rect 298154 267709 298160 267721
rect 317008 267709 317014 267721
rect 298154 267681 317014 267709
rect 298154 267669 298160 267681
rect 317008 267669 317014 267681
rect 317066 267669 317072 267721
rect 317296 267669 317302 267721
rect 317354 267709 317360 267721
rect 318448 267709 318454 267721
rect 317354 267681 318454 267709
rect 317354 267669 317360 267681
rect 318448 267669 318454 267681
rect 318506 267669 318512 267721
rect 318544 267669 318550 267721
rect 318602 267709 318608 267721
rect 318602 267681 328862 267709
rect 318602 267669 318608 267681
rect 289456 267595 289462 267647
rect 289514 267635 289520 267647
rect 289514 267607 300158 267635
rect 289514 267595 289520 267607
rect 267856 267521 267862 267573
rect 267914 267561 267920 267573
rect 287920 267561 287926 267573
rect 267914 267533 287926 267561
rect 267914 267521 267920 267533
rect 287920 267521 287926 267533
rect 287978 267521 287984 267573
rect 290320 267521 290326 267573
rect 290378 267561 290384 267573
rect 300016 267561 300022 267573
rect 290378 267533 300022 267561
rect 290378 267521 290384 267533
rect 300016 267521 300022 267533
rect 300074 267521 300080 267573
rect 300130 267561 300158 267607
rect 300400 267595 300406 267647
rect 300458 267635 300464 267647
rect 328720 267635 328726 267647
rect 300458 267607 328726 267635
rect 300458 267595 300464 267607
rect 328720 267595 328726 267607
rect 328778 267595 328784 267647
rect 328834 267635 328862 267681
rect 328912 267669 328918 267721
rect 328970 267709 328976 267721
rect 349840 267709 349846 267721
rect 328970 267681 349846 267709
rect 328970 267669 328976 267681
rect 349840 267669 349846 267681
rect 349898 267669 349904 267721
rect 352240 267669 352246 267721
rect 352298 267709 352304 267721
rect 356848 267709 356854 267721
rect 352298 267681 356854 267709
rect 352298 267669 352304 267681
rect 356848 267669 356854 267681
rect 356906 267669 356912 267721
rect 356944 267669 356950 267721
rect 357002 267709 357008 267721
rect 366736 267709 366742 267721
rect 357002 267681 366742 267709
rect 357002 267669 357008 267681
rect 366736 267669 366742 267681
rect 366794 267669 366800 267721
rect 366832 267669 366838 267721
rect 366890 267709 366896 267721
rect 369328 267709 369334 267721
rect 366890 267681 369334 267709
rect 366890 267669 366896 267681
rect 369328 267669 369334 267681
rect 369386 267669 369392 267721
rect 369442 267681 377342 267709
rect 330640 267635 330646 267647
rect 328834 267607 330646 267635
rect 330640 267595 330646 267607
rect 330698 267595 330704 267647
rect 332560 267595 332566 267647
rect 332618 267635 332624 267647
rect 337648 267635 337654 267647
rect 332618 267607 337654 267635
rect 332618 267595 332624 267607
rect 337648 267595 337654 267607
rect 337706 267595 337712 267647
rect 353680 267635 353686 267647
rect 338338 267607 353686 267635
rect 338338 267561 338366 267607
rect 353680 267595 353686 267607
rect 353738 267595 353744 267647
rect 354256 267595 354262 267647
rect 354314 267635 354320 267647
rect 366640 267635 366646 267647
rect 354314 267607 366646 267635
rect 354314 267595 354320 267607
rect 366640 267595 366646 267607
rect 366698 267595 366704 267647
rect 366928 267595 366934 267647
rect 366986 267635 366992 267647
rect 369442 267635 369470 267681
rect 366986 267607 369470 267635
rect 366986 267595 366992 267607
rect 372880 267595 372886 267647
rect 372938 267635 372944 267647
rect 377200 267635 377206 267647
rect 372938 267607 377206 267635
rect 372938 267595 372944 267607
rect 377200 267595 377206 267607
rect 377258 267595 377264 267647
rect 377314 267635 377342 267681
rect 377488 267669 377494 267721
rect 377546 267709 377552 267721
rect 379984 267709 379990 267721
rect 377546 267681 379990 267709
rect 377546 267669 377552 267681
rect 379984 267669 379990 267681
rect 380042 267669 380048 267721
rect 380080 267669 380086 267721
rect 380138 267709 380144 267721
rect 383056 267709 383062 267721
rect 380138 267681 383062 267709
rect 380138 267669 380144 267681
rect 383056 267669 383062 267681
rect 383114 267669 383120 267721
rect 515440 267709 515446 267721
rect 384034 267681 515446 267709
rect 377314 267607 378686 267635
rect 347152 267561 347158 267573
rect 300130 267533 338366 267561
rect 338434 267533 347158 267561
rect 265744 267447 265750 267499
rect 265802 267487 265808 267499
rect 317200 267487 317206 267499
rect 265802 267459 317206 267487
rect 265802 267447 265808 267459
rect 317200 267447 317206 267459
rect 317258 267447 317264 267499
rect 317680 267447 317686 267499
rect 317738 267487 317744 267499
rect 327760 267487 327766 267499
rect 317738 267459 327766 267487
rect 317738 267447 317744 267459
rect 327760 267447 327766 267459
rect 327818 267447 327824 267499
rect 337456 267487 337462 267499
rect 328066 267459 337462 267487
rect 291472 267373 291478 267425
rect 291530 267413 291536 267425
rect 299920 267413 299926 267425
rect 291530 267385 299926 267413
rect 291530 267373 291536 267385
rect 299920 267373 299926 267385
rect 299978 267373 299984 267425
rect 300016 267373 300022 267425
rect 300074 267413 300080 267425
rect 327952 267413 327958 267425
rect 300074 267385 327958 267413
rect 300074 267373 300080 267385
rect 327952 267373 327958 267385
rect 328010 267373 328016 267425
rect 258832 267299 258838 267351
rect 258890 267339 258896 267351
rect 321424 267339 321430 267351
rect 258890 267311 321430 267339
rect 258890 267299 258896 267311
rect 321424 267299 321430 267311
rect 321482 267299 321488 267351
rect 321520 267299 321526 267351
rect 321578 267339 321584 267351
rect 328066 267339 328094 267459
rect 337456 267447 337462 267459
rect 337514 267447 337520 267499
rect 338434 267487 338462 267533
rect 347152 267521 347158 267533
rect 347210 267521 347216 267573
rect 347824 267521 347830 267573
rect 347882 267561 347888 267573
rect 348976 267561 348982 267573
rect 347882 267533 348982 267561
rect 347882 267521 347888 267533
rect 348976 267521 348982 267533
rect 349034 267521 349040 267573
rect 356944 267561 356950 267573
rect 356002 267533 356950 267561
rect 337570 267459 338462 267487
rect 328336 267373 328342 267425
rect 328394 267413 328400 267425
rect 337570 267413 337598 267459
rect 338800 267447 338806 267499
rect 338858 267487 338864 267499
rect 348496 267487 348502 267499
rect 338858 267459 348502 267487
rect 338858 267447 338864 267459
rect 348496 267447 348502 267459
rect 348554 267447 348560 267499
rect 349840 267487 349846 267499
rect 348610 267459 349846 267487
rect 328394 267385 337598 267413
rect 328394 267373 328400 267385
rect 337936 267373 337942 267425
rect 337994 267413 338000 267425
rect 343696 267413 343702 267425
rect 337994 267385 343702 267413
rect 337994 267373 338000 267385
rect 343696 267373 343702 267385
rect 343754 267373 343760 267425
rect 348208 267373 348214 267425
rect 348266 267413 348272 267425
rect 348610 267413 348638 267459
rect 349840 267447 349846 267459
rect 349898 267447 349904 267499
rect 350704 267447 350710 267499
rect 350762 267487 350768 267499
rect 356002 267487 356030 267533
rect 356944 267521 356950 267533
rect 357002 267521 357008 267573
rect 361552 267521 361558 267573
rect 361610 267561 361616 267573
rect 377104 267561 377110 267573
rect 361610 267533 377110 267561
rect 361610 267521 361616 267533
rect 377104 267521 377110 267533
rect 377162 267521 377168 267573
rect 378658 267561 378686 267607
rect 378736 267595 378742 267647
rect 378794 267635 378800 267647
rect 384034 267635 384062 267681
rect 515440 267669 515446 267681
rect 515498 267669 515504 267721
rect 391984 267635 391990 267647
rect 378794 267607 384062 267635
rect 384130 267607 391990 267635
rect 378794 267595 378800 267607
rect 384130 267561 384158 267607
rect 391984 267595 391990 267607
rect 392042 267595 392048 267647
rect 396592 267595 396598 267647
rect 396650 267635 396656 267647
rect 397168 267635 397174 267647
rect 396650 267607 397174 267635
rect 396650 267595 396656 267607
rect 397168 267595 397174 267607
rect 397226 267595 397232 267647
rect 397264 267595 397270 267647
rect 397322 267635 397328 267647
rect 411856 267635 411862 267647
rect 397322 267607 411862 267635
rect 397322 267595 397328 267607
rect 411856 267595 411862 267607
rect 411914 267595 411920 267647
rect 378658 267533 384158 267561
rect 384208 267521 384214 267573
rect 384266 267561 384272 267573
rect 384266 267533 397886 267561
rect 384266 267521 384272 267533
rect 350762 267459 356030 267487
rect 350762 267447 350768 267459
rect 356848 267447 356854 267499
rect 356906 267487 356912 267499
rect 356906 267459 366590 267487
rect 356906 267447 356912 267459
rect 348266 267385 348638 267413
rect 348266 267373 348272 267385
rect 348688 267373 348694 267425
rect 348746 267413 348752 267425
rect 366448 267413 366454 267425
rect 348746 267385 366454 267413
rect 348746 267373 348752 267385
rect 366448 267373 366454 267385
rect 366506 267373 366512 267425
rect 321578 267311 328094 267339
rect 321578 267299 321584 267311
rect 328240 267299 328246 267351
rect 328298 267339 328304 267351
rect 347824 267339 347830 267351
rect 328298 267311 347830 267339
rect 328298 267299 328304 267311
rect 347824 267299 347830 267311
rect 347882 267299 347888 267351
rect 348496 267299 348502 267351
rect 348554 267339 348560 267351
rect 358672 267339 358678 267351
rect 348554 267311 358678 267339
rect 348554 267299 348560 267311
rect 358672 267299 358678 267311
rect 358730 267299 358736 267351
rect 267568 267225 267574 267277
rect 267626 267265 267632 267277
rect 268048 267265 268054 267277
rect 267626 267237 268054 267265
rect 267626 267225 267632 267237
rect 268048 267225 268054 267237
rect 268106 267225 268112 267277
rect 292528 267225 292534 267277
rect 292586 267265 292592 267277
rect 299824 267265 299830 267277
rect 292586 267237 299830 267265
rect 292586 267225 292592 267237
rect 299824 267225 299830 267237
rect 299882 267225 299888 267277
rect 299920 267225 299926 267277
rect 299978 267265 299984 267277
rect 348688 267265 348694 267277
rect 299978 267237 348694 267265
rect 299978 267225 299984 267237
rect 348688 267225 348694 267237
rect 348746 267225 348752 267277
rect 359056 267265 359062 267277
rect 348802 267237 359062 267265
rect 251632 267151 251638 267203
rect 251690 267191 251696 267203
rect 315184 267191 315190 267203
rect 251690 267163 315190 267191
rect 251690 267151 251696 267163
rect 315184 267151 315190 267163
rect 315242 267151 315248 267203
rect 317104 267151 317110 267203
rect 317162 267191 317168 267203
rect 317776 267191 317782 267203
rect 317162 267163 317782 267191
rect 317162 267151 317168 267163
rect 317776 267151 317782 267163
rect 317834 267151 317840 267203
rect 317890 267163 318110 267191
rect 293584 267077 293590 267129
rect 293642 267117 293648 267129
rect 299728 267117 299734 267129
rect 293642 267089 299734 267117
rect 293642 267077 293648 267089
rect 299728 267077 299734 267089
rect 299786 267077 299792 267129
rect 299824 267077 299830 267129
rect 299882 267117 299888 267129
rect 317890 267117 317918 267163
rect 299882 267089 317918 267117
rect 318082 267117 318110 267163
rect 318160 267151 318166 267203
rect 318218 267191 318224 267203
rect 328240 267191 328246 267203
rect 318218 267163 328246 267191
rect 318218 267151 318224 267163
rect 328240 267151 328246 267163
rect 328298 267151 328304 267203
rect 328432 267151 328438 267203
rect 328490 267191 328496 267203
rect 337936 267191 337942 267203
rect 328490 267163 337942 267191
rect 328490 267151 328496 267163
rect 337936 267151 337942 267163
rect 337994 267151 338000 267203
rect 338032 267151 338038 267203
rect 338090 267191 338096 267203
rect 348208 267191 348214 267203
rect 338090 267163 348214 267191
rect 338090 267151 338096 267163
rect 348208 267151 348214 267163
rect 348266 267151 348272 267203
rect 348592 267151 348598 267203
rect 348650 267191 348656 267203
rect 348802 267191 348830 267237
rect 359056 267225 359062 267237
rect 359114 267225 359120 267277
rect 359152 267225 359158 267277
rect 359210 267265 359216 267277
rect 366562 267265 366590 267459
rect 366640 267447 366646 267499
rect 366698 267487 366704 267499
rect 367888 267487 367894 267499
rect 366698 267459 367894 267487
rect 366698 267447 366704 267459
rect 367888 267447 367894 267459
rect 367946 267447 367952 267499
rect 368176 267447 368182 267499
rect 368234 267487 368240 267499
rect 397744 267487 397750 267499
rect 368234 267459 397750 267487
rect 368234 267447 368240 267459
rect 397744 267447 397750 267459
rect 397802 267447 397808 267499
rect 397858 267487 397886 267533
rect 397936 267521 397942 267573
rect 397994 267561 398000 267573
rect 408784 267561 408790 267573
rect 397994 267533 408790 267561
rect 397994 267521 398000 267533
rect 408784 267521 408790 267533
rect 408842 267521 408848 267573
rect 406000 267487 406006 267499
rect 397858 267459 406006 267487
rect 406000 267447 406006 267459
rect 406058 267447 406064 267499
rect 367408 267373 367414 267425
rect 367466 267413 367472 267425
rect 367466 267385 377534 267413
rect 367466 267373 367472 267385
rect 366736 267299 366742 267351
rect 366794 267339 366800 267351
rect 368176 267339 368182 267351
rect 366794 267311 368182 267339
rect 366794 267299 366800 267311
rect 368176 267299 368182 267311
rect 368234 267299 368240 267351
rect 368464 267299 368470 267351
rect 368522 267339 368528 267351
rect 377392 267339 377398 267351
rect 368522 267311 377398 267339
rect 368522 267299 368528 267311
rect 377392 267299 377398 267311
rect 377450 267299 377456 267351
rect 377506 267339 377534 267385
rect 377584 267373 377590 267425
rect 377642 267413 377648 267425
rect 377642 267385 378686 267413
rect 377642 267373 377648 267385
rect 378544 267339 378550 267351
rect 377506 267311 378550 267339
rect 378544 267299 378550 267311
rect 378602 267299 378608 267351
rect 378658 267339 378686 267385
rect 378928 267373 378934 267425
rect 378986 267413 378992 267425
rect 392944 267413 392950 267425
rect 378986 267385 392950 267413
rect 378986 267373 378992 267385
rect 392944 267373 392950 267385
rect 393002 267373 393008 267425
rect 399568 267413 399574 267425
rect 396706 267385 399574 267413
rect 387760 267339 387766 267351
rect 378658 267311 387766 267339
rect 387760 267299 387766 267311
rect 387818 267299 387824 267351
rect 388816 267299 388822 267351
rect 388874 267339 388880 267351
rect 396706 267339 396734 267385
rect 399568 267373 399574 267385
rect 399626 267373 399632 267425
rect 408976 267373 408982 267425
rect 409034 267413 409040 267425
rect 426256 267413 426262 267425
rect 409034 267385 426262 267413
rect 409034 267373 409040 267385
rect 426256 267373 426262 267385
rect 426314 267373 426320 267425
rect 388874 267311 396734 267339
rect 388874 267299 388880 267311
rect 396784 267299 396790 267351
rect 396842 267339 396848 267351
rect 413776 267339 413782 267351
rect 396842 267311 413782 267339
rect 396842 267299 396848 267311
rect 413776 267299 413782 267311
rect 413834 267299 413840 267351
rect 367984 267265 367990 267277
rect 359210 267237 366494 267265
rect 366562 267237 367990 267265
rect 359210 267225 359216 267237
rect 348650 267163 348830 267191
rect 348650 267151 348656 267163
rect 348976 267151 348982 267203
rect 349034 267191 349040 267203
rect 354256 267191 354262 267203
rect 349034 267163 354262 267191
rect 349034 267151 349040 267163
rect 354256 267151 354262 267163
rect 354314 267151 354320 267203
rect 355024 267151 355030 267203
rect 355082 267191 355088 267203
rect 366160 267191 366166 267203
rect 355082 267163 366166 267191
rect 355082 267151 355088 267163
rect 366160 267151 366166 267163
rect 366218 267151 366224 267203
rect 318082 267089 328718 267117
rect 299882 267077 299888 267089
rect 244240 267003 244246 267055
rect 244298 267043 244304 267055
rect 317296 267043 317302 267055
rect 244298 267015 317302 267043
rect 244298 267003 244304 267015
rect 317296 267003 317302 267015
rect 317354 267003 317360 267055
rect 317968 267003 317974 267055
rect 318026 267043 318032 267055
rect 326224 267043 326230 267055
rect 318026 267015 326230 267043
rect 318026 267003 318032 267015
rect 326224 267003 326230 267015
rect 326282 267003 326288 267055
rect 326320 267003 326326 267055
rect 326378 267043 326384 267055
rect 326378 267015 327518 267043
rect 326378 267003 326384 267015
rect 237424 266929 237430 266981
rect 237482 266969 237488 266981
rect 318352 266969 318358 266981
rect 237482 266941 318358 266969
rect 237482 266929 237488 266941
rect 318352 266929 318358 266941
rect 318410 266929 318416 266981
rect 318448 266929 318454 266981
rect 318506 266969 318512 266981
rect 318832 266969 318838 266981
rect 318506 266941 318838 266969
rect 318506 266929 318512 266941
rect 318832 266929 318838 266941
rect 318890 266929 318896 266981
rect 318928 266929 318934 266981
rect 318986 266969 318992 266981
rect 327376 266969 327382 266981
rect 318986 266941 327382 266969
rect 318986 266929 318992 266941
rect 327376 266929 327382 266941
rect 327434 266929 327440 266981
rect 327490 266969 327518 267015
rect 327568 267003 327574 267055
rect 327626 267043 327632 267055
rect 327952 267043 327958 267055
rect 327626 267015 327958 267043
rect 327626 267003 327632 267015
rect 327952 267003 327958 267015
rect 328010 267003 328016 267055
rect 328240 267003 328246 267055
rect 328298 267043 328304 267055
rect 328690 267043 328718 267089
rect 329008 267077 329014 267129
rect 329066 267117 329072 267129
rect 331888 267117 331894 267129
rect 329066 267089 331894 267117
rect 329066 267077 329072 267089
rect 331888 267077 331894 267089
rect 331946 267077 331952 267129
rect 366352 267117 366358 267129
rect 332002 267089 348254 267117
rect 332002 267043 332030 267089
rect 328298 267015 328574 267043
rect 328690 267015 332030 267043
rect 328298 267003 328304 267015
rect 328336 266969 328342 266981
rect 327490 266941 328342 266969
rect 328336 266929 328342 266941
rect 328394 266929 328400 266981
rect 328546 266969 328574 267015
rect 337168 267003 337174 267055
rect 337226 267043 337232 267055
rect 348226 267043 348254 267089
rect 348418 267089 366358 267117
rect 348418 267043 348446 267089
rect 366352 267077 366358 267089
rect 366410 267077 366416 267129
rect 366466 267117 366494 267237
rect 367984 267225 367990 267237
rect 368042 267225 368048 267277
rect 368368 267225 368374 267277
rect 368426 267265 368432 267277
rect 368752 267265 368758 267277
rect 368426 267237 368758 267265
rect 368426 267225 368432 267237
rect 368752 267225 368758 267237
rect 368810 267225 368816 267277
rect 369040 267225 369046 267277
rect 369098 267265 369104 267277
rect 374416 267265 374422 267277
rect 369098 267237 374422 267265
rect 369098 267225 369104 267237
rect 374416 267225 374422 267237
rect 374474 267225 374480 267277
rect 374800 267265 374806 267277
rect 374530 267237 374806 267265
rect 374224 267191 374230 267203
rect 367522 267163 374230 267191
rect 367522 267117 367550 267163
rect 374224 267151 374230 267163
rect 374282 267151 374288 267203
rect 374530 267191 374558 267237
rect 374800 267225 374806 267237
rect 374858 267225 374864 267277
rect 377104 267225 377110 267277
rect 377162 267265 377168 267277
rect 409072 267265 409078 267277
rect 377162 267237 409078 267265
rect 377162 267225 377168 267237
rect 409072 267225 409078 267237
rect 409130 267225 409136 267277
rect 374338 267163 374558 267191
rect 374626 267163 388958 267191
rect 366466 267089 367550 267117
rect 367888 267077 367894 267129
rect 367946 267117 367952 267129
rect 374338 267117 374366 267163
rect 367946 267089 374366 267117
rect 367946 267077 367952 267089
rect 374416 267077 374422 267129
rect 374474 267117 374480 267129
rect 374626 267117 374654 267163
rect 374474 267089 374654 267117
rect 374474 267077 374480 267089
rect 374800 267077 374806 267129
rect 374858 267117 374864 267129
rect 377488 267117 377494 267129
rect 374858 267089 377494 267117
rect 374858 267077 374864 267089
rect 377488 267077 377494 267089
rect 377546 267077 377552 267129
rect 377680 267077 377686 267129
rect 377738 267117 377744 267129
rect 386224 267117 386230 267129
rect 377738 267089 386230 267117
rect 377738 267077 377744 267089
rect 386224 267077 386230 267089
rect 386282 267077 386288 267129
rect 388930 267117 388958 267163
rect 389008 267151 389014 267203
rect 389066 267191 389072 267203
rect 412528 267191 412534 267203
rect 389066 267163 412534 267191
rect 389066 267151 389072 267163
rect 412528 267151 412534 267163
rect 412586 267151 412592 267203
rect 393040 267117 393046 267129
rect 388930 267089 393046 267117
rect 393040 267077 393046 267089
rect 393098 267077 393104 267129
rect 398320 267077 398326 267129
rect 398378 267117 398384 267129
rect 421456 267117 421462 267129
rect 398378 267089 421462 267117
rect 398378 267077 398384 267089
rect 421456 267077 421462 267089
rect 421514 267077 421520 267129
rect 337226 267015 348158 267043
rect 348226 267015 348446 267043
rect 337226 267003 337232 267015
rect 329968 266969 329974 266981
rect 328546 266941 329974 266969
rect 329968 266929 329974 266941
rect 330026 266929 330032 266981
rect 330064 266929 330070 266981
rect 330122 266969 330128 266981
rect 337360 266969 337366 266981
rect 330122 266941 337366 266969
rect 330122 266929 330128 266941
rect 337360 266929 337366 266941
rect 337418 266929 337424 266981
rect 337456 266929 337462 266981
rect 337514 266969 337520 266981
rect 348016 266969 348022 266981
rect 337514 266941 348022 266969
rect 337514 266929 337520 266941
rect 348016 266929 348022 266941
rect 348074 266929 348080 266981
rect 348130 266969 348158 267015
rect 349840 267003 349846 267055
rect 349898 267043 349904 267055
rect 366256 267043 366262 267055
rect 349898 267015 366262 267043
rect 349898 267003 349904 267015
rect 366256 267003 366262 267015
rect 366314 267003 366320 267055
rect 366370 267015 367742 267043
rect 349360 266969 349366 266981
rect 348130 266941 349366 266969
rect 349360 266929 349366 266941
rect 349418 266929 349424 266981
rect 353968 266929 353974 266981
rect 354026 266969 354032 266981
rect 366370 266969 366398 267015
rect 354026 266941 366398 266969
rect 354026 266929 354032 266941
rect 366544 266929 366550 266981
rect 366602 266969 366608 266981
rect 367600 266969 367606 266981
rect 366602 266941 367606 266969
rect 366602 266929 366608 266941
rect 367600 266929 367606 266941
rect 367658 266929 367664 266981
rect 367714 266969 367742 267015
rect 367984 267003 367990 267055
rect 368042 267043 368048 267055
rect 397264 267043 397270 267055
rect 368042 267015 397270 267043
rect 368042 267003 368048 267015
rect 397264 267003 397270 267015
rect 397322 267003 397328 267055
rect 399280 267003 399286 267055
rect 399338 267043 399344 267055
rect 408880 267043 408886 267055
rect 399338 267015 408886 267043
rect 399338 267003 399344 267015
rect 408880 267003 408886 267015
rect 408938 267003 408944 267055
rect 408976 266969 408982 266981
rect 367714 266941 408982 266969
rect 408976 266929 408982 266941
rect 409034 266929 409040 266981
rect 413392 266969 413398 266981
rect 409090 266941 413398 266969
rect 293776 266855 293782 266907
rect 293834 266895 293840 266907
rect 293834 266867 299678 266895
rect 293834 266855 293840 266867
rect 294256 266781 294262 266833
rect 294314 266821 294320 266833
rect 299650 266821 299678 266867
rect 299728 266855 299734 266907
rect 299786 266895 299792 266907
rect 377872 266895 377878 266907
rect 299786 266867 377878 266895
rect 299786 266855 299792 266867
rect 377872 266855 377878 266867
rect 377930 266855 377936 266907
rect 377968 266855 377974 266907
rect 378026 266895 378032 266907
rect 384208 266895 384214 266907
rect 378026 266867 384214 266895
rect 378026 266855 378032 266867
rect 384208 266855 384214 266867
rect 384266 266855 384272 266907
rect 391024 266895 391030 266907
rect 389122 266867 391030 266895
rect 369136 266821 369142 266833
rect 294314 266793 299534 266821
rect 299650 266793 369142 266821
rect 294314 266781 294320 266793
rect 287632 266707 287638 266759
rect 287690 266747 287696 266759
rect 296656 266747 296662 266759
rect 287690 266719 296662 266747
rect 287690 266707 287696 266719
rect 296656 266707 296662 266719
rect 296714 266707 296720 266759
rect 299506 266747 299534 266793
rect 369136 266781 369142 266793
rect 369194 266781 369200 266833
rect 369328 266781 369334 266833
rect 369386 266821 369392 266833
rect 369386 266793 378974 266821
rect 369386 266781 369392 266793
rect 378736 266747 378742 266759
rect 299506 266719 378742 266747
rect 378736 266707 378742 266719
rect 378794 266707 378800 266759
rect 378946 266747 378974 266793
rect 379024 266781 379030 266833
rect 379082 266821 379088 266833
rect 385456 266821 385462 266833
rect 379082 266793 385462 266821
rect 379082 266781 379088 266793
rect 385456 266781 385462 266793
rect 385514 266781 385520 266833
rect 389122 266747 389150 266867
rect 391024 266855 391030 266867
rect 391082 266855 391088 266907
rect 393040 266855 393046 266907
rect 393098 266895 393104 266907
rect 404464 266895 404470 266907
rect 393098 266867 404470 266895
rect 393098 266855 393104 266867
rect 404464 266855 404470 266867
rect 404522 266855 404528 266907
rect 406096 266855 406102 266907
rect 406154 266895 406160 266907
rect 407152 266895 407158 266907
rect 406154 266867 407158 266895
rect 406154 266855 406160 266867
rect 407152 266855 407158 266867
rect 407210 266855 407216 266907
rect 408496 266855 408502 266907
rect 408554 266895 408560 266907
rect 409090 266895 409118 266941
rect 413392 266929 413398 266941
rect 413450 266929 413456 266981
rect 408554 266867 409118 266895
rect 408554 266855 408560 266867
rect 397744 266781 397750 266833
rect 397802 266821 397808 266833
rect 403216 266821 403222 266833
rect 397802 266793 403222 266821
rect 397802 266781 397808 266793
rect 403216 266781 403222 266793
rect 403274 266781 403280 266833
rect 408592 266781 408598 266833
rect 408650 266821 408656 266833
rect 413680 266821 413686 266833
rect 408650 266793 413686 266821
rect 408650 266781 408656 266793
rect 413680 266781 413686 266793
rect 413738 266781 413744 266833
rect 389584 266747 389590 266759
rect 378946 266719 389150 266747
rect 389314 266719 389590 266747
rect 230032 266633 230038 266685
rect 230090 266673 230096 266685
rect 318160 266673 318166 266685
rect 230090 266645 318166 266673
rect 230090 266633 230096 266645
rect 318160 266633 318166 266645
rect 318218 266633 318224 266685
rect 318544 266633 318550 266685
rect 318602 266673 318608 266685
rect 326416 266673 326422 266685
rect 318602 266645 326422 266673
rect 318602 266633 318608 266645
rect 326416 266633 326422 266645
rect 326474 266633 326480 266685
rect 326512 266633 326518 266685
rect 326570 266673 326576 266685
rect 328048 266673 328054 266685
rect 326570 266645 328054 266673
rect 326570 266633 326576 266645
rect 328048 266633 328054 266645
rect 328106 266633 328112 266685
rect 337264 266673 337270 266685
rect 328450 266645 337270 266673
rect 295312 266559 295318 266611
rect 295370 266599 295376 266611
rect 328240 266599 328246 266611
rect 295370 266571 328246 266599
rect 295370 266559 295376 266571
rect 328240 266559 328246 266571
rect 328298 266559 328304 266611
rect 215728 266485 215734 266537
rect 215786 266525 215792 266537
rect 309808 266525 309814 266537
rect 215786 266497 309814 266525
rect 215786 266485 215792 266497
rect 309808 266485 309814 266497
rect 309866 266485 309872 266537
rect 310000 266485 310006 266537
rect 310058 266525 310064 266537
rect 312976 266525 312982 266537
rect 310058 266497 312982 266525
rect 310058 266485 310064 266497
rect 312976 266485 312982 266497
rect 313034 266485 313040 266537
rect 315088 266485 315094 266537
rect 315146 266525 315152 266537
rect 328450 266525 328478 266645
rect 337264 266633 337270 266645
rect 337322 266633 337328 266685
rect 337648 266633 337654 266685
rect 337706 266673 337712 266685
rect 367408 266673 367414 266685
rect 337706 266645 367414 266673
rect 337706 266633 337712 266645
rect 367408 266633 367414 266645
rect 367466 266633 367472 266685
rect 367600 266633 367606 266685
rect 367658 266673 367664 266685
rect 389314 266673 389342 266719
rect 389584 266707 389590 266719
rect 389642 266707 389648 266759
rect 393040 266707 393046 266759
rect 393098 266747 393104 266759
rect 407344 266747 407350 266759
rect 393098 266719 407350 266747
rect 393098 266707 393104 266719
rect 407344 266707 407350 266719
rect 407402 266707 407408 266759
rect 408688 266707 408694 266759
rect 408746 266747 408752 266759
rect 409648 266747 409654 266759
rect 408746 266719 409654 266747
rect 408746 266707 408752 266719
rect 409648 266707 409654 266719
rect 409706 266707 409712 266759
rect 367658 266645 389342 266673
rect 367658 266633 367664 266645
rect 389776 266633 389782 266685
rect 389834 266673 389840 266685
rect 433360 266673 433366 266685
rect 389834 266645 433366 266673
rect 389834 266633 389840 266645
rect 433360 266633 433366 266645
rect 433418 266633 433424 266685
rect 328912 266559 328918 266611
rect 328970 266599 328976 266611
rect 377680 266599 377686 266611
rect 328970 266571 377686 266599
rect 328970 266559 328976 266571
rect 377680 266559 377686 266571
rect 377738 266559 377744 266611
rect 377872 266559 377878 266611
rect 377930 266599 377936 266611
rect 378448 266599 378454 266611
rect 377930 266571 378454 266599
rect 377930 266559 377936 266571
rect 378448 266559 378454 266571
rect 378506 266559 378512 266611
rect 378544 266559 378550 266611
rect 378602 266599 378608 266611
rect 393040 266599 393046 266611
rect 378602 266571 393046 266599
rect 378602 266559 378608 266571
rect 393040 266559 393046 266571
rect 393098 266559 393104 266611
rect 406864 266559 406870 266611
rect 406922 266599 406928 266611
rect 407728 266599 407734 266611
rect 406922 266571 407734 266599
rect 406922 266559 406928 266571
rect 407728 266559 407734 266571
rect 407786 266559 407792 266611
rect 409072 266559 409078 266611
rect 409130 266599 409136 266611
rect 410320 266599 410326 266611
rect 409130 266571 410326 266599
rect 409130 266559 409136 266571
rect 410320 266559 410326 266571
rect 410378 266559 410384 266611
rect 315146 266497 328478 266525
rect 315146 266485 315152 266497
rect 328528 266485 328534 266537
rect 328586 266525 328592 266537
rect 338800 266525 338806 266537
rect 328586 266497 338806 266525
rect 328586 266485 328592 266497
rect 338800 266485 338806 266497
rect 338858 266485 338864 266537
rect 347824 266485 347830 266537
rect 347882 266525 347888 266537
rect 348592 266525 348598 266537
rect 347882 266497 348598 266525
rect 347882 266485 347888 266497
rect 348592 266485 348598 266497
rect 348650 266485 348656 266537
rect 349072 266485 349078 266537
rect 349130 266525 349136 266537
rect 357520 266525 357526 266537
rect 349130 266497 357526 266525
rect 349130 266485 349136 266497
rect 357520 266485 357526 266497
rect 357578 266485 357584 266537
rect 358288 266485 358294 266537
rect 358346 266525 358352 266537
rect 367408 266525 367414 266537
rect 358346 266497 367414 266525
rect 358346 266485 358352 266497
rect 367408 266485 367414 266497
rect 367466 266485 367472 266537
rect 367600 266485 367606 266537
rect 367658 266525 367664 266537
rect 447664 266525 447670 266537
rect 367658 266497 447670 266525
rect 367658 266485 367664 266497
rect 447664 266485 447670 266497
rect 447722 266485 447728 266537
rect 270640 266411 270646 266463
rect 270698 266451 270704 266463
rect 287920 266451 287926 266463
rect 270698 266423 287926 266451
rect 270698 266411 270704 266423
rect 287920 266411 287926 266423
rect 287978 266411 287984 266463
rect 295984 266411 295990 266463
rect 296042 266451 296048 266463
rect 389392 266451 389398 266463
rect 296042 266423 389398 266451
rect 296042 266411 296048 266423
rect 389392 266411 389398 266423
rect 389450 266411 389456 266463
rect 399088 266411 399094 266463
rect 399146 266451 399152 266463
rect 400240 266451 400246 266463
rect 399146 266423 400246 266451
rect 399146 266411 399152 266423
rect 400240 266411 400246 266423
rect 400298 266411 400304 266463
rect 400720 266411 400726 266463
rect 400778 266451 400784 266463
rect 406096 266451 406102 266463
rect 400778 266423 406102 266451
rect 400778 266411 400784 266423
rect 406096 266411 406102 266423
rect 406154 266411 406160 266463
rect 406576 266411 406582 266463
rect 406634 266451 406640 266463
rect 408592 266451 408598 266463
rect 406634 266423 408598 266451
rect 406634 266411 406640 266423
rect 408592 266411 408598 266423
rect 408650 266411 408656 266463
rect 287632 266337 287638 266389
rect 287690 266377 287696 266389
rect 296752 266377 296758 266389
rect 287690 266349 296758 266377
rect 287690 266337 287696 266349
rect 296752 266337 296758 266349
rect 296810 266337 296816 266389
rect 296848 266337 296854 266389
rect 296906 266377 296912 266389
rect 296906 266349 399230 266377
rect 296906 266337 296912 266349
rect 208528 266263 208534 266315
rect 208586 266303 208592 266315
rect 310000 266303 310006 266315
rect 208586 266275 310006 266303
rect 208586 266263 208592 266275
rect 310000 266263 310006 266275
rect 310058 266263 310064 266315
rect 310096 266263 310102 266315
rect 310154 266303 310160 266315
rect 317104 266303 317110 266315
rect 310154 266275 317110 266303
rect 310154 266263 310160 266275
rect 317104 266263 317110 266275
rect 317162 266263 317168 266315
rect 317200 266263 317206 266315
rect 317258 266303 317264 266315
rect 317584 266303 317590 266315
rect 317258 266275 317590 266303
rect 317258 266263 317264 266275
rect 317584 266263 317590 266275
rect 317642 266263 317648 266315
rect 317968 266263 317974 266315
rect 318026 266303 318032 266315
rect 318256 266303 318262 266315
rect 318026 266275 318262 266303
rect 318026 266263 318032 266275
rect 318256 266263 318262 266275
rect 318314 266263 318320 266315
rect 318928 266303 318934 266315
rect 318370 266275 318934 266303
rect 298000 266189 298006 266241
rect 298058 266229 298064 266241
rect 318160 266229 318166 266241
rect 298058 266201 318166 266229
rect 298058 266189 298064 266201
rect 318160 266189 318166 266201
rect 318218 266189 318224 266241
rect 201424 266115 201430 266167
rect 201482 266155 201488 266167
rect 310096 266155 310102 266167
rect 201482 266127 310102 266155
rect 201482 266115 201488 266127
rect 310096 266115 310102 266127
rect 310154 266115 310160 266167
rect 310192 266115 310198 266167
rect 310250 266155 310256 266167
rect 312880 266155 312886 266167
rect 310250 266127 312886 266155
rect 310250 266115 310256 266127
rect 312880 266115 312886 266127
rect 312938 266115 312944 266167
rect 312976 266115 312982 266167
rect 313034 266155 313040 266167
rect 318370 266155 318398 266275
rect 318928 266263 318934 266275
rect 318986 266263 318992 266315
rect 322480 266263 322486 266315
rect 322538 266303 322544 266315
rect 328624 266303 328630 266315
rect 322538 266275 328630 266303
rect 322538 266263 322544 266275
rect 328624 266263 328630 266275
rect 328682 266263 328688 266315
rect 328816 266263 328822 266315
rect 328874 266303 328880 266315
rect 346576 266303 346582 266315
rect 328874 266275 346582 266303
rect 328874 266263 328880 266275
rect 346576 266263 346582 266275
rect 346634 266263 346640 266315
rect 348016 266263 348022 266315
rect 348074 266303 348080 266315
rect 349840 266303 349846 266315
rect 348074 266275 349846 266303
rect 348074 266263 348080 266275
rect 349840 266263 349846 266275
rect 349898 266263 349904 266315
rect 349936 266263 349942 266315
rect 349994 266303 350000 266315
rect 357808 266303 357814 266315
rect 349994 266275 357814 266303
rect 349994 266263 350000 266275
rect 357808 266263 357814 266275
rect 357866 266263 357872 266315
rect 366448 266263 366454 266315
rect 366506 266303 366512 266315
rect 367312 266303 367318 266315
rect 366506 266275 367318 266303
rect 366506 266263 366512 266275
rect 367312 266263 367318 266275
rect 367370 266263 367376 266315
rect 367408 266263 367414 266315
rect 367466 266303 367472 266315
rect 393904 266303 393910 266315
rect 367466 266275 393910 266303
rect 367466 266263 367472 266275
rect 393904 266263 393910 266275
rect 393962 266263 393968 266315
rect 318448 266189 318454 266241
rect 318506 266229 318512 266241
rect 398320 266229 398326 266241
rect 318506 266201 398326 266229
rect 318506 266189 318512 266201
rect 398320 266189 398326 266201
rect 398378 266189 398384 266241
rect 399202 266229 399230 266349
rect 399568 266337 399574 266389
rect 399626 266377 399632 266389
rect 413200 266377 413206 266389
rect 399626 266349 413206 266377
rect 399626 266337 399632 266349
rect 413200 266337 413206 266349
rect 413258 266337 413264 266389
rect 501616 266337 501622 266389
rect 501674 266377 501680 266389
rect 569872 266377 569878 266389
rect 501674 266349 569878 266377
rect 501674 266337 501680 266349
rect 569872 266337 569878 266349
rect 569930 266337 569936 266389
rect 399376 266263 399382 266315
rect 399434 266303 399440 266315
rect 461968 266303 461974 266315
rect 399434 266275 461974 266303
rect 399434 266263 399440 266275
rect 461968 266263 461974 266275
rect 462026 266263 462032 266315
rect 414352 266229 414358 266241
rect 399202 266201 414358 266229
rect 414352 266189 414358 266201
rect 414410 266189 414416 266241
rect 313034 266127 318398 266155
rect 313034 266115 313040 266127
rect 318832 266115 318838 266167
rect 318890 266155 318896 266167
rect 331696 266155 331702 266167
rect 318890 266127 331702 266155
rect 318890 266115 318896 266127
rect 331696 266115 331702 266127
rect 331754 266115 331760 266167
rect 331888 266115 331894 266167
rect 331946 266155 331952 266167
rect 349936 266155 349942 266167
rect 331946 266127 349942 266155
rect 331946 266115 331952 266127
rect 349936 266115 349942 266127
rect 349994 266115 350000 266167
rect 351280 266115 351286 266167
rect 351338 266155 351344 266167
rect 359152 266155 359158 266167
rect 351338 266127 359158 266155
rect 351338 266115 351344 266127
rect 359152 266115 359158 266127
rect 359210 266115 359216 266167
rect 360016 266115 360022 266167
rect 360074 266155 360080 266167
rect 476176 266155 476182 266167
rect 360074 266127 476182 266155
rect 360074 266115 360080 266127
rect 476176 266115 476182 266127
rect 476234 266115 476240 266167
rect 298576 266041 298582 266093
rect 298634 266081 298640 266093
rect 428656 266081 428662 266093
rect 298634 266053 428662 266081
rect 298634 266041 298640 266053
rect 428656 266041 428662 266053
rect 428714 266041 428720 266093
rect 299728 265967 299734 266019
rect 299786 266007 299792 266019
rect 435664 266007 435670 266019
rect 299786 265979 435670 266007
rect 299786 265967 299792 265979
rect 435664 265967 435670 265979
rect 435722 265967 435728 266019
rect 300304 265893 300310 265945
rect 300362 265933 300368 265945
rect 442864 265933 442870 265945
rect 300362 265905 442870 265933
rect 300362 265893 300368 265905
rect 442864 265893 442870 265905
rect 442922 265893 442928 265945
rect 288784 265819 288790 265871
rect 288842 265859 288848 265871
rect 300400 265859 300406 265871
rect 288842 265831 300406 265859
rect 288842 265819 288848 265831
rect 300400 265819 300406 265831
rect 300458 265819 300464 265871
rect 301264 265819 301270 265871
rect 301322 265859 301328 265871
rect 449968 265859 449974 265871
rect 301322 265831 449974 265859
rect 301322 265819 301328 265831
rect 449968 265819 449974 265831
rect 450026 265819 450032 265871
rect 287248 265745 287254 265797
rect 287306 265785 287312 265797
rect 298096 265785 298102 265797
rect 287306 265757 298102 265785
rect 287306 265745 287312 265757
rect 298096 265745 298102 265757
rect 298154 265745 298160 265797
rect 302320 265745 302326 265797
rect 302378 265785 302384 265797
rect 457168 265785 457174 265797
rect 302378 265757 457174 265785
rect 302378 265745 302384 265757
rect 457168 265745 457174 265757
rect 457226 265745 457232 265797
rect 302992 265671 302998 265723
rect 303050 265711 303056 265723
rect 312208 265711 312214 265723
rect 303050 265683 312214 265711
rect 303050 265671 303056 265683
rect 312208 265671 312214 265683
rect 312266 265671 312272 265723
rect 312880 265671 312886 265723
rect 312938 265711 312944 265723
rect 337168 265711 337174 265723
rect 312938 265683 337174 265711
rect 312938 265671 312944 265683
rect 337168 265671 337174 265683
rect 337226 265671 337232 265723
rect 337552 265671 337558 265723
rect 337610 265711 337616 265723
rect 464272 265711 464278 265723
rect 337610 265683 464278 265711
rect 337610 265671 337616 265683
rect 464272 265671 464278 265683
rect 464330 265671 464336 265723
rect 304048 265597 304054 265649
rect 304106 265637 304112 265649
rect 471376 265637 471382 265649
rect 304106 265609 471382 265637
rect 304106 265597 304112 265609
rect 471376 265597 471382 265609
rect 471434 265597 471440 265649
rect 257584 265523 257590 265575
rect 257642 265563 257648 265575
rect 269872 265563 269878 265575
rect 257642 265535 269878 265563
rect 257642 265523 257648 265535
rect 269872 265523 269878 265535
rect 269930 265523 269936 265575
rect 304720 265523 304726 265575
rect 304778 265563 304784 265575
rect 478576 265563 478582 265575
rect 304778 265535 478582 265563
rect 304778 265523 304784 265535
rect 478576 265523 478582 265535
rect 478634 265523 478640 265575
rect 306736 265449 306742 265501
rect 306794 265489 306800 265501
rect 492880 265489 492886 265501
rect 306794 265461 492886 265489
rect 306794 265449 306800 265461
rect 492880 265449 492886 265461
rect 492938 265449 492944 265501
rect 307312 265375 307318 265427
rect 307370 265415 307376 265427
rect 499888 265415 499894 265427
rect 307370 265387 499894 265415
rect 307370 265375 307376 265387
rect 499888 265375 499894 265387
rect 499946 265375 499952 265427
rect 308224 265301 308230 265353
rect 308282 265341 308288 265353
rect 507088 265341 507094 265353
rect 308282 265313 507094 265341
rect 308282 265301 308288 265313
rect 507088 265301 507094 265313
rect 507146 265301 507152 265353
rect 225328 265227 225334 265279
rect 225386 265267 225392 265279
rect 273616 265267 273622 265279
rect 225386 265239 273622 265267
rect 225386 265227 225392 265239
rect 273616 265227 273622 265239
rect 273674 265227 273680 265279
rect 308848 265227 308854 265279
rect 308906 265267 308912 265279
rect 510640 265267 510646 265279
rect 308906 265239 510646 265267
rect 308906 265227 308912 265239
rect 510640 265227 510646 265239
rect 510698 265227 510704 265279
rect 221680 265153 221686 265205
rect 221738 265193 221744 265205
rect 273136 265193 273142 265205
rect 221738 265165 273142 265193
rect 221738 265153 221744 265165
rect 273136 265153 273142 265165
rect 273194 265153 273200 265205
rect 309328 265153 309334 265205
rect 309386 265193 309392 265205
rect 514288 265193 514294 265205
rect 309386 265165 514294 265193
rect 309386 265153 309392 265165
rect 514288 265153 514294 265165
rect 514346 265153 514352 265205
rect 223120 265079 223126 265131
rect 223178 265119 223184 265131
rect 329008 265119 329014 265131
rect 223178 265091 329014 265119
rect 223178 265079 223184 265091
rect 329008 265079 329014 265091
rect 329066 265079 329072 265131
rect 329680 265079 329686 265131
rect 329738 265119 329744 265131
rect 332368 265119 332374 265131
rect 329738 265091 332374 265119
rect 329738 265079 329744 265091
rect 332368 265079 332374 265091
rect 332426 265079 332432 265131
rect 349840 265079 349846 265131
rect 349898 265119 349904 265131
rect 372976 265119 372982 265131
rect 349898 265091 372982 265119
rect 349898 265079 349904 265091
rect 372976 265079 372982 265091
rect 373034 265079 373040 265131
rect 376912 265079 376918 265131
rect 376970 265119 376976 265131
rect 611824 265119 611830 265131
rect 376970 265091 611830 265119
rect 376970 265079 376976 265091
rect 611824 265079 611830 265091
rect 611882 265079 611888 265131
rect 197872 265005 197878 265057
rect 197930 265045 197936 265057
rect 325840 265045 325846 265057
rect 197930 265017 325846 265045
rect 197930 265005 197936 265017
rect 325840 265005 325846 265017
rect 325898 265005 325904 265057
rect 326608 265005 326614 265057
rect 326666 265045 326672 265057
rect 333136 265045 333142 265057
rect 326666 265017 333142 265045
rect 326666 265005 326672 265017
rect 333136 265005 333142 265017
rect 333194 265005 333200 265057
rect 356848 265005 356854 265057
rect 356906 265045 356912 265057
rect 367600 265045 367606 265057
rect 356906 265017 367606 265045
rect 356906 265005 356912 265017
rect 367600 265005 367606 265017
rect 367658 265005 367664 265057
rect 368560 265045 368566 265057
rect 368482 265017 368566 265045
rect 81808 264931 81814 264983
rect 81866 264971 81872 264983
rect 90640 264971 90646 264983
rect 81866 264943 90646 264971
rect 81866 264931 81872 264943
rect 90640 264931 90646 264943
rect 90698 264931 90704 264983
rect 309808 264931 309814 264983
rect 309866 264971 309872 264983
rect 318352 264971 318358 264983
rect 309866 264943 318358 264971
rect 309866 264931 309872 264943
rect 318352 264931 318358 264943
rect 318410 264931 318416 264983
rect 318448 264931 318454 264983
rect 318506 264971 318512 264983
rect 318736 264971 318742 264983
rect 318506 264943 318742 264971
rect 318506 264931 318512 264943
rect 318736 264931 318742 264943
rect 318794 264931 318800 264983
rect 324112 264931 324118 264983
rect 324170 264971 324176 264983
rect 329296 264971 329302 264983
rect 324170 264943 329302 264971
rect 324170 264931 324176 264943
rect 329296 264931 329302 264943
rect 329354 264931 329360 264983
rect 347728 264931 347734 264983
rect 347786 264971 347792 264983
rect 368482 264971 368510 265017
rect 368560 265005 368566 265017
rect 368618 265005 368624 265057
rect 369136 265005 369142 265057
rect 369194 265045 369200 265057
rect 378640 265045 378646 265057
rect 369194 265017 378646 265045
rect 369194 265005 369200 265017
rect 378640 265005 378646 265017
rect 378698 265005 378704 265057
rect 379504 265005 379510 265057
rect 379562 265045 379568 265057
rect 633136 265045 633142 265057
rect 379562 265017 633142 265045
rect 379562 265005 379568 265017
rect 633136 265005 633142 265017
rect 633194 265005 633200 265057
rect 347786 264943 368510 264971
rect 347786 264931 347792 264943
rect 369520 264931 369526 264983
rect 369578 264971 369584 264983
rect 369578 264943 382526 264971
rect 369578 264931 369584 264943
rect 343696 264857 343702 264909
rect 343754 264897 343760 264909
rect 382384 264897 382390 264909
rect 343754 264869 382390 264897
rect 343754 264857 343760 264869
rect 382384 264857 382390 264869
rect 382442 264857 382448 264909
rect 382498 264897 382526 264943
rect 388624 264931 388630 264983
rect 388682 264971 388688 264983
rect 413200 264971 413206 264983
rect 388682 264943 413206 264971
rect 388682 264931 388688 264943
rect 413200 264931 413206 264943
rect 413258 264931 413264 264983
rect 455152 264931 455158 264983
rect 455210 264971 455216 264983
rect 475120 264971 475126 264983
rect 455210 264943 475126 264971
rect 455210 264931 455216 264943
rect 475120 264931 475126 264943
rect 475178 264931 475184 264983
rect 483856 264931 483862 264983
rect 483914 264971 483920 264983
rect 511120 264971 511126 264983
rect 483914 264943 511126 264971
rect 483914 264931 483920 264943
rect 511120 264931 511126 264943
rect 511178 264931 511184 264983
rect 551056 264897 551062 264909
rect 382498 264869 551062 264897
rect 551056 264857 551062 264869
rect 551114 264857 551120 264909
rect 158608 264487 158614 264539
rect 158666 264527 158672 264539
rect 161200 264527 161206 264539
rect 158666 264499 161206 264527
rect 158666 264487 158672 264499
rect 161200 264487 161206 264499
rect 161258 264487 161264 264539
rect 42256 264265 42262 264317
rect 42314 264305 42320 264317
rect 50512 264305 50518 264317
rect 42314 264277 50518 264305
rect 42314 264265 42320 264277
rect 50512 264265 50518 264277
rect 50570 264265 50576 264317
rect 77776 263599 77782 263651
rect 77834 263639 77840 263651
rect 87760 263639 87766 263651
rect 77834 263611 87766 263639
rect 77834 263599 77840 263611
rect 87760 263599 87766 263611
rect 87818 263599 87824 263651
rect 42640 263229 42646 263281
rect 42698 263269 42704 263281
rect 53392 263269 53398 263281
rect 42698 263241 53398 263269
rect 42698 263229 42704 263241
rect 53392 263229 53398 263241
rect 53450 263229 53456 263281
rect 42640 262267 42646 262319
rect 42698 262307 42704 262319
rect 56176 262307 56182 262319
rect 42698 262279 56182 262307
rect 42698 262267 42704 262279
rect 56176 262267 56182 262279
rect 56234 262267 56240 262319
rect 87760 260713 87766 260765
rect 87818 260753 87824 260765
rect 93328 260753 93334 260765
rect 87818 260725 93334 260753
rect 87818 260713 87824 260725
rect 93328 260713 93334 260725
rect 93386 260713 93392 260765
rect 90640 260639 90646 260691
rect 90698 260679 90704 260691
rect 102544 260679 102550 260691
rect 90698 260651 102550 260679
rect 90698 260639 90704 260651
rect 102544 260639 102550 260651
rect 102602 260639 102608 260691
rect 639280 256347 639286 256399
rect 639338 256387 639344 256399
rect 679792 256387 679798 256399
rect 639338 256359 679798 256387
rect 639338 256347 639344 256359
rect 679792 256347 679798 256359
rect 679850 256347 679856 256399
rect 93328 256273 93334 256325
rect 93386 256313 93392 256325
rect 97840 256313 97846 256325
rect 93386 256285 97846 256313
rect 93386 256273 93392 256285
rect 97840 256273 97846 256285
rect 97898 256273 97904 256325
rect 44560 255089 44566 255141
rect 44618 255129 44624 255141
rect 60400 255129 60406 255141
rect 44618 255101 60406 255129
rect 44618 255089 44624 255101
rect 60400 255089 60406 255101
rect 60458 255089 60464 255141
rect 632080 253501 632086 253513
rect 627874 253473 632086 253501
rect 625168 253387 625174 253439
rect 625226 253427 625232 253439
rect 627874 253427 627902 253473
rect 632080 253461 632086 253473
rect 632138 253461 632144 253513
rect 625226 253399 627902 253427
rect 625226 253387 625232 253399
rect 100144 252943 100150 252995
rect 100202 252983 100208 252995
rect 100720 252983 100726 252995
rect 100202 252955 100726 252983
rect 100202 252943 100208 252955
rect 100720 252943 100726 252955
rect 100778 252943 100784 252995
rect 191440 252425 191446 252477
rect 191498 252465 191504 252477
rect 193264 252465 193270 252477
rect 191498 252437 193270 252465
rect 191498 252425 191504 252437
rect 193264 252425 193270 252437
rect 193322 252425 193328 252477
rect 53776 252055 53782 252107
rect 53834 252095 53840 252107
rect 210640 252095 210646 252107
rect 53834 252067 210646 252095
rect 53834 252055 53840 252067
rect 210640 252055 210646 252067
rect 210698 252055 210704 252107
rect 45040 251981 45046 252033
rect 45098 252021 45104 252033
rect 206800 252021 206806 252033
rect 45098 251993 206806 252021
rect 45098 251981 45104 251993
rect 206800 251981 206806 251993
rect 206858 251981 206864 252033
rect 497488 251611 497494 251663
rect 497546 251651 497552 251663
rect 501616 251651 501622 251663
rect 497546 251623 501622 251651
rect 497546 251611 497552 251623
rect 501616 251611 501622 251623
rect 501674 251611 501680 251663
rect 674992 251611 674998 251663
rect 675050 251651 675056 251663
rect 676912 251651 676918 251663
rect 675050 251623 676918 251651
rect 675050 251611 675056 251623
rect 676912 251611 676918 251623
rect 676970 251611 676976 251663
rect 675088 251537 675094 251589
rect 675146 251577 675152 251589
rect 676816 251577 676822 251589
rect 675146 251549 676822 251577
rect 675146 251537 675152 251549
rect 676816 251537 676822 251549
rect 676874 251537 676880 251589
rect 674512 250945 674518 250997
rect 674570 250985 674576 250997
rect 675376 250985 675382 250997
rect 674570 250957 675382 250985
rect 674570 250945 674576 250957
rect 675376 250945 675382 250957
rect 675434 250945 675440 250997
rect 674608 250353 674614 250405
rect 674666 250393 674672 250405
rect 675472 250393 675478 250405
rect 674666 250365 675478 250393
rect 674666 250353 674672 250365
rect 675472 250353 675478 250365
rect 675530 250353 675536 250405
rect 42160 249835 42166 249887
rect 42218 249875 42224 249887
rect 42640 249875 42646 249887
rect 42218 249847 42646 249875
rect 42218 249835 42224 249847
rect 42640 249835 42646 249847
rect 42698 249835 42704 249887
rect 674128 249539 674134 249591
rect 674186 249579 674192 249591
rect 675376 249579 675382 249591
rect 674186 249551 675382 249579
rect 674186 249539 674192 249551
rect 675376 249539 675382 249551
rect 675434 249539 675440 249591
rect 613456 249095 613462 249147
rect 613514 249135 613520 249147
rect 625168 249135 625174 249147
rect 613514 249107 625174 249135
rect 613514 249095 613520 249107
rect 625168 249095 625174 249107
rect 625226 249095 625232 249147
rect 673936 247911 673942 247963
rect 673994 247951 674000 247963
rect 675376 247951 675382 247963
rect 673994 247923 675382 247951
rect 673994 247911 674000 247923
rect 675376 247911 675382 247923
rect 675434 247911 675440 247963
rect 205840 247393 205846 247445
rect 205898 247433 205904 247445
rect 205898 247405 403358 247433
rect 205898 247393 205904 247405
rect 211600 247319 211606 247371
rect 211658 247359 211664 247371
rect 211658 247331 396350 247359
rect 211658 247319 211664 247331
rect 211792 247245 211798 247297
rect 211850 247285 211856 247297
rect 211850 247257 396254 247285
rect 211850 247245 211856 247257
rect 212176 247171 212182 247223
rect 212234 247211 212240 247223
rect 212234 247183 388670 247211
rect 212234 247171 212240 247183
rect 211984 247097 211990 247149
rect 212042 247137 212048 247149
rect 212042 247109 378686 247137
rect 212042 247097 212048 247109
rect 267490 247035 267806 247063
rect 90736 246949 90742 247001
rect 90794 246989 90800 247001
rect 100240 246989 100246 247001
rect 90794 246961 100246 246989
rect 90794 246949 90800 246961
rect 100240 246949 100246 246961
rect 100298 246949 100304 247001
rect 187888 246949 187894 247001
rect 187946 246989 187952 247001
rect 201520 246989 201526 247001
rect 187946 246961 201526 246989
rect 187946 246949 187952 246961
rect 201520 246949 201526 246961
rect 201578 246949 201584 247001
rect 63280 246875 63286 246927
rect 63338 246915 63344 246927
rect 204976 246915 204982 246927
rect 63338 246887 204982 246915
rect 63338 246875 63344 246887
rect 204976 246875 204982 246887
rect 205034 246875 205040 246927
rect 56080 246801 56086 246853
rect 56138 246841 56144 246853
rect 204688 246841 204694 246853
rect 56138 246813 204694 246841
rect 56138 246801 56144 246813
rect 204688 246801 204694 246813
rect 204746 246801 204752 246853
rect 211600 246801 211606 246853
rect 211658 246841 211664 246853
rect 211658 246813 212894 246841
rect 211658 246801 211664 246813
rect 53488 246727 53494 246779
rect 53546 246767 53552 246779
rect 204784 246767 204790 246779
rect 53546 246739 204790 246767
rect 53546 246727 53552 246739
rect 204784 246727 204790 246739
rect 204842 246727 204848 246779
rect 212656 246767 212662 246779
rect 210946 246739 212662 246767
rect 56272 246653 56278 246705
rect 56330 246693 56336 246705
rect 210160 246693 210166 246705
rect 56330 246665 210166 246693
rect 56330 246653 56336 246665
rect 210160 246653 210166 246665
rect 210218 246653 210224 246705
rect 53680 246579 53686 246631
rect 53738 246619 53744 246631
rect 90736 246619 90742 246631
rect 53738 246591 90742 246619
rect 53738 246579 53744 246591
rect 90736 246579 90742 246591
rect 90794 246579 90800 246631
rect 100240 246579 100246 246631
rect 100298 246619 100304 246631
rect 210946 246619 210974 246739
rect 212656 246727 212662 246739
rect 212714 246727 212720 246779
rect 212866 246767 212894 246813
rect 228226 246813 243422 246841
rect 228226 246779 228254 246813
rect 221584 246767 221590 246779
rect 212866 246739 221590 246767
rect 221584 246727 221590 246739
rect 221642 246727 221648 246779
rect 228208 246727 228214 246779
rect 228266 246727 228272 246779
rect 229648 246727 229654 246779
rect 229706 246767 229712 246779
rect 243088 246767 243094 246779
rect 229706 246739 243094 246767
rect 229706 246727 229712 246739
rect 243088 246727 243094 246739
rect 243146 246727 243152 246779
rect 243394 246767 243422 246813
rect 267490 246779 267518 247035
rect 267778 246989 267806 247035
rect 289954 247035 311198 247063
rect 267778 246961 288446 246989
rect 270850 246813 280958 246841
rect 246160 246767 246166 246779
rect 243394 246739 246166 246767
rect 246160 246727 246166 246739
rect 246218 246727 246224 246779
rect 254032 246727 254038 246779
rect 254090 246767 254096 246779
rect 254090 246739 266750 246767
rect 254090 246727 254096 246739
rect 211120 246653 211126 246705
rect 211178 246693 211184 246705
rect 211178 246665 226142 246693
rect 211178 246653 211184 246665
rect 100298 246591 210974 246619
rect 100298 246579 100304 246591
rect 211024 246579 211030 246631
rect 211082 246619 211088 246631
rect 226000 246619 226006 246631
rect 211082 246591 226006 246619
rect 211082 246579 211088 246591
rect 226000 246579 226006 246591
rect 226058 246579 226064 246631
rect 226114 246619 226142 246665
rect 226384 246653 226390 246705
rect 226442 246693 226448 246705
rect 243376 246693 243382 246705
rect 226442 246665 243382 246693
rect 226442 246653 226448 246665
rect 243376 246653 243382 246665
rect 243434 246653 243440 246705
rect 248272 246653 248278 246705
rect 248330 246693 248336 246705
rect 266608 246693 266614 246705
rect 248330 246665 266614 246693
rect 248330 246653 248336 246665
rect 266608 246653 266614 246665
rect 266666 246653 266672 246705
rect 266722 246693 266750 246739
rect 267472 246727 267478 246779
rect 267530 246727 267536 246779
rect 269296 246727 269302 246779
rect 269354 246767 269360 246779
rect 270850 246767 270878 246813
rect 269354 246739 270878 246767
rect 280930 246767 280958 246813
rect 288418 246779 288446 246961
rect 288610 246887 289790 246915
rect 288304 246767 288310 246779
rect 280930 246739 288310 246767
rect 269354 246727 269360 246739
rect 288304 246727 288310 246739
rect 288362 246727 288368 246779
rect 288400 246727 288406 246779
rect 288458 246727 288464 246779
rect 288610 246693 288638 246887
rect 289762 246841 289790 246887
rect 289954 246841 289982 247035
rect 289762 246813 289982 246841
rect 290146 246961 310046 246989
rect 290146 246779 290174 246961
rect 291106 246887 309854 246915
rect 291106 246779 291134 246887
rect 292642 246813 309758 246841
rect 292642 246779 292670 246813
rect 309730 246779 309758 246813
rect 309826 246779 309854 246887
rect 310018 246779 310046 246961
rect 311170 246779 311198 247035
rect 326338 246887 350366 246915
rect 326338 246779 326366 246887
rect 339778 246813 348926 246841
rect 290128 246727 290134 246779
rect 290186 246727 290192 246779
rect 291088 246727 291094 246779
rect 291146 246727 291152 246779
rect 292624 246727 292630 246779
rect 292682 246727 292688 246779
rect 309712 246727 309718 246779
rect 309770 246727 309776 246779
rect 309808 246727 309814 246779
rect 309866 246727 309872 246779
rect 310000 246727 310006 246779
rect 310058 246727 310064 246779
rect 311152 246727 311158 246779
rect 311210 246727 311216 246779
rect 326320 246727 326326 246779
rect 326378 246727 326384 246779
rect 266722 246665 288638 246693
rect 290032 246653 290038 246705
rect 290090 246693 290096 246705
rect 292144 246693 292150 246705
rect 290090 246665 292150 246693
rect 290090 246653 290096 246665
rect 292144 246653 292150 246665
rect 292202 246653 292208 246705
rect 297136 246653 297142 246705
rect 297194 246693 297200 246705
rect 304624 246693 304630 246705
rect 297194 246665 304630 246693
rect 297194 246653 297200 246665
rect 304624 246653 304630 246665
rect 304682 246653 304688 246705
rect 328528 246693 328534 246705
rect 305602 246665 328534 246693
rect 247696 246619 247702 246631
rect 226114 246591 247702 246619
rect 247696 246579 247702 246591
rect 247754 246579 247760 246631
rect 247792 246579 247798 246631
rect 247850 246619 247856 246631
rect 247850 246591 267806 246619
rect 247850 246579 247856 246591
rect 53296 246505 53302 246557
rect 53354 246545 53360 246557
rect 90640 246545 90646 246557
rect 53354 246517 90646 246545
rect 53354 246505 53360 246517
rect 90640 246505 90646 246517
rect 90698 246505 90704 246557
rect 100528 246505 100534 246557
rect 100586 246545 100592 246557
rect 212272 246545 212278 246557
rect 100586 246517 212278 246545
rect 100586 246505 100592 246517
rect 212272 246505 212278 246517
rect 212330 246505 212336 246557
rect 221584 246505 221590 246557
rect 221642 246545 221648 246557
rect 229648 246545 229654 246557
rect 221642 246517 229654 246545
rect 221642 246505 221648 246517
rect 229648 246505 229654 246517
rect 229706 246505 229712 246557
rect 229936 246505 229942 246557
rect 229994 246545 230000 246557
rect 243184 246545 243190 246557
rect 229994 246517 243190 246545
rect 229994 246505 230000 246517
rect 243184 246505 243190 246517
rect 243242 246505 243248 246557
rect 267472 246545 267478 246557
rect 247810 246517 267478 246545
rect 53200 246431 53206 246483
rect 53258 246471 53264 246483
rect 53258 246443 100382 246471
rect 53258 246431 53264 246443
rect 44656 246357 44662 246409
rect 44714 246397 44720 246409
rect 100240 246397 100246 246409
rect 44714 246369 100246 246397
rect 44714 246357 44720 246369
rect 100240 246357 100246 246369
rect 100298 246357 100304 246409
rect 100354 246397 100382 246443
rect 100546 246443 205022 246471
rect 100546 246397 100574 246443
rect 100354 246369 100574 246397
rect 100624 246357 100630 246409
rect 100682 246397 100688 246409
rect 204880 246397 204886 246409
rect 100682 246369 204886 246397
rect 100682 246357 100688 246369
rect 204880 246357 204886 246369
rect 204938 246357 204944 246409
rect 204994 246397 205022 246443
rect 210544 246431 210550 246483
rect 210602 246471 210608 246483
rect 228304 246471 228310 246483
rect 210602 246443 228310 246471
rect 210602 246431 210608 246443
rect 228304 246431 228310 246443
rect 228362 246431 228368 246483
rect 228688 246431 228694 246483
rect 228746 246471 228752 246483
rect 247810 246471 247838 246517
rect 267472 246505 267478 246517
rect 267530 246505 267536 246557
rect 267778 246545 267806 246591
rect 268816 246579 268822 246631
rect 268874 246619 268880 246631
rect 280816 246619 280822 246631
rect 268874 246591 280822 246619
rect 268874 246579 268880 246591
rect 280816 246579 280822 246591
rect 280874 246579 280880 246631
rect 288400 246579 288406 246631
rect 288458 246619 288464 246631
rect 290128 246619 290134 246631
rect 288458 246591 290134 246619
rect 288458 246579 288464 246591
rect 290128 246579 290134 246591
rect 290186 246579 290192 246631
rect 290992 246579 290998 246631
rect 291050 246619 291056 246631
rect 291568 246619 291574 246631
rect 291050 246591 291574 246619
rect 291050 246579 291056 246591
rect 291568 246579 291574 246591
rect 291626 246579 291632 246631
rect 291952 246579 291958 246631
rect 292010 246619 292016 246631
rect 305602 246619 305630 246665
rect 328528 246653 328534 246665
rect 328586 246653 328592 246705
rect 329008 246653 329014 246705
rect 329066 246693 329072 246705
rect 339280 246693 339286 246705
rect 329066 246665 339286 246693
rect 329066 246653 329072 246665
rect 339280 246653 339286 246665
rect 339338 246653 339344 246705
rect 292010 246591 305630 246619
rect 292010 246579 292016 246591
rect 307984 246579 307990 246631
rect 308042 246619 308048 246631
rect 309424 246619 309430 246631
rect 308042 246591 309430 246619
rect 308042 246579 308048 246591
rect 309424 246579 309430 246591
rect 309482 246579 309488 246631
rect 324016 246579 324022 246631
rect 324074 246619 324080 246631
rect 339778 246619 339806 246813
rect 348898 246779 348926 246813
rect 350338 246779 350366 246887
rect 350434 246887 369950 246915
rect 348112 246727 348118 246779
rect 348170 246767 348176 246779
rect 348592 246767 348598 246779
rect 348170 246739 348598 246767
rect 348170 246727 348176 246739
rect 348592 246727 348598 246739
rect 348650 246727 348656 246779
rect 348880 246727 348886 246779
rect 348938 246727 348944 246779
rect 350320 246727 350326 246779
rect 350378 246727 350384 246779
rect 350434 246693 350462 246887
rect 339970 246665 350462 246693
rect 350530 246813 369854 246841
rect 324074 246591 339806 246619
rect 324074 246579 324080 246591
rect 339856 246579 339862 246631
rect 339914 246619 339920 246631
rect 339970 246619 339998 246665
rect 339914 246591 339998 246619
rect 339914 246579 339920 246591
rect 340144 246579 340150 246631
rect 340202 246619 340208 246631
rect 350128 246619 350134 246631
rect 340202 246591 350134 246619
rect 340202 246579 340208 246591
rect 350128 246579 350134 246591
rect 350186 246579 350192 246631
rect 267856 246545 267862 246557
rect 267778 246517 267862 246545
rect 267856 246505 267862 246517
rect 267914 246505 267920 246557
rect 269200 246505 269206 246557
rect 269258 246545 269264 246557
rect 287824 246545 287830 246557
rect 269258 246517 287830 246545
rect 269258 246505 269264 246517
rect 287824 246505 287830 246517
rect 287882 246505 287888 246557
rect 287920 246505 287926 246557
rect 287978 246545 287984 246557
rect 292624 246545 292630 246557
rect 287978 246517 292630 246545
rect 287978 246505 287984 246517
rect 292624 246505 292630 246517
rect 292682 246505 292688 246557
rect 297616 246505 297622 246557
rect 297674 246545 297680 246557
rect 297904 246545 297910 246557
rect 297674 246517 297910 246545
rect 297674 246505 297680 246517
rect 297904 246505 297910 246517
rect 297962 246505 297968 246557
rect 300208 246505 300214 246557
rect 300266 246545 300272 246557
rect 302320 246545 302326 246557
rect 300266 246517 302326 246545
rect 300266 246505 300272 246517
rect 302320 246505 302326 246517
rect 302378 246505 302384 246557
rect 307504 246505 307510 246557
rect 307562 246545 307568 246557
rect 307562 246517 308030 246545
rect 307562 246505 307568 246517
rect 228746 246443 247838 246471
rect 228746 246431 228752 246443
rect 248176 246431 248182 246483
rect 248234 246471 248240 246483
rect 248234 246443 267902 246471
rect 248234 246431 248240 246443
rect 204994 246369 210494 246397
rect 44752 246283 44758 246335
rect 44810 246323 44816 246335
rect 209680 246323 209686 246335
rect 44810 246295 209686 246323
rect 44810 246283 44816 246295
rect 209680 246283 209686 246295
rect 209738 246283 209744 246335
rect 60400 246209 60406 246261
rect 60458 246249 60464 246261
rect 161296 246249 161302 246261
rect 60458 246221 161302 246249
rect 60458 246209 60464 246221
rect 161296 246209 161302 246221
rect 161354 246209 161360 246261
rect 181552 246209 181558 246261
rect 181610 246249 181616 246261
rect 202576 246249 202582 246261
rect 181610 246221 202582 246249
rect 181610 246209 181616 246221
rect 202576 246209 202582 246221
rect 202634 246209 202640 246261
rect 210466 246249 210494 246369
rect 210736 246357 210742 246409
rect 210794 246397 210800 246409
rect 266512 246397 266518 246409
rect 210794 246369 266518 246397
rect 210794 246357 210800 246369
rect 266512 246357 266518 246369
rect 266570 246357 266576 246409
rect 266608 246357 266614 246409
rect 266666 246397 266672 246409
rect 267760 246397 267766 246409
rect 266666 246369 267766 246397
rect 266666 246357 266672 246369
rect 267760 246357 267766 246369
rect 267818 246357 267824 246409
rect 267874 246397 267902 246443
rect 267952 246431 267958 246483
rect 268010 246471 268016 246483
rect 288016 246471 288022 246483
rect 268010 246443 288022 246471
rect 268010 246431 268016 246443
rect 288016 246431 288022 246443
rect 288074 246431 288080 246483
rect 288304 246431 288310 246483
rect 288362 246471 288368 246483
rect 290608 246471 290614 246483
rect 288362 246443 290614 246471
rect 288362 246431 288368 246443
rect 290608 246431 290614 246443
rect 290666 246431 290672 246483
rect 308002 246471 308030 246517
rect 308080 246505 308086 246557
rect 308138 246545 308144 246557
rect 326320 246545 326326 246557
rect 308138 246517 326326 246545
rect 308138 246505 308144 246517
rect 326320 246505 326326 246517
rect 326378 246505 326384 246557
rect 328912 246505 328918 246557
rect 328970 246545 328976 246557
rect 350530 246545 350558 246813
rect 369826 246779 369854 246813
rect 369922 246779 369950 246887
rect 378658 246779 378686 247109
rect 388642 247063 388670 247183
rect 388642 247035 393374 247063
rect 393346 246779 393374 247035
rect 369808 246727 369814 246779
rect 369866 246727 369872 246779
rect 369904 246727 369910 246779
rect 369962 246727 369968 246779
rect 378640 246727 378646 246779
rect 378698 246727 378704 246779
rect 389488 246727 389494 246779
rect 389546 246767 389552 246779
rect 393040 246767 393046 246779
rect 389546 246739 393046 246767
rect 389546 246727 389552 246739
rect 393040 246727 393046 246739
rect 393098 246727 393104 246779
rect 393328 246727 393334 246779
rect 393386 246727 393392 246779
rect 352336 246653 352342 246705
rect 352394 246693 352400 246705
rect 377200 246693 377206 246705
rect 352394 246665 377206 246693
rect 352394 246653 352400 246665
rect 377200 246653 377206 246665
rect 377258 246653 377264 246705
rect 388240 246653 388246 246705
rect 388298 246693 388304 246705
rect 389008 246693 389014 246705
rect 388298 246665 389014 246693
rect 388298 246653 388304 246665
rect 389008 246653 389014 246665
rect 389066 246653 389072 246705
rect 392560 246653 392566 246705
rect 392618 246693 392624 246705
rect 393424 246693 393430 246705
rect 392618 246665 393430 246693
rect 392618 246653 392624 246665
rect 393424 246653 393430 246665
rect 393482 246653 393488 246705
rect 396226 246693 396254 247257
rect 396130 246665 396254 246693
rect 396322 246693 396350 247331
rect 403330 246779 403358 247405
rect 674032 247245 674038 247297
rect 674090 247285 674096 247297
rect 675472 247285 675478 247297
rect 674090 247257 675478 247285
rect 674090 247245 674096 247257
rect 675472 247245 675478 247257
rect 675530 247245 675536 247297
rect 403312 246727 403318 246779
rect 403370 246727 403376 246779
rect 674320 246727 674326 246779
rect 674378 246767 674384 246779
rect 675376 246767 675382 246779
rect 674378 246739 675382 246767
rect 674378 246727 674384 246739
rect 675376 246727 675382 246739
rect 675434 246727 675440 246779
rect 403792 246693 403798 246705
rect 396322 246665 403798 246693
rect 368464 246579 368470 246631
rect 368522 246619 368528 246631
rect 369040 246619 369046 246631
rect 368522 246591 369046 246619
rect 368522 246579 368528 246591
rect 369040 246579 369046 246591
rect 369098 246579 369104 246631
rect 369808 246579 369814 246631
rect 369866 246619 369872 246631
rect 370672 246619 370678 246631
rect 369866 246591 370678 246619
rect 369866 246579 369872 246591
rect 370672 246579 370678 246591
rect 370730 246579 370736 246631
rect 388528 246579 388534 246631
rect 388586 246619 388592 246631
rect 388586 246591 390014 246619
rect 388586 246579 388592 246591
rect 328970 246517 350558 246545
rect 328970 246505 328976 246517
rect 350608 246505 350614 246557
rect 350666 246545 350672 246557
rect 369424 246545 369430 246557
rect 350666 246517 369430 246545
rect 350666 246505 350672 246517
rect 369424 246505 369430 246517
rect 369482 246505 369488 246557
rect 369712 246505 369718 246557
rect 369770 246545 369776 246557
rect 389776 246545 389782 246557
rect 369770 246517 389782 246545
rect 369770 246505 369776 246517
rect 389776 246505 389782 246517
rect 389834 246505 389840 246557
rect 308002 246443 308222 246471
rect 287920 246397 287926 246409
rect 267874 246369 287926 246397
rect 287920 246357 287926 246369
rect 287978 246357 287984 246409
rect 288112 246357 288118 246409
rect 288170 246397 288176 246409
rect 308080 246397 308086 246409
rect 288170 246369 308086 246397
rect 288170 246357 288176 246369
rect 308080 246357 308086 246369
rect 308138 246357 308144 246409
rect 308194 246397 308222 246443
rect 310000 246431 310006 246483
rect 310058 246471 310064 246483
rect 347536 246471 347542 246483
rect 310058 246443 347542 246471
rect 310058 246431 310064 246443
rect 347536 246431 347542 246443
rect 347594 246431 347600 246483
rect 350320 246431 350326 246483
rect 350378 246471 350384 246483
rect 389488 246471 389494 246483
rect 350378 246443 369086 246471
rect 350378 246431 350384 246443
rect 309616 246397 309622 246409
rect 308194 246369 309622 246397
rect 309616 246357 309622 246369
rect 309674 246357 309680 246409
rect 309712 246357 309718 246409
rect 309770 246397 309776 246409
rect 368368 246397 368374 246409
rect 309770 246369 368374 246397
rect 309770 246357 309776 246369
rect 368368 246357 368374 246369
rect 368426 246357 368432 246409
rect 369058 246397 369086 246443
rect 369250 246443 389494 246471
rect 369250 246397 369278 246443
rect 389488 246431 389494 246443
rect 389546 246431 389552 246483
rect 389986 246471 390014 246591
rect 396130 246545 396158 246665
rect 403792 246653 403798 246665
rect 403850 246653 403856 246705
rect 404368 246545 404374 246557
rect 396130 246517 404374 246545
rect 404368 246505 404374 246517
rect 404426 246505 404432 246557
rect 405136 246471 405142 246483
rect 389986 246443 405142 246471
rect 405136 246431 405142 246443
rect 405194 246431 405200 246483
rect 369058 246369 369278 246397
rect 378640 246357 378646 246409
rect 378698 246397 378704 246409
rect 378698 246369 383294 246397
rect 378698 246357 378704 246369
rect 211312 246283 211318 246335
rect 211370 246323 211376 246335
rect 228208 246323 228214 246335
rect 211370 246295 228214 246323
rect 211370 246283 211376 246295
rect 228208 246283 228214 246295
rect 228266 246283 228272 246335
rect 228304 246283 228310 246335
rect 228362 246323 228368 246335
rect 229936 246323 229942 246335
rect 228362 246295 229942 246323
rect 228362 246283 228368 246295
rect 229936 246283 229942 246295
rect 229994 246283 230000 246335
rect 247696 246283 247702 246335
rect 247754 246323 247760 246335
rect 324016 246323 324022 246335
rect 247754 246295 324022 246323
rect 247754 246283 247760 246295
rect 324016 246283 324022 246295
rect 324074 246283 324080 246335
rect 327088 246283 327094 246335
rect 327146 246323 327152 246335
rect 327146 246295 329054 246323
rect 327146 246283 327152 246295
rect 211888 246249 211894 246261
rect 210466 246221 211894 246249
rect 211888 246209 211894 246221
rect 211946 246209 211952 246261
rect 222448 246209 222454 246261
rect 222506 246249 222512 246261
rect 269296 246249 269302 246261
rect 222506 246221 269302 246249
rect 222506 246209 222512 246221
rect 269296 246209 269302 246221
rect 269354 246209 269360 246261
rect 271600 246209 271606 246261
rect 271658 246249 271664 246261
rect 287344 246249 287350 246261
rect 271658 246221 287350 246249
rect 271658 246209 271664 246221
rect 287344 246209 287350 246221
rect 287402 246209 287408 246261
rect 288112 246209 288118 246261
rect 288170 246249 288176 246261
rect 307504 246249 307510 246261
rect 288170 246221 307510 246249
rect 288170 246209 288176 246221
rect 307504 246209 307510 246221
rect 307562 246209 307568 246261
rect 308176 246209 308182 246261
rect 308234 246249 308240 246261
rect 308234 246221 309758 246249
rect 308234 246209 308240 246221
rect 161392 246135 161398 246187
rect 161450 246175 161456 246187
rect 181456 246175 181462 246187
rect 161450 246147 181462 246175
rect 161450 246135 161456 246147
rect 181456 246135 181462 246147
rect 181514 246135 181520 246187
rect 226000 246135 226006 246187
rect 226058 246175 226064 246187
rect 228688 246175 228694 246187
rect 226058 246147 228694 246175
rect 226058 246135 226064 246147
rect 228688 246135 228694 246147
rect 228746 246135 228752 246187
rect 243088 246135 243094 246187
rect 243146 246175 243152 246187
rect 248272 246175 248278 246187
rect 243146 246147 248278 246175
rect 243146 246135 243152 246147
rect 248272 246135 248278 246147
rect 248330 246135 248336 246187
rect 263440 246135 263446 246187
rect 263498 246175 263504 246187
rect 277936 246175 277942 246187
rect 263498 246147 277942 246175
rect 263498 246135 263504 246147
rect 277936 246135 277942 246147
rect 277994 246135 278000 246187
rect 280816 246135 280822 246187
rect 280874 246175 280880 246187
rect 287824 246175 287830 246187
rect 280874 246147 287830 246175
rect 280874 246135 280880 246147
rect 287824 246135 287830 246147
rect 287882 246135 287888 246187
rect 288016 246135 288022 246187
rect 288074 246175 288080 246187
rect 307888 246175 307894 246187
rect 288074 246147 307894 246175
rect 288074 246135 288080 246147
rect 307888 246135 307894 246147
rect 307946 246135 307952 246187
rect 309730 246175 309758 246221
rect 309808 246209 309814 246261
rect 309866 246249 309872 246261
rect 328912 246249 328918 246261
rect 309866 246221 328918 246249
rect 309866 246209 309872 246221
rect 328912 246209 328918 246221
rect 328970 246209 328976 246261
rect 329026 246249 329054 246295
rect 339280 246283 339286 246335
rect 339338 246323 339344 246335
rect 339856 246323 339862 246335
rect 339338 246295 339862 246323
rect 339338 246283 339344 246295
rect 339856 246283 339862 246295
rect 339914 246283 339920 246335
rect 339952 246283 339958 246335
rect 340010 246323 340016 246335
rect 347248 246323 347254 246335
rect 340010 246295 347254 246323
rect 340010 246283 340016 246295
rect 347248 246283 347254 246295
rect 347306 246283 347312 246335
rect 350128 246283 350134 246335
rect 350186 246323 350192 246335
rect 350186 246295 367550 246323
rect 350186 246283 350192 246295
rect 352336 246249 352342 246261
rect 329026 246221 352342 246249
rect 352336 246209 352342 246221
rect 352394 246209 352400 246261
rect 367522 246249 367550 246295
rect 367600 246283 367606 246335
rect 367658 246323 367664 246335
rect 367658 246295 383198 246323
rect 367658 246283 367664 246295
rect 367522 246221 383102 246249
rect 383074 246187 383102 246221
rect 383170 246187 383198 246295
rect 383266 246249 383294 246369
rect 383344 246357 383350 246409
rect 383402 246397 383408 246409
rect 383584 246397 383590 246409
rect 383402 246369 383590 246397
rect 383402 246357 383408 246369
rect 383584 246357 383590 246369
rect 383642 246357 383648 246409
rect 391984 246249 391990 246261
rect 383266 246221 391990 246249
rect 391984 246209 391990 246221
rect 392042 246209 392048 246261
rect 393040 246209 393046 246261
rect 393098 246249 393104 246261
rect 409168 246249 409174 246261
rect 393098 246221 409174 246249
rect 393098 246209 393104 246221
rect 409168 246209 409174 246221
rect 409226 246209 409232 246261
rect 340144 246175 340150 246187
rect 309730 246147 340150 246175
rect 340144 246135 340150 246147
rect 340202 246135 340208 246187
rect 340240 246135 340246 246187
rect 340298 246175 340304 246187
rect 347344 246175 347350 246187
rect 340298 246147 347350 246175
rect 340298 246135 340304 246147
rect 347344 246135 347350 246147
rect 347402 246135 347408 246187
rect 347536 246135 347542 246187
rect 347594 246175 347600 246187
rect 350608 246175 350614 246187
rect 347594 246147 350614 246175
rect 347594 246135 347600 246147
rect 350608 246135 350614 246147
rect 350666 246135 350672 246187
rect 367984 246135 367990 246187
rect 368042 246175 368048 246187
rect 370192 246175 370198 246187
rect 368042 246147 370198 246175
rect 368042 246135 368048 246147
rect 370192 246135 370198 246147
rect 370250 246135 370256 246187
rect 383056 246135 383062 246187
rect 383114 246135 383120 246187
rect 383152 246135 383158 246187
rect 383210 246135 383216 246187
rect 393328 246135 393334 246187
rect 393386 246175 393392 246187
rect 403888 246175 403894 246187
rect 393386 246147 403894 246175
rect 393386 246135 393392 246147
rect 403888 246135 403894 246147
rect 403946 246135 403952 246187
rect 41296 246061 41302 246113
rect 41354 246101 41360 246113
rect 43312 246101 43318 246113
rect 41354 246073 43318 246101
rect 41354 246061 41360 246073
rect 43312 246061 43318 246073
rect 43370 246101 43376 246113
rect 504016 246101 504022 246113
rect 43370 246073 504022 246101
rect 43370 246061 43376 246073
rect 504016 246061 504022 246073
rect 504074 246061 504080 246113
rect 43408 245987 43414 246039
rect 43466 246027 43472 246039
rect 43466 245999 339998 246027
rect 43466 245987 43472 245999
rect 243184 245913 243190 245965
rect 243242 245953 243248 245965
rect 248176 245953 248182 245965
rect 243242 245925 248182 245953
rect 243242 245913 243248 245925
rect 248176 245913 248182 245925
rect 248234 245913 248240 245965
rect 263824 245913 263830 245965
rect 263882 245953 263888 245965
rect 263882 245925 277886 245953
rect 263882 245913 263888 245925
rect 181360 245839 181366 245891
rect 181418 245839 181424 245891
rect 246160 245839 246166 245891
rect 246218 245879 246224 245891
rect 248368 245879 248374 245891
rect 246218 245851 248374 245879
rect 246218 245839 246224 245851
rect 248368 245839 248374 245851
rect 248426 245839 248432 245891
rect 263056 245839 263062 245891
rect 263114 245879 263120 245891
rect 277744 245879 277750 245891
rect 263114 245851 277750 245879
rect 263114 245839 263120 245851
rect 277744 245839 277750 245851
rect 277802 245839 277808 245891
rect 277858 245879 277886 245925
rect 277936 245913 277942 245965
rect 277994 245953 278000 245965
rect 339856 245953 339862 245965
rect 277994 245925 339862 245953
rect 277994 245913 278000 245925
rect 339856 245913 339862 245925
rect 339914 245913 339920 245965
rect 339970 245953 339998 245999
rect 347344 245987 347350 246039
rect 347402 246027 347408 246039
rect 509776 246027 509782 246039
rect 347402 245999 509782 246027
rect 347402 245987 347408 245999
rect 509776 245987 509782 245999
rect 509834 245987 509840 246039
rect 340240 245953 340246 245965
rect 339970 245925 340246 245953
rect 340240 245913 340246 245925
rect 340298 245913 340304 245965
rect 347248 245913 347254 245965
rect 347306 245953 347312 245965
rect 368080 245953 368086 245965
rect 347306 245925 368086 245953
rect 347306 245913 347312 245925
rect 368080 245913 368086 245925
rect 368138 245913 368144 245965
rect 368368 245913 368374 245965
rect 368426 245953 368432 245965
rect 369712 245953 369718 245965
rect 368426 245925 369718 245953
rect 368426 245913 368432 245925
rect 369712 245913 369718 245925
rect 369770 245913 369776 245965
rect 391984 245913 391990 245965
rect 392042 245953 392048 245965
rect 400912 245953 400918 245965
rect 392042 245925 400918 245953
rect 392042 245913 392048 245925
rect 400912 245913 400918 245925
rect 400970 245913 400976 245965
rect 367504 245879 367510 245891
rect 277858 245851 367510 245879
rect 367504 245839 367510 245851
rect 367562 245839 367568 245891
rect 383152 245839 383158 245891
rect 383210 245879 383216 245891
rect 401488 245879 401494 245891
rect 383210 245851 401494 245879
rect 383210 245839 383216 245851
rect 401488 245839 401494 245851
rect 401546 245839 401552 245891
rect 181378 245521 181406 245839
rect 251824 245765 251830 245817
rect 251882 245805 251888 245817
rect 356656 245805 356662 245817
rect 251882 245777 356662 245805
rect 251882 245765 251888 245777
rect 356656 245765 356662 245777
rect 356714 245765 356720 245817
rect 368560 245765 368566 245817
rect 368618 245805 368624 245817
rect 388720 245805 388726 245817
rect 368618 245777 388726 245805
rect 368618 245765 368624 245777
rect 388720 245765 388726 245777
rect 388778 245765 388784 245817
rect 202576 245691 202582 245743
rect 202634 245731 202640 245743
rect 213136 245731 213142 245743
rect 202634 245703 213142 245731
rect 202634 245691 202640 245703
rect 213136 245691 213142 245703
rect 213194 245691 213200 245743
rect 216880 245691 216886 245743
rect 216938 245731 216944 245743
rect 228208 245731 228214 245743
rect 216938 245703 228214 245731
rect 216938 245691 216944 245703
rect 228208 245691 228214 245703
rect 228266 245691 228272 245743
rect 243376 245691 243382 245743
rect 243434 245731 243440 245743
rect 254032 245731 254038 245743
rect 243434 245703 254038 245731
rect 243434 245691 243440 245703
rect 254032 245691 254038 245703
rect 254090 245691 254096 245743
rect 254128 245691 254134 245743
rect 254186 245731 254192 245743
rect 358000 245731 358006 245743
rect 254186 245703 358006 245731
rect 254186 245691 254192 245703
rect 358000 245691 358006 245703
rect 358058 245691 358064 245743
rect 383056 245691 383062 245743
rect 383114 245731 383120 245743
rect 392944 245731 392950 245743
rect 383114 245703 392950 245731
rect 383114 245691 383120 245703
rect 392944 245691 392950 245703
rect 393002 245691 393008 245743
rect 266512 245617 266518 245669
rect 266570 245657 266576 245669
rect 269200 245657 269206 245669
rect 266570 245629 269206 245657
rect 266570 245617 266576 245629
rect 269200 245617 269206 245629
rect 269258 245617 269264 245669
rect 277744 245617 277750 245669
rect 277802 245657 277808 245669
rect 369232 245657 369238 245669
rect 277802 245629 369238 245657
rect 277802 245617 277808 245629
rect 369232 245617 369238 245629
rect 369290 245617 369296 245669
rect 227536 245543 227542 245595
rect 227594 245583 227600 245595
rect 247984 245583 247990 245595
rect 227594 245555 247990 245583
rect 227594 245543 227600 245555
rect 247984 245543 247990 245555
rect 248042 245543 248048 245595
rect 262672 245543 262678 245595
rect 262730 245583 262736 245595
rect 369808 245583 369814 245595
rect 262730 245555 369814 245583
rect 262730 245543 262736 245555
rect 369808 245543 369814 245555
rect 369866 245543 369872 245595
rect 181360 245469 181366 245521
rect 181418 245469 181424 245521
rect 253360 245469 253366 245521
rect 253418 245509 253424 245521
rect 357616 245509 357622 245521
rect 253418 245481 357622 245509
rect 253418 245469 253424 245481
rect 357616 245469 357622 245481
rect 357674 245469 357680 245521
rect 202192 245395 202198 245447
rect 202250 245435 202256 245447
rect 222448 245435 222454 245447
rect 202250 245407 222454 245435
rect 202250 245395 202256 245407
rect 222448 245395 222454 245407
rect 222506 245395 222512 245447
rect 252400 245395 252406 245447
rect 252458 245435 252464 245447
rect 357136 245435 357142 245447
rect 252458 245407 357142 245435
rect 252458 245395 252464 245407
rect 357136 245395 357142 245407
rect 357194 245395 357200 245447
rect 168592 245321 168598 245373
rect 168650 245361 168656 245373
rect 181264 245361 181270 245373
rect 168650 245333 181270 245361
rect 168650 245321 168656 245333
rect 181264 245321 181270 245333
rect 181322 245321 181328 245373
rect 261808 245321 261814 245373
rect 261866 245361 261872 245373
rect 372016 245361 372022 245373
rect 261866 245333 372022 245361
rect 261866 245321 261872 245333
rect 372016 245321 372022 245333
rect 372074 245321 372080 245373
rect 260848 245247 260854 245299
rect 260906 245287 260912 245299
rect 374032 245287 374038 245299
rect 260906 245259 374038 245287
rect 260906 245247 260912 245259
rect 374032 245247 374038 245259
rect 374090 245247 374096 245299
rect 211792 245173 211798 245225
rect 211850 245213 211856 245225
rect 247600 245213 247606 245225
rect 211850 245185 247606 245213
rect 211850 245173 211856 245185
rect 247600 245173 247606 245185
rect 247658 245173 247664 245225
rect 261232 245173 261238 245225
rect 261290 245213 261296 245225
rect 372880 245213 372886 245225
rect 261290 245185 372886 245213
rect 261290 245173 261296 245185
rect 372880 245173 372886 245185
rect 372938 245173 372944 245225
rect 389776 245173 389782 245225
rect 389834 245213 389840 245225
rect 407056 245213 407062 245225
rect 389834 245185 407062 245213
rect 389834 245173 389840 245185
rect 407056 245173 407062 245185
rect 407114 245173 407120 245225
rect 211984 245099 211990 245151
rect 212042 245139 212048 245151
rect 227440 245139 227446 245151
rect 212042 245111 227446 245139
rect 212042 245099 212048 245111
rect 227440 245099 227446 245111
rect 227498 245099 227504 245151
rect 260368 245099 260374 245151
rect 260426 245139 260432 245151
rect 375760 245139 375766 245151
rect 260426 245111 375766 245139
rect 260426 245099 260432 245111
rect 375760 245099 375766 245111
rect 375818 245099 375824 245151
rect 227056 245025 227062 245077
rect 227114 245065 227120 245077
rect 227920 245065 227926 245077
rect 227114 245037 227926 245065
rect 227114 245025 227120 245037
rect 227920 245025 227926 245037
rect 227978 245025 227984 245077
rect 246448 245025 246454 245077
rect 246506 245065 246512 245077
rect 248080 245065 248086 245077
rect 246506 245037 248086 245065
rect 246506 245025 246512 245037
rect 248080 245025 248086 245037
rect 248138 245025 248144 245077
rect 260464 245025 260470 245077
rect 260522 245065 260528 245077
rect 374608 245065 374614 245077
rect 260522 245037 374614 245065
rect 260522 245025 260528 245037
rect 374608 245025 374614 245037
rect 374666 245025 374672 245077
rect 42352 244951 42358 245003
rect 42410 244991 42416 245003
rect 214192 244991 214198 245003
rect 42410 244963 214198 244991
rect 42410 244951 42416 244963
rect 214192 244951 214198 244963
rect 214250 244951 214256 245003
rect 216496 244951 216502 245003
rect 216554 244991 216560 245003
rect 358480 244991 358486 245003
rect 216554 244963 358486 244991
rect 216554 244951 216560 244963
rect 358480 244951 358486 244963
rect 358538 244951 358544 245003
rect 210160 244877 210166 244929
rect 210218 244917 210224 244929
rect 214096 244917 214102 244929
rect 210218 244889 214102 244917
rect 210218 244877 210224 244889
rect 214096 244877 214102 244889
rect 214154 244877 214160 244929
rect 247696 244877 247702 244929
rect 247754 244917 247760 244929
rect 268240 244917 268246 244929
rect 247754 244889 268246 244917
rect 247754 244877 247760 244889
rect 268240 244877 268246 244889
rect 268298 244877 268304 244929
rect 292336 244917 292342 244929
rect 268354 244889 292342 244917
rect 97936 244803 97942 244855
rect 97994 244843 98000 244855
rect 97994 244815 109406 244843
rect 97994 244803 98000 244815
rect 109378 244769 109406 244815
rect 193264 244803 193270 244855
rect 193322 244843 193328 244855
rect 193322 244815 195902 244843
rect 193322 244803 193328 244815
rect 144592 244769 144598 244781
rect 109378 244741 144598 244769
rect 144592 244729 144598 244741
rect 144650 244729 144656 244781
rect 195874 244769 195902 244815
rect 209680 244803 209686 244855
rect 209738 244843 209744 244855
rect 213520 244843 213526 244855
rect 209738 244815 213526 244843
rect 209738 244803 209744 244815
rect 213520 244803 213526 244815
rect 213578 244803 213584 244855
rect 247984 244803 247990 244855
rect 248042 244843 248048 244855
rect 268354 244843 268382 244889
rect 292336 244877 292342 244889
rect 292394 244877 292400 244929
rect 299536 244877 299542 244929
rect 299594 244917 299600 244929
rect 307696 244917 307702 244929
rect 299594 244889 307702 244917
rect 299594 244877 299600 244889
rect 307696 244877 307702 244889
rect 307754 244877 307760 244929
rect 307792 244877 307798 244929
rect 307850 244917 307856 244929
rect 309136 244917 309142 244929
rect 307850 244889 309142 244917
rect 307850 244877 307856 244889
rect 309136 244877 309142 244889
rect 309194 244877 309200 244929
rect 309616 244877 309622 244929
rect 309674 244917 309680 244929
rect 328240 244917 328246 244929
rect 309674 244889 328246 244917
rect 309674 244877 309680 244889
rect 328240 244877 328246 244889
rect 328298 244877 328304 244929
rect 328528 244877 328534 244929
rect 328586 244917 328592 244929
rect 368464 244917 368470 244929
rect 328586 244889 368470 244917
rect 328586 244877 328592 244889
rect 368464 244877 368470 244889
rect 368522 244877 368528 244929
rect 389776 244917 389782 244929
rect 368578 244889 389782 244917
rect 308080 244843 308086 244855
rect 248042 244815 268382 244843
rect 269314 244815 308086 244843
rect 248042 244803 248048 244815
rect 198928 244769 198934 244781
rect 195874 244741 198934 244769
rect 198928 244729 198934 244741
rect 198986 244729 198992 244781
rect 227632 244729 227638 244781
rect 227690 244769 227696 244781
rect 228112 244769 228118 244781
rect 227690 244741 228118 244769
rect 227690 244729 227696 244741
rect 228112 244729 228118 244741
rect 228170 244729 228176 244781
rect 248080 244729 248086 244781
rect 248138 244769 248144 244781
rect 267856 244769 267862 244781
rect 248138 244741 267862 244769
rect 248138 244729 248144 244741
rect 267856 244729 267862 244741
rect 267914 244729 267920 244781
rect 268816 244769 268822 244781
rect 268162 244741 268822 244769
rect 102544 244655 102550 244707
rect 102602 244695 102608 244707
rect 142960 244695 142966 244707
rect 102602 244667 142966 244695
rect 102602 244655 102608 244667
rect 142960 244655 142966 244667
rect 143018 244655 143024 244707
rect 259216 244655 259222 244707
rect 259274 244695 259280 244707
rect 268162 244695 268190 244741
rect 268816 244729 268822 244741
rect 268874 244729 268880 244781
rect 259274 244667 268190 244695
rect 259274 244655 259280 244667
rect 268240 244655 268246 244707
rect 268298 244695 268304 244707
rect 269314 244695 269342 244815
rect 308080 244803 308086 244815
rect 308138 244803 308144 244855
rect 328624 244843 328630 244855
rect 309058 244815 328630 244843
rect 278032 244729 278038 244781
rect 278090 244769 278096 244781
rect 298000 244769 298006 244781
rect 278090 244741 298006 244769
rect 278090 244729 278096 244741
rect 298000 244729 298006 244741
rect 298058 244729 298064 244781
rect 298096 244729 298102 244781
rect 298154 244769 298160 244781
rect 309058 244769 309086 244815
rect 328624 244803 328630 244815
rect 328682 244803 328688 244855
rect 348208 244803 348214 244855
rect 348266 244843 348272 244855
rect 368578 244843 368606 244889
rect 389776 244877 389782 244889
rect 389834 244877 389840 244929
rect 348266 244815 368606 244843
rect 348266 244803 348272 244815
rect 368848 244803 368854 244855
rect 368906 244843 368912 244855
rect 388528 244843 388534 244855
rect 368906 244815 388534 244843
rect 368906 244803 368912 244815
rect 388528 244803 388534 244815
rect 388586 244803 388592 244855
rect 608176 244803 608182 244855
rect 608234 244843 608240 244855
rect 613456 244843 613462 244855
rect 608234 244815 613462 244843
rect 608234 244803 608240 244815
rect 613456 244803 613462 244815
rect 613514 244803 613520 244855
rect 298154 244741 309086 244769
rect 298154 244729 298160 244741
rect 309136 244729 309142 244781
rect 309194 244769 309200 244781
rect 327952 244769 327958 244781
rect 309194 244741 327958 244769
rect 309194 244729 309200 244741
rect 327952 244729 327958 244741
rect 328010 244729 328016 244781
rect 328048 244729 328054 244781
rect 328106 244769 328112 244781
rect 338608 244769 338614 244781
rect 328106 244741 338614 244769
rect 328106 244729 328112 244741
rect 338608 244729 338614 244741
rect 338666 244729 338672 244781
rect 268298 244667 269342 244695
rect 268298 244655 268304 244667
rect 277744 244655 277750 244707
rect 277802 244695 277808 244707
rect 318160 244695 318166 244707
rect 277802 244667 318166 244695
rect 277802 244655 277808 244667
rect 318160 244655 318166 244667
rect 318218 244655 318224 244707
rect 326800 244655 326806 244707
rect 326858 244695 326864 244707
rect 329008 244695 329014 244707
rect 326858 244667 329014 244695
rect 326858 244655 326864 244667
rect 329008 244655 329014 244667
rect 329066 244655 329072 244707
rect 389776 244655 389782 244707
rect 389834 244695 389840 244707
rect 404368 244695 404374 244707
rect 389834 244667 404374 244695
rect 389834 244655 389840 244667
rect 404368 244655 404374 244667
rect 404426 244655 404432 244707
rect 138160 244581 138166 244633
rect 138218 244621 138224 244633
rect 205744 244621 205750 244633
rect 138218 244593 205750 244621
rect 138218 244581 138224 244593
rect 205744 244581 205750 244593
rect 205802 244581 205808 244633
rect 235120 244581 235126 244633
rect 235178 244621 235184 244633
rect 267184 244621 267190 244633
rect 235178 244593 267190 244621
rect 235178 244581 235184 244593
rect 267184 244581 267190 244593
rect 267242 244581 267248 244633
rect 277840 244581 277846 244633
rect 277898 244621 277904 244633
rect 318256 244621 318262 244633
rect 277898 244593 318262 244621
rect 277898 244581 277904 244593
rect 318256 244581 318262 244593
rect 318314 244581 318320 244633
rect 135280 244507 135286 244559
rect 135338 244547 135344 244559
rect 206992 244547 206998 244559
rect 135338 244519 206998 244547
rect 135338 244507 135344 244519
rect 206992 244507 206998 244519
rect 207050 244507 207056 244559
rect 242224 244507 242230 244559
rect 242282 244547 242288 244559
rect 257776 244547 257782 244559
rect 242282 244519 257782 244547
rect 242282 244507 242288 244519
rect 257776 244507 257782 244519
rect 257834 244507 257840 244559
rect 262000 244507 262006 244559
rect 262058 244547 262064 244559
rect 338128 244547 338134 244559
rect 262058 244519 338134 244547
rect 262058 244507 262064 244519
rect 338128 244507 338134 244519
rect 338186 244507 338192 244559
rect 132400 244433 132406 244485
rect 132458 244473 132464 244485
rect 205456 244473 205462 244485
rect 132458 244445 205462 244473
rect 132458 244433 132464 244445
rect 205456 244433 205462 244445
rect 205514 244433 205520 244485
rect 277936 244433 277942 244485
rect 277994 244473 278000 244485
rect 328048 244473 328054 244485
rect 277994 244445 328054 244473
rect 277994 244433 278000 244445
rect 328048 244433 328054 244445
rect 328106 244433 328112 244485
rect 42064 244359 42070 244411
rect 42122 244399 42128 244411
rect 42544 244399 42550 244411
rect 42122 244371 42550 244399
rect 42122 244359 42128 244371
rect 42544 244359 42550 244371
rect 42602 244359 42608 244411
rect 126640 244359 126646 244411
rect 126698 244399 126704 244411
rect 205264 244399 205270 244411
rect 126698 244371 205270 244399
rect 126698 244359 126704 244371
rect 205264 244359 205270 244371
rect 205322 244359 205328 244411
rect 260560 244359 260566 244411
rect 260618 244399 260624 244411
rect 308752 244399 308758 244411
rect 260618 244371 308758 244399
rect 260618 244359 260624 244371
rect 308752 244359 308758 244371
rect 308810 244359 308816 244411
rect 123760 244285 123766 244337
rect 123818 244325 123824 244337
rect 205072 244325 205078 244337
rect 123818 244297 205078 244325
rect 123818 244285 123824 244297
rect 205072 244285 205078 244297
rect 205130 244285 205136 244337
rect 258928 244285 258934 244337
rect 258986 244325 258992 244337
rect 336688 244325 336694 244337
rect 258986 244297 336694 244325
rect 258986 244285 258992 244297
rect 336688 244285 336694 244297
rect 336746 244285 336752 244337
rect 674800 244285 674806 244337
rect 674858 244325 674864 244337
rect 675280 244325 675286 244337
rect 674858 244297 675286 244325
rect 674858 244285 674864 244297
rect 675280 244285 675286 244297
rect 675338 244285 675344 244337
rect 120880 244211 120886 244263
rect 120938 244251 120944 244263
rect 205648 244251 205654 244263
rect 120938 244223 205654 244251
rect 120938 244211 120944 244223
rect 205648 244211 205654 244223
rect 205706 244211 205712 244263
rect 257200 244211 257206 244263
rect 257258 244251 257264 244263
rect 335920 244251 335926 244263
rect 257258 244223 335926 244251
rect 257258 244211 257264 244223
rect 335920 244211 335926 244223
rect 335978 244211 335984 244263
rect 383056 244211 383062 244263
rect 383114 244251 383120 244263
rect 383440 244251 383446 244263
rect 383114 244223 383446 244251
rect 383114 244211 383120 244223
rect 383440 244211 383446 244223
rect 383498 244211 383504 244263
rect 118000 244137 118006 244189
rect 118058 244177 118064 244189
rect 204496 244177 204502 244189
rect 118058 244149 204502 244177
rect 118058 244137 118064 244149
rect 204496 244137 204502 244149
rect 204554 244137 204560 244189
rect 211504 244137 211510 244189
rect 211562 244177 211568 244189
rect 267856 244177 267862 244189
rect 211562 244149 267862 244177
rect 211562 244137 211568 244149
rect 267856 244137 267862 244149
rect 267914 244137 267920 244189
rect 267952 244137 267958 244189
rect 268010 244177 268016 244189
rect 297904 244177 297910 244189
rect 268010 244149 297910 244177
rect 268010 244137 268016 244149
rect 297904 244137 297910 244149
rect 297962 244137 297968 244189
rect 298000 244137 298006 244189
rect 298058 244177 298064 244189
rect 309904 244177 309910 244189
rect 298058 244149 309910 244177
rect 298058 244137 298064 244149
rect 309904 244137 309910 244149
rect 309962 244137 309968 244189
rect 312400 244137 312406 244189
rect 312458 244177 312464 244189
rect 368752 244177 368758 244189
rect 312458 244149 368758 244177
rect 312458 244137 312464 244149
rect 368752 244137 368758 244149
rect 368810 244137 368816 244189
rect 112240 244063 112246 244115
rect 112298 244103 112304 244115
rect 206416 244103 206422 244115
rect 112298 244075 206422 244103
rect 112298 244063 112304 244075
rect 206416 244063 206422 244075
rect 206474 244063 206480 244115
rect 251344 244063 251350 244115
rect 251402 244103 251408 244115
rect 356272 244103 356278 244115
rect 251402 244075 356278 244103
rect 251402 244063 251408 244075
rect 356272 244063 356278 244075
rect 356330 244063 356336 244115
rect 109360 243989 109366 244041
rect 109418 244029 109424 244041
rect 206224 244029 206230 244041
rect 109418 244001 206230 244029
rect 109418 243989 109424 244001
rect 206224 243989 206230 244001
rect 206282 243989 206288 244041
rect 249616 243989 249622 244041
rect 249674 244029 249680 244041
rect 355792 244029 355798 244041
rect 249674 244001 355798 244029
rect 249674 243989 249680 244001
rect 355792 243989 355798 244001
rect 355850 243989 355856 244041
rect 106480 243915 106486 243967
rect 106538 243955 106544 243967
rect 204592 243955 204598 243967
rect 106538 243927 204598 243955
rect 106538 243915 106544 243927
rect 204592 243915 204598 243927
rect 204650 243915 204656 243967
rect 257776 243915 257782 243967
rect 257834 243955 257840 243967
rect 352144 243955 352150 243967
rect 257834 243927 352150 243955
rect 257834 243915 257840 243927
rect 352144 243915 352150 243927
rect 352202 243915 352208 243967
rect 103600 243841 103606 243893
rect 103658 243881 103664 243893
rect 206608 243881 206614 243893
rect 103658 243853 206614 243881
rect 103658 243841 103664 243853
rect 206608 243841 206614 243853
rect 206666 243841 206672 243893
rect 243280 243841 243286 243893
rect 243338 243881 243344 243893
rect 352624 243881 352630 243893
rect 243338 243853 352630 243881
rect 243338 243841 243344 243853
rect 352624 243841 352630 243853
rect 352682 243841 352688 243893
rect 100144 243767 100150 243819
rect 100202 243807 100208 243819
rect 206512 243807 206518 243819
rect 100202 243779 206518 243807
rect 100202 243767 100208 243779
rect 206512 243767 206518 243779
rect 206570 243767 206576 243819
rect 244720 243767 244726 243819
rect 244778 243807 244784 243819
rect 353584 243807 353590 243819
rect 244778 243779 353590 243807
rect 244778 243767 244784 243779
rect 353584 243767 353590 243779
rect 353642 243767 353648 243819
rect 94960 243693 94966 243745
rect 95018 243733 95024 243745
rect 206320 243733 206326 243745
rect 95018 243705 206326 243733
rect 95018 243693 95024 243705
rect 206320 243693 206326 243705
rect 206378 243693 206384 243745
rect 246352 243693 246358 243745
rect 246410 243733 246416 243745
rect 299488 243733 299494 243745
rect 246410 243705 299494 243733
rect 246410 243693 246416 243705
rect 299488 243693 299494 243705
rect 299546 243693 299552 243745
rect 299650 243705 299774 243733
rect 92080 243619 92086 243671
rect 92138 243659 92144 243671
rect 206032 243659 206038 243671
rect 92138 243631 206038 243659
rect 92138 243619 92144 243631
rect 206032 243619 206038 243631
rect 206090 243619 206096 243671
rect 247312 243619 247318 243671
rect 247370 243659 247376 243671
rect 299650 243659 299678 243705
rect 247370 243631 299678 243659
rect 299746 243659 299774 243705
rect 307696 243693 307702 243745
rect 307754 243733 307760 243745
rect 354352 243733 354358 243745
rect 307754 243705 354358 243733
rect 307754 243693 307760 243705
rect 354352 243693 354358 243705
rect 354410 243693 354416 243745
rect 354832 243659 354838 243671
rect 299746 243631 354838 243659
rect 247370 243619 247376 243631
rect 354832 243619 354838 243631
rect 354890 243619 354896 243671
rect 86320 243545 86326 243597
rect 86378 243585 86384 243597
rect 206704 243585 206710 243597
rect 86378 243557 206710 243585
rect 86378 243545 86384 243557
rect 206704 243545 206710 243557
rect 206762 243545 206768 243597
rect 237136 243545 237142 243597
rect 237194 243585 237200 243597
rect 349936 243585 349942 243597
rect 237194 243557 349942 243585
rect 237194 243545 237200 243557
rect 349936 243545 349942 243557
rect 349994 243545 350000 243597
rect 80560 243471 80566 243523
rect 80618 243511 80624 243523
rect 206896 243511 206902 243523
rect 80618 243483 206902 243511
rect 80618 243471 80624 243483
rect 206896 243471 206902 243483
rect 206954 243471 206960 243523
rect 240496 243471 240502 243523
rect 240554 243511 240560 243523
rect 296656 243511 296662 243523
rect 240554 243483 296662 243511
rect 240554 243471 240560 243483
rect 296656 243471 296662 243483
rect 296714 243471 296720 243523
rect 297136 243471 297142 243523
rect 297194 243511 297200 243523
rect 351472 243511 351478 243523
rect 297194 243483 351478 243511
rect 297194 243471 297200 243483
rect 351472 243471 351478 243483
rect 351530 243471 351536 243523
rect 77680 243397 77686 243449
rect 77738 243437 77744 243449
rect 205168 243437 205174 243449
rect 77738 243409 205174 243437
rect 77738 243397 77744 243409
rect 205168 243397 205174 243409
rect 205226 243397 205232 243449
rect 230608 243397 230614 243449
rect 230666 243437 230672 243449
rect 346672 243437 346678 243449
rect 230666 243409 346678 243437
rect 230666 243397 230672 243409
rect 346672 243397 346678 243409
rect 346730 243397 346736 243449
rect 69040 243323 69046 243375
rect 69098 243363 69104 243375
rect 206128 243363 206134 243375
rect 69098 243335 206134 243363
rect 69098 243323 69104 243335
rect 206128 243323 206134 243335
rect 206186 243323 206192 243375
rect 227824 243323 227830 243375
rect 227882 243363 227888 243375
rect 296656 243363 296662 243375
rect 227882 243335 296662 243363
rect 227882 243323 227888 243335
rect 296656 243323 296662 243335
rect 296714 243323 296720 243375
rect 297136 243323 297142 243375
rect 297194 243363 297200 243375
rect 345520 243363 345526 243375
rect 297194 243335 345526 243363
rect 297194 243323 297200 243335
rect 345520 243323 345526 243335
rect 345578 243323 345584 243375
rect 235600 243249 235606 243301
rect 235658 243289 235664 243301
rect 266128 243289 266134 243301
rect 235658 243261 266134 243289
rect 235658 243249 235664 243261
rect 266128 243249 266134 243261
rect 266186 243249 266192 243301
rect 270160 243249 270166 243301
rect 270218 243289 270224 243301
rect 296752 243289 296758 243301
rect 270218 243261 296758 243289
rect 270218 243249 270224 243261
rect 296752 243249 296758 243261
rect 296810 243249 296816 243301
rect 297232 243249 297238 243301
rect 297290 243289 297296 243301
rect 323056 243289 323062 243301
rect 297290 243261 323062 243289
rect 297290 243249 297296 243261
rect 323056 243249 323062 243261
rect 323114 243249 323120 243301
rect 282160 243175 282166 243227
rect 282218 243215 282224 243227
rect 296656 243215 296662 243227
rect 282218 243187 296662 243215
rect 282218 243175 282224 243187
rect 296656 243175 296662 243187
rect 296714 243175 296720 243227
rect 296944 243175 296950 243227
rect 297002 243215 297008 243227
rect 308368 243215 308374 243227
rect 297002 243187 308374 243215
rect 297002 243175 297008 243187
rect 308368 243175 308374 243187
rect 308426 243175 308432 243227
rect 308752 243175 308758 243227
rect 308810 243215 308816 243227
rect 337264 243215 337270 243227
rect 308810 243187 337270 243215
rect 308810 243175 308816 243187
rect 337264 243175 337270 243187
rect 337322 243175 337328 243227
rect 266992 243101 266998 243153
rect 267050 243141 267056 243153
rect 279760 243141 279766 243153
rect 267050 243113 279766 243141
rect 267050 243101 267056 243113
rect 279760 243101 279766 243113
rect 279818 243101 279824 243153
rect 279952 243101 279958 243153
rect 280010 243141 280016 243153
rect 296752 243141 296758 243153
rect 280010 243113 296758 243141
rect 280010 243101 280016 243113
rect 296752 243101 296758 243113
rect 296810 243101 296816 243153
rect 309424 243141 309430 243153
rect 296866 243113 309430 243141
rect 267088 243027 267094 243079
rect 267146 243067 267152 243079
rect 277840 243067 277846 243079
rect 267146 243039 277846 243067
rect 267146 243027 267152 243039
rect 277840 243027 277846 243039
rect 277898 243027 277904 243079
rect 287344 243027 287350 243079
rect 287402 243067 287408 243079
rect 296866 243067 296894 243113
rect 309424 243101 309430 243113
rect 309482 243101 309488 243153
rect 318160 243101 318166 243153
rect 318218 243141 318224 243153
rect 339568 243141 339574 243153
rect 318218 243113 339574 243141
rect 318218 243101 318224 243113
rect 339568 243101 339574 243113
rect 339626 243101 339632 243153
rect 287402 243039 296894 243067
rect 287402 243027 287408 243039
rect 318256 243027 318262 243079
rect 318314 243067 318320 243079
rect 340336 243067 340342 243079
rect 318314 243039 340342 243067
rect 318314 243027 318320 243039
rect 340336 243027 340342 243039
rect 340394 243027 340400 243079
rect 267472 242953 267478 243005
rect 267530 242993 267536 243005
rect 304144 242993 304150 243005
rect 267530 242965 304150 242993
rect 267530 242953 267536 242965
rect 304144 242953 304150 242965
rect 304202 242953 304208 243005
rect 675184 242953 675190 243005
rect 675242 242993 675248 243005
rect 675376 242993 675382 243005
rect 675242 242965 675382 242993
rect 675242 242953 675248 242965
rect 675376 242953 675382 242965
rect 675434 242953 675440 243005
rect 265072 242879 265078 242931
rect 265130 242919 265136 242931
rect 277744 242919 277750 242931
rect 265130 242891 277750 242919
rect 265130 242879 265136 242891
rect 277744 242879 277750 242891
rect 277802 242879 277808 242931
rect 284656 242879 284662 242931
rect 284714 242919 284720 242931
rect 298096 242919 298102 242931
rect 284714 242891 298102 242919
rect 284714 242879 284720 242891
rect 298096 242879 298102 242891
rect 298154 242879 298160 242931
rect 263728 242805 263734 242857
rect 263786 242845 263792 242857
rect 277936 242845 277942 242857
rect 263786 242817 277942 242845
rect 263786 242805 263792 242817
rect 277936 242805 277942 242817
rect 277994 242805 278000 242857
rect 301264 242845 301270 242857
rect 293698 242817 301270 242845
rect 270832 242731 270838 242783
rect 270890 242771 270896 242783
rect 293392 242771 293398 242783
rect 270890 242743 293398 242771
rect 270890 242731 270896 242743
rect 293392 242731 293398 242743
rect 293450 242731 293456 242783
rect 293488 242731 293494 242783
rect 293546 242771 293552 242783
rect 293698 242771 293726 242817
rect 301264 242805 301270 242817
rect 301322 242805 301328 242857
rect 293546 242743 293726 242771
rect 293546 242731 293552 242743
rect 293872 242731 293878 242783
rect 293930 242771 293936 242783
rect 293930 242743 297854 242771
rect 293930 242731 293936 242743
rect 297826 242697 297854 242743
rect 297904 242731 297910 242783
rect 297962 242771 297968 242783
rect 316432 242771 316438 242783
rect 297962 242743 316438 242771
rect 297962 242731 297968 242743
rect 316432 242731 316438 242743
rect 316490 242731 316496 242783
rect 320848 242697 320854 242709
rect 297826 242669 320854 242697
rect 320848 242657 320854 242669
rect 320906 242657 320912 242709
rect 264880 242583 264886 242635
rect 264938 242623 264944 242635
rect 278032 242623 278038 242635
rect 264938 242595 278038 242623
rect 264938 242583 264944 242595
rect 278032 242583 278038 242595
rect 278090 242583 278096 242635
rect 284752 242583 284758 242635
rect 284810 242623 284816 242635
rect 317104 242623 317110 242635
rect 284810 242595 317110 242623
rect 284810 242583 284816 242595
rect 317104 242583 317110 242595
rect 317162 242583 317168 242635
rect 267856 242509 267862 242561
rect 267914 242549 267920 242561
rect 287440 242549 287446 242561
rect 267914 242521 287446 242549
rect 267914 242509 267920 242521
rect 287440 242509 287446 242521
rect 287498 242509 287504 242561
rect 287536 242509 287542 242561
rect 287594 242549 287600 242561
rect 293488 242549 293494 242561
rect 287594 242521 293494 242549
rect 287594 242509 287600 242521
rect 293488 242509 293494 242521
rect 293546 242509 293552 242561
rect 297904 242509 297910 242561
rect 297962 242549 297968 242561
rect 319120 242549 319126 242561
rect 297962 242521 319126 242549
rect 297962 242509 297968 242521
rect 319120 242509 319126 242521
rect 319178 242509 319184 242561
rect 269680 242435 269686 242487
rect 269738 242475 269744 242487
rect 269738 242447 290750 242475
rect 269738 242435 269744 242447
rect 274480 242361 274486 242413
rect 274538 242401 274544 242413
rect 289456 242401 289462 242413
rect 274538 242373 289462 242401
rect 274538 242361 274544 242373
rect 289456 242361 289462 242373
rect 289514 242361 289520 242413
rect 269200 242287 269206 242339
rect 269258 242327 269264 242339
rect 287536 242327 287542 242339
rect 269258 242299 287542 242327
rect 269258 242287 269264 242299
rect 287536 242287 287542 242299
rect 287594 242287 287600 242339
rect 290722 242327 290750 242447
rect 293968 242435 293974 242487
rect 294026 242475 294032 242487
rect 297520 242475 297526 242487
rect 294026 242447 297526 242475
rect 294026 242435 294032 242447
rect 297520 242435 297526 242447
rect 297578 242435 297584 242487
rect 298096 242435 298102 242487
rect 298154 242475 298160 242487
rect 317968 242475 317974 242487
rect 298154 242447 317974 242475
rect 298154 242435 298160 242447
rect 317968 242435 317974 242447
rect 318026 242435 318032 242487
rect 290800 242361 290806 242413
rect 290858 242401 290864 242413
rect 321328 242401 321334 242413
rect 290858 242373 321334 242401
rect 290858 242361 290864 242373
rect 321328 242361 321334 242373
rect 321386 242361 321392 242413
rect 675088 242361 675094 242413
rect 675146 242401 675152 242413
rect 675376 242401 675382 242413
rect 675146 242373 675382 242401
rect 675146 242361 675152 242373
rect 675376 242361 675382 242373
rect 675434 242361 675440 242413
rect 299248 242327 299254 242339
rect 290722 242299 299254 242327
rect 299248 242287 299254 242299
rect 299306 242287 299312 242339
rect 299632 242287 299638 242339
rect 299690 242327 299696 242339
rect 323440 242327 323446 242339
rect 299690 242299 323446 242327
rect 299690 242287 299696 242299
rect 323440 242287 323446 242299
rect 323498 242287 323504 242339
rect 141136 242213 141142 242265
rect 141194 242253 141200 242265
rect 161104 242253 161110 242265
rect 141194 242225 161110 242253
rect 141194 242213 141200 242225
rect 161104 242213 161110 242225
rect 161162 242213 161168 242265
rect 288976 242213 288982 242265
rect 289034 242253 289040 242265
rect 292336 242253 292342 242265
rect 289034 242225 292342 242253
rect 289034 242213 289040 242225
rect 292336 242213 292342 242225
rect 292394 242213 292400 242265
rect 292432 242213 292438 242265
rect 292490 242253 292496 242265
rect 321904 242253 321910 242265
rect 292490 242225 321910 242253
rect 292490 242213 292496 242225
rect 321904 242213 321910 242225
rect 321962 242213 321968 242265
rect 270448 242139 270454 242191
rect 270506 242179 270512 242191
rect 297616 242179 297622 242191
rect 270506 242151 297622 242179
rect 270506 242139 270512 242151
rect 297616 242139 297622 242151
rect 297674 242139 297680 242191
rect 298000 242139 298006 242191
rect 298058 242179 298064 242191
rect 305392 242179 305398 242191
rect 298058 242151 305398 242179
rect 298058 242139 298064 242151
rect 305392 242139 305398 242151
rect 305450 242139 305456 242191
rect 317968 242139 317974 242191
rect 318026 242179 318032 242191
rect 335632 242179 335638 242191
rect 318026 242151 335638 242179
rect 318026 242139 318032 242151
rect 335632 242139 335638 242151
rect 335690 242139 335696 242191
rect 40048 242065 40054 242117
rect 40106 242105 40112 242117
rect 42352 242105 42358 242117
rect 40106 242077 42358 242105
rect 40106 242065 40112 242077
rect 42352 242065 42358 242077
rect 42410 242065 42416 242117
rect 157936 242065 157942 242117
rect 157994 242105 158000 242117
rect 157994 242077 161246 242105
rect 157994 242065 158000 242077
rect 40144 241991 40150 242043
rect 40202 242031 40208 242043
rect 43120 242031 43126 242043
rect 40202 242003 43126 242031
rect 40202 241991 40208 242003
rect 43120 241991 43126 242003
rect 43178 241991 43184 242043
rect 161104 241991 161110 242043
rect 161162 241991 161168 242043
rect 161218 242031 161246 242077
rect 284272 242065 284278 242117
rect 284330 242105 284336 242117
rect 297904 242105 297910 242117
rect 284330 242077 297910 242105
rect 284330 242065 284336 242077
rect 297904 242065 297910 242077
rect 297962 242065 297968 242117
rect 298192 242065 298198 242117
rect 298250 242105 298256 242117
rect 316912 242105 316918 242117
rect 298250 242077 316918 242105
rect 298250 242065 298256 242077
rect 316912 242065 316918 242077
rect 316970 242065 316976 242117
rect 319600 242065 319606 242117
rect 319658 242105 319664 242117
rect 333424 242105 333430 242117
rect 319658 242077 333430 242105
rect 319658 242065 319664 242077
rect 333424 242065 333430 242077
rect 333482 242065 333488 242117
rect 177040 242031 177046 242043
rect 161218 242003 177046 242031
rect 177040 241991 177046 242003
rect 177098 241991 177104 242043
rect 205840 242031 205846 242043
rect 191458 242003 205846 242031
rect 37360 241917 37366 241969
rect 37418 241957 37424 241969
rect 42928 241957 42934 241969
rect 37418 241929 42934 241957
rect 37418 241917 37424 241929
rect 42928 241917 42934 241929
rect 42986 241917 42992 241969
rect 44560 241917 44566 241969
rect 44618 241957 44624 241969
rect 141136 241957 141142 241969
rect 44618 241929 141142 241957
rect 44618 241917 44624 241929
rect 141136 241917 141142 241929
rect 141194 241917 141200 241969
rect 161122 241957 161150 241991
rect 191458 241957 191486 242003
rect 205840 241991 205846 242003
rect 205898 241991 205904 242043
rect 292240 242031 292246 242043
rect 289090 242003 292246 242031
rect 288976 241957 288982 241969
rect 161122 241929 191486 241957
rect 241858 241929 288982 241957
rect 238480 241843 238486 241895
rect 238538 241883 238544 241895
rect 241858 241883 241886 241929
rect 288976 241917 288982 241929
rect 289034 241917 289040 241969
rect 238538 241855 241886 241883
rect 238538 241843 238544 241855
rect 250288 241843 250294 241895
rect 250346 241883 250352 241895
rect 273040 241883 273046 241895
rect 250346 241855 273046 241883
rect 250346 241843 250352 241855
rect 273040 241843 273046 241855
rect 273098 241843 273104 241895
rect 273136 241843 273142 241895
rect 273194 241883 273200 241895
rect 281872 241883 281878 241895
rect 273194 241855 281878 241883
rect 273194 241843 273200 241855
rect 281872 241843 281878 241855
rect 281930 241843 281936 241895
rect 283408 241843 283414 241895
rect 283466 241883 283472 241895
rect 289090 241883 289118 242003
rect 292240 241991 292246 242003
rect 292298 241991 292304 242043
rect 293584 241991 293590 242043
rect 293642 242031 293648 242043
rect 299632 242031 299638 242043
rect 293642 242003 299638 242031
rect 293642 241991 293648 242003
rect 299632 241991 299638 242003
rect 299690 241991 299696 242043
rect 290512 241917 290518 241969
rect 290570 241957 290576 241969
rect 291568 241957 291574 241969
rect 290570 241929 291574 241957
rect 290570 241917 290576 241929
rect 291568 241917 291574 241929
rect 291626 241917 291632 241969
rect 292336 241917 292342 241969
rect 292394 241957 292400 241969
rect 350512 241957 350518 241969
rect 292394 241929 350518 241957
rect 292394 241917 292400 241929
rect 350512 241917 350518 241929
rect 350570 241917 350576 241969
rect 360112 241917 360118 241969
rect 360170 241957 360176 241969
rect 371824 241957 371830 241969
rect 360170 241929 371830 241957
rect 360170 241917 360176 241929
rect 371824 241917 371830 241929
rect 371882 241917 371888 241969
rect 283466 241855 289118 241883
rect 283466 241843 283472 241855
rect 289168 241843 289174 241895
rect 289226 241883 289232 241895
rect 299728 241883 299734 241895
rect 289226 241855 299734 241883
rect 289226 241843 289232 241855
rect 299728 241843 299734 241855
rect 299786 241843 299792 241895
rect 306736 241843 306742 241895
rect 306794 241883 306800 241895
rect 309136 241883 309142 241895
rect 306794 241855 309142 241883
rect 306794 241843 306800 241855
rect 309136 241843 309142 241855
rect 309194 241843 309200 241895
rect 314224 241843 314230 241895
rect 314282 241883 314288 241895
rect 329968 241883 329974 241895
rect 314282 241855 329974 241883
rect 314282 241843 314288 241855
rect 329968 241843 329974 241855
rect 330026 241843 330032 241895
rect 338320 241843 338326 241895
rect 338378 241883 338384 241895
rect 378352 241883 378358 241895
rect 338378 241855 378358 241883
rect 338378 241843 338384 241855
rect 378352 241843 378358 241855
rect 378410 241843 378416 241895
rect 395824 241883 395830 241895
rect 378466 241855 395830 241883
rect 217552 241769 217558 241821
rect 217610 241809 217616 241821
rect 234736 241809 234742 241821
rect 217610 241781 234742 241809
rect 217610 241769 217616 241781
rect 234736 241769 234742 241781
rect 234794 241769 234800 241821
rect 248560 241769 248566 241821
rect 248618 241809 248624 241821
rect 273904 241809 273910 241821
rect 248618 241781 273910 241809
rect 248618 241769 248624 241781
rect 273904 241769 273910 241781
rect 273962 241769 273968 241821
rect 274000 241769 274006 241821
rect 274058 241809 274064 241821
rect 287056 241809 287062 241821
rect 274058 241781 287062 241809
rect 274058 241769 274064 241781
rect 287056 241769 287062 241781
rect 287114 241769 287120 241821
rect 290512 241809 290518 241821
rect 287170 241781 290518 241809
rect 219280 241695 219286 241747
rect 219338 241735 219344 241747
rect 233968 241735 233974 241747
rect 219338 241707 233974 241735
rect 219338 241695 219344 241707
rect 233968 241695 233974 241707
rect 234026 241695 234032 241747
rect 255088 241695 255094 241747
rect 255146 241735 255152 241747
rect 255146 241707 274046 241735
rect 255146 241695 255152 241707
rect 215440 241621 215446 241673
rect 215498 241661 215504 241673
rect 272944 241661 272950 241673
rect 215498 241633 272950 241661
rect 215498 241621 215504 241633
rect 272944 241621 272950 241633
rect 273002 241621 273008 241673
rect 273040 241621 273046 241673
rect 273098 241661 273104 241673
rect 273808 241661 273814 241673
rect 273098 241633 273814 241661
rect 273098 241621 273104 241633
rect 273808 241621 273814 241633
rect 273866 241621 273872 241673
rect 274018 241661 274046 241707
rect 274096 241695 274102 241747
rect 274154 241735 274160 241747
rect 287170 241735 287198 241781
rect 290512 241769 290518 241781
rect 290570 241769 290576 241821
rect 290608 241769 290614 241821
rect 290666 241809 290672 241821
rect 290666 241781 298238 241809
rect 290666 241769 290672 241781
rect 274154 241707 287198 241735
rect 274154 241695 274160 241707
rect 287344 241695 287350 241747
rect 287402 241735 287408 241747
rect 298096 241735 298102 241747
rect 287402 241707 298102 241735
rect 287402 241695 287408 241707
rect 298096 241695 298102 241707
rect 298154 241695 298160 241747
rect 289168 241661 289174 241673
rect 274018 241633 289174 241661
rect 289168 241621 289174 241633
rect 289226 241621 289232 241673
rect 289360 241621 289366 241673
rect 289418 241661 289424 241673
rect 296464 241661 296470 241673
rect 289418 241633 296470 241661
rect 289418 241621 289424 241633
rect 296464 241621 296470 241633
rect 296522 241621 296528 241673
rect 298210 241661 298238 241781
rect 307600 241769 307606 241821
rect 307658 241809 307664 241821
rect 309808 241809 309814 241821
rect 307658 241781 309814 241809
rect 307658 241769 307664 241781
rect 309808 241769 309814 241781
rect 309866 241769 309872 241821
rect 314416 241809 314422 241821
rect 312130 241781 314422 241809
rect 305584 241695 305590 241747
rect 305642 241735 305648 241747
rect 308464 241735 308470 241747
rect 305642 241707 308470 241735
rect 305642 241695 305648 241707
rect 308464 241695 308470 241707
rect 308522 241695 308528 241747
rect 312130 241661 312158 241781
rect 314416 241769 314422 241781
rect 314474 241769 314480 241821
rect 315184 241769 315190 241821
rect 315242 241809 315248 241821
rect 374416 241809 374422 241821
rect 315242 241781 374422 241809
rect 315242 241769 315248 241781
rect 374416 241769 374422 241781
rect 374474 241769 374480 241821
rect 378466 241809 378494 241855
rect 395824 241843 395830 241855
rect 395882 241843 395888 241895
rect 376930 241781 378494 241809
rect 328144 241735 328150 241747
rect 298210 241633 312158 241661
rect 314338 241707 328150 241735
rect 220432 241547 220438 241599
rect 220490 241587 220496 241599
rect 233392 241587 233398 241599
rect 220490 241559 233398 241587
rect 220490 241547 220496 241559
rect 233392 241547 233398 241559
rect 233450 241547 233456 241599
rect 237712 241547 237718 241599
rect 237770 241587 237776 241599
rect 261616 241587 261622 241599
rect 237770 241559 261622 241587
rect 237770 241547 237776 241559
rect 261616 241547 261622 241559
rect 261674 241547 261680 241599
rect 262000 241547 262006 241599
rect 262058 241587 262064 241599
rect 314338 241587 314366 241707
rect 328144 241695 328150 241707
rect 328202 241695 328208 241747
rect 328240 241695 328246 241747
rect 328298 241735 328304 241747
rect 339760 241735 339766 241747
rect 328298 241707 339766 241735
rect 328298 241695 328304 241707
rect 339760 241695 339766 241707
rect 339818 241695 339824 241747
rect 339856 241695 339862 241747
rect 339914 241735 339920 241747
rect 360112 241735 360118 241747
rect 339914 241707 360118 241735
rect 339914 241695 339920 241707
rect 360112 241695 360118 241707
rect 360170 241695 360176 241747
rect 314416 241621 314422 241673
rect 314474 241661 314480 241673
rect 316048 241661 316054 241673
rect 314474 241633 316054 241661
rect 314474 241621 314480 241633
rect 316048 241621 316054 241633
rect 316106 241621 316112 241673
rect 316624 241621 316630 241673
rect 316682 241661 316688 241673
rect 375088 241661 375094 241673
rect 316682 241633 375094 241661
rect 316682 241621 316688 241633
rect 375088 241621 375094 241633
rect 375146 241621 375152 241673
rect 325168 241587 325174 241599
rect 262058 241559 314366 241587
rect 314434 241559 325174 241587
rect 262058 241547 262064 241559
rect 223216 241473 223222 241525
rect 223274 241513 223280 241525
rect 232144 241513 232150 241525
rect 223274 241485 232150 241513
rect 223274 241473 223280 241485
rect 232144 241473 232150 241485
rect 232202 241473 232208 241525
rect 236944 241473 236950 241525
rect 237002 241513 237008 241525
rect 263344 241513 263350 241525
rect 237002 241485 263350 241513
rect 237002 241473 237008 241485
rect 263344 241473 263350 241485
rect 263402 241473 263408 241525
rect 264304 241473 264310 241525
rect 264362 241513 264368 241525
rect 271984 241513 271990 241525
rect 264362 241485 271990 241513
rect 264362 241473 264368 241485
rect 271984 241473 271990 241485
rect 272042 241473 272048 241525
rect 277936 241473 277942 241525
rect 277994 241513 278000 241525
rect 314224 241513 314230 241525
rect 277994 241485 314230 241513
rect 277994 241473 278000 241485
rect 314224 241473 314230 241485
rect 314282 241473 314288 241525
rect 213904 241399 213910 241451
rect 213962 241439 213968 241451
rect 229168 241439 229174 241451
rect 213962 241411 229174 241439
rect 213962 241399 213968 241411
rect 229168 241399 229174 241411
rect 229226 241399 229232 241451
rect 252784 241399 252790 241451
rect 252842 241439 252848 241451
rect 314434 241439 314462 241559
rect 325168 241547 325174 241559
rect 325226 241547 325232 241599
rect 325264 241547 325270 241599
rect 325322 241587 325328 241599
rect 328240 241587 328246 241599
rect 325322 241559 328246 241587
rect 325322 241547 325328 241559
rect 328240 241547 328246 241559
rect 328298 241547 328304 241599
rect 331504 241547 331510 241599
rect 331562 241587 331568 241599
rect 331562 241559 339134 241587
rect 331562 241547 331568 241559
rect 336496 241513 336502 241525
rect 318370 241485 336502 241513
rect 252842 241411 314462 241439
rect 252842 241399 252848 241411
rect 314512 241399 314518 241451
rect 314570 241439 314576 241451
rect 318370 241439 318398 241485
rect 336496 241473 336502 241485
rect 336554 241473 336560 241525
rect 339106 241513 339134 241559
rect 339184 241547 339190 241599
rect 339242 241587 339248 241599
rect 356560 241587 356566 241599
rect 339242 241559 356566 241587
rect 339242 241547 339248 241559
rect 356560 241547 356566 241559
rect 356618 241547 356624 241599
rect 361936 241547 361942 241599
rect 361994 241587 362000 241599
rect 373936 241587 373942 241599
rect 361994 241559 373942 241587
rect 361994 241547 362000 241559
rect 373936 241547 373942 241559
rect 373994 241547 374000 241599
rect 359344 241513 359350 241525
rect 339106 241485 359350 241513
rect 359344 241473 359350 241485
rect 359402 241473 359408 241525
rect 360976 241473 360982 241525
rect 361034 241513 361040 241525
rect 376930 241513 376958 241781
rect 379216 241769 379222 241821
rect 379274 241809 379280 241821
rect 409264 241809 409270 241821
rect 379274 241781 409270 241809
rect 379274 241769 379280 241781
rect 409264 241769 409270 241781
rect 409322 241769 409328 241821
rect 377008 241695 377014 241747
rect 377066 241735 377072 241747
rect 404944 241735 404950 241747
rect 377066 241707 404950 241735
rect 377066 241695 377072 241707
rect 404944 241695 404950 241707
rect 405002 241695 405008 241747
rect 379600 241621 379606 241673
rect 379658 241661 379664 241673
rect 409936 241661 409942 241673
rect 379658 241633 409942 241661
rect 379658 241621 379664 241633
rect 409936 241621 409942 241633
rect 409994 241621 410000 241673
rect 674224 241547 674230 241599
rect 674282 241587 674288 241599
rect 675472 241587 675478 241599
rect 674282 241559 675478 241587
rect 674282 241547 674288 241559
rect 675472 241547 675478 241559
rect 675530 241547 675536 241599
rect 361034 241485 376958 241513
rect 361034 241473 361040 241485
rect 380080 241473 380086 241525
rect 380138 241513 380144 241525
rect 383536 241513 383542 241525
rect 380138 241485 383542 241513
rect 380138 241473 380144 241485
rect 383536 241473 383542 241485
rect 383594 241473 383600 241525
rect 383632 241473 383638 241525
rect 383690 241513 383696 241525
rect 385552 241513 385558 241525
rect 383690 241485 385558 241513
rect 383690 241473 383696 241485
rect 385552 241473 385558 241485
rect 385610 241473 385616 241525
rect 329584 241439 329590 241451
rect 314570 241411 318398 241439
rect 318466 241411 329590 241439
rect 314570 241399 314576 241411
rect 277744 241325 277750 241377
rect 277802 241365 277808 241377
rect 314608 241365 314614 241377
rect 277802 241337 314614 241365
rect 277802 241325 277808 241337
rect 314608 241325 314614 241337
rect 314666 241325 314672 241377
rect 317776 241325 317782 241377
rect 317834 241365 317840 241377
rect 318466 241365 318494 241411
rect 329584 241399 329590 241411
rect 329642 241399 329648 241451
rect 333712 241399 333718 241451
rect 333770 241439 333776 241451
rect 362896 241439 362902 241451
rect 333770 241411 362902 241439
rect 333770 241399 333776 241411
rect 362896 241399 362902 241411
rect 362954 241399 362960 241451
rect 363184 241399 363190 241451
rect 363242 241439 363248 241451
rect 400144 241439 400150 241451
rect 363242 241411 400150 241439
rect 363242 241399 363248 241411
rect 400144 241399 400150 241411
rect 400202 241399 400208 241451
rect 317834 241337 318494 241365
rect 317834 241325 317840 241337
rect 327376 241325 327382 241377
rect 327434 241365 327440 241377
rect 332944 241365 332950 241377
rect 327434 241337 332950 241365
rect 327434 241325 327440 241337
rect 332944 241325 332950 241337
rect 333002 241325 333008 241377
rect 333328 241325 333334 241377
rect 333386 241365 333392 241377
rect 363280 241365 363286 241377
rect 333386 241337 363286 241365
rect 333386 241325 333392 241337
rect 363280 241325 363286 241337
rect 363338 241325 363344 241377
rect 364144 241325 364150 241377
rect 364202 241365 364208 241377
rect 401872 241365 401878 241377
rect 364202 241337 401878 241365
rect 364202 241325 364208 241337
rect 401872 241325 401878 241337
rect 401930 241325 401936 241377
rect 277840 241251 277846 241303
rect 277898 241291 277904 241303
rect 277898 241263 317534 241291
rect 277898 241251 277904 241263
rect 224080 241177 224086 241229
rect 224138 241217 224144 241229
rect 231760 241217 231766 241229
rect 224138 241189 231766 241217
rect 224138 241177 224144 241189
rect 231760 241177 231766 241189
rect 231818 241177 231824 241229
rect 233296 241177 233302 241229
rect 233354 241217 233360 241229
rect 238672 241217 238678 241229
rect 233354 241189 238678 241217
rect 233354 241177 233360 241189
rect 238672 241177 238678 241189
rect 238730 241177 238736 241229
rect 255952 241177 255958 241229
rect 256010 241217 256016 241229
rect 310480 241217 310486 241229
rect 256010 241189 310486 241217
rect 256010 241177 256016 241189
rect 310480 241177 310486 241189
rect 310538 241177 310544 241229
rect 317506 241217 317534 241263
rect 317872 241251 317878 241303
rect 317930 241291 317936 241303
rect 330160 241291 330166 241303
rect 317930 241263 330166 241291
rect 317930 241251 317936 241263
rect 330160 241251 330166 241263
rect 330218 241251 330224 241303
rect 331024 241251 331030 241303
rect 331082 241291 331088 241303
rect 358288 241291 358294 241303
rect 331082 241263 358294 241291
rect 331082 241251 331088 241263
rect 358288 241251 358294 241263
rect 358346 241251 358352 241303
rect 362032 241251 362038 241303
rect 362090 241291 362096 241303
rect 373552 241291 373558 241303
rect 362090 241263 373558 241291
rect 362090 241251 362096 241263
rect 373552 241251 373558 241263
rect 373610 241251 373616 241303
rect 373936 241251 373942 241303
rect 373994 241291 374000 241303
rect 397456 241291 397462 241303
rect 373994 241263 397462 241291
rect 373994 241251 374000 241263
rect 397456 241251 397462 241263
rect 397514 241251 397520 241303
rect 331696 241217 331702 241229
rect 317506 241189 331702 241217
rect 331696 241177 331702 241189
rect 331754 241177 331760 241229
rect 363760 241177 363766 241229
rect 363818 241217 363824 241229
rect 400720 241217 400726 241229
rect 363818 241189 400726 241217
rect 363818 241177 363824 241189
rect 400720 241177 400726 241189
rect 400778 241177 400784 241229
rect 225232 241103 225238 241155
rect 225290 241143 225296 241155
rect 231184 241143 231190 241155
rect 225290 241115 231190 241143
rect 225290 241103 225296 241115
rect 231184 241103 231190 241115
rect 231242 241103 231248 241155
rect 250672 241143 250678 241155
rect 237586 241115 250678 241143
rect 222544 241029 222550 241081
rect 222602 241069 222608 241081
rect 232528 241069 232534 241081
rect 222602 241041 232534 241069
rect 222602 241029 222608 241041
rect 232528 241029 232534 241041
rect 232586 241029 232592 241081
rect 216688 240955 216694 241007
rect 216746 240995 216752 241007
rect 236176 240995 236182 241007
rect 216746 240967 236182 240995
rect 216746 240955 216752 240967
rect 236176 240955 236182 240967
rect 236234 240955 236240 241007
rect 227344 240881 227350 240933
rect 227402 240921 227408 240933
rect 230320 240921 230326 240933
rect 227402 240893 230326 240921
rect 227402 240881 227408 240893
rect 230320 240881 230326 240893
rect 230378 240881 230384 240933
rect 212752 240807 212758 240859
rect 212810 240847 212816 240859
rect 233200 240847 233206 240859
rect 212810 240819 233206 240847
rect 212810 240807 212816 240819
rect 233200 240807 233206 240819
rect 233258 240807 233264 240859
rect 219280 240733 219286 240785
rect 219338 240773 219344 240785
rect 237586 240773 237614 241115
rect 250672 241103 250678 241115
rect 250730 241103 250736 241155
rect 254992 241103 254998 241155
rect 255050 241143 255056 241155
rect 314512 241143 314518 241155
rect 255050 241115 314518 241143
rect 255050 241103 255056 241115
rect 314512 241103 314518 241115
rect 314570 241103 314576 241155
rect 314608 241103 314614 241155
rect 314666 241143 314672 241155
rect 332752 241143 332758 241155
rect 314666 241115 332758 241143
rect 314666 241103 314672 241115
rect 332752 241103 332758 241115
rect 332810 241103 332816 241155
rect 364240 241103 364246 241155
rect 364298 241143 364304 241155
rect 402736 241143 402742 241155
rect 364298 241115 402742 241143
rect 364298 241103 364304 241115
rect 402736 241103 402742 241115
rect 402794 241103 402800 241155
rect 249808 241069 249814 241081
rect 219338 240745 237614 240773
rect 237682 241041 249814 241069
rect 219338 240733 219344 240745
rect 41776 240585 41782 240637
rect 41834 240585 41840 240637
rect 219664 240585 219670 240637
rect 219722 240625 219728 240637
rect 237682 240625 237710 241041
rect 249808 241029 249814 241041
rect 249866 241029 249872 241081
rect 254224 241029 254230 241081
rect 254282 241069 254288 241081
rect 337840 241069 337846 241081
rect 254282 241041 337846 241069
rect 254282 241029 254288 241041
rect 337840 241029 337846 241041
rect 337898 241029 337904 241081
rect 362896 241029 362902 241081
rect 362954 241069 362960 241081
rect 364336 241069 364342 241081
rect 362954 241041 364342 241069
rect 362954 241029 362960 241041
rect 364336 241029 364342 241041
rect 364394 241029 364400 241081
rect 373552 241029 373558 241081
rect 373610 241069 373616 241081
rect 398416 241069 398422 241081
rect 373610 241041 398422 241069
rect 373610 241029 373616 241041
rect 398416 241029 398422 241041
rect 398474 241029 398480 241081
rect 244432 240955 244438 241007
rect 244490 240995 244496 241007
rect 326896 240995 326902 241007
rect 244490 240967 326902 240995
rect 244490 240955 244496 240967
rect 326896 240955 326902 240967
rect 326954 240955 326960 241007
rect 326992 240955 326998 241007
rect 327050 240995 327056 241007
rect 338320 240995 338326 241007
rect 327050 240967 338326 240995
rect 327050 240955 327056 240967
rect 338320 240955 338326 240967
rect 338378 240955 338384 241007
rect 362416 240955 362422 241007
rect 362474 240995 362480 241007
rect 398992 240995 398998 241007
rect 362474 240967 398998 240995
rect 362474 240955 362480 240967
rect 398992 240955 398998 240967
rect 399050 240955 399056 241007
rect 237904 240881 237910 240933
rect 237962 240921 237968 240933
rect 252880 240921 252886 240933
rect 237962 240893 252886 240921
rect 237962 240881 237968 240893
rect 252880 240881 252886 240893
rect 252938 240881 252944 240933
rect 253744 240881 253750 240933
rect 253802 240921 253808 240933
rect 339376 240921 339382 240933
rect 253802 240893 339382 240921
rect 253802 240881 253808 240893
rect 339376 240881 339382 240893
rect 339434 240881 339440 240933
rect 339472 240881 339478 240933
rect 339530 240921 339536 240933
rect 362224 240921 362230 240933
rect 339530 240893 362230 240921
rect 339530 240881 339536 240893
rect 362224 240881 362230 240893
rect 362282 240881 362288 240933
rect 365968 240881 365974 240933
rect 366026 240921 366032 240933
rect 406096 240921 406102 240933
rect 366026 240893 406102 240921
rect 366026 240881 366032 240893
rect 406096 240881 406102 240893
rect 406154 240881 406160 240933
rect 237808 240807 237814 240859
rect 237866 240847 237872 240859
rect 252016 240847 252022 240859
rect 237866 240819 252022 240847
rect 237866 240807 237872 240819
rect 252016 240807 252022 240819
rect 252074 240807 252080 240859
rect 252304 240807 252310 240859
rect 252362 240847 252368 240859
rect 342640 240847 342646 240859
rect 252362 240819 342646 240847
rect 252362 240807 252368 240819
rect 342640 240807 342646 240819
rect 342698 240807 342704 240859
rect 366352 240807 366358 240859
rect 366410 240847 366416 240859
rect 407152 240847 407158 240859
rect 366410 240819 407158 240847
rect 366410 240807 366416 240819
rect 407152 240807 407158 240819
rect 407210 240807 407216 240859
rect 251536 240733 251542 240785
rect 251594 240773 251600 240785
rect 344176 240773 344182 240785
rect 251594 240745 344182 240773
rect 251594 240733 251600 240745
rect 344176 240733 344182 240745
rect 344234 240733 344240 240785
rect 365008 240733 365014 240785
rect 365066 240773 365072 240785
rect 404464 240773 404470 240785
rect 365066 240745 404470 240773
rect 365066 240733 365072 240745
rect 404464 240733 404470 240745
rect 404522 240733 404528 240785
rect 249808 240659 249814 240711
rect 249866 240699 249872 240711
rect 347440 240699 347446 240711
rect 249866 240671 347446 240699
rect 249866 240659 249872 240671
rect 347440 240659 347446 240671
rect 347498 240659 347504 240711
rect 367216 240659 367222 240711
rect 367274 240699 367280 240711
rect 408880 240699 408886 240711
rect 367274 240671 408886 240699
rect 367274 240659 367280 240671
rect 408880 240659 408886 240671
rect 408938 240659 408944 240711
rect 219722 240597 237710 240625
rect 219722 240585 219728 240597
rect 250576 240585 250582 240637
rect 250634 240625 250640 240637
rect 345712 240625 345718 240637
rect 250634 240597 345718 240625
rect 250634 240585 250640 240597
rect 345712 240585 345718 240597
rect 345770 240585 345776 240637
rect 364624 240585 364630 240637
rect 364682 240625 364688 240637
rect 403408 240625 403414 240637
rect 364682 240597 403414 240625
rect 364682 240585 364688 240597
rect 403408 240585 403414 240597
rect 403466 240585 403472 240637
rect 41794 240415 41822 240585
rect 220624 240511 220630 240563
rect 220682 240551 220688 240563
rect 247888 240551 247894 240563
rect 220682 240523 247894 240551
rect 220682 240511 220688 240523
rect 247888 240511 247894 240523
rect 247946 240511 247952 240563
rect 248368 240511 248374 240563
rect 248426 240551 248432 240563
rect 350416 240551 350422 240563
rect 248426 240523 350422 240551
rect 248426 240511 248432 240523
rect 350416 240511 350422 240523
rect 350474 240511 350480 240563
rect 365392 240511 365398 240563
rect 365450 240551 365456 240563
rect 405232 240551 405238 240563
rect 365450 240523 405238 240551
rect 365450 240511 365456 240523
rect 405232 240511 405238 240523
rect 405290 240511 405296 240563
rect 674992 240511 674998 240563
rect 675050 240551 675056 240563
rect 675472 240551 675478 240563
rect 675050 240523 675478 240551
rect 675050 240511 675056 240523
rect 675472 240511 675478 240523
rect 675530 240511 675536 240563
rect 144592 240437 144598 240489
rect 144650 240477 144656 240489
rect 162736 240477 162742 240489
rect 144650 240449 162742 240477
rect 144650 240437 144656 240449
rect 162736 240437 162742 240449
rect 162794 240437 162800 240489
rect 220240 240437 220246 240489
rect 220298 240477 220304 240489
rect 248656 240477 248662 240489
rect 220298 240449 248662 240477
rect 220298 240437 220304 240449
rect 248656 240437 248662 240449
rect 248714 240437 248720 240489
rect 249328 240437 249334 240489
rect 249386 240477 249392 240489
rect 349168 240477 349174 240489
rect 249386 240449 349174 240477
rect 249386 240437 249392 240449
rect 349168 240437 349174 240449
rect 349226 240437 349232 240489
rect 366448 240437 366454 240489
rect 366506 240477 366512 240489
rect 407728 240477 407734 240489
rect 366506 240449 407734 240477
rect 366506 240437 366512 240449
rect 407728 240437 407734 240449
rect 407786 240437 407792 240489
rect 41776 240363 41782 240415
rect 41834 240363 41840 240415
rect 218512 240363 218518 240415
rect 218570 240403 218576 240415
rect 237808 240403 237814 240415
rect 218570 240375 237814 240403
rect 218570 240363 218576 240375
rect 237808 240363 237814 240375
rect 237866 240363 237872 240415
rect 238960 240363 238966 240415
rect 239018 240403 239024 240415
rect 263920 240403 263926 240415
rect 239018 240375 263926 240403
rect 239018 240363 239024 240375
rect 263920 240363 263926 240375
rect 263978 240363 263984 240415
rect 275728 240363 275734 240415
rect 275786 240403 275792 240415
rect 283024 240403 283030 240415
rect 275786 240375 283030 240403
rect 275786 240363 275792 240375
rect 283024 240363 283030 240375
rect 283082 240363 283088 240415
rect 313360 240363 313366 240415
rect 313418 240403 313424 240415
rect 370288 240403 370294 240415
rect 313418 240375 370294 240403
rect 313418 240363 313424 240375
rect 370288 240363 370294 240375
rect 370346 240363 370352 240415
rect 378256 240363 378262 240415
rect 378314 240403 378320 240415
rect 408208 240403 408214 240415
rect 378314 240375 408214 240403
rect 378314 240363 378320 240375
rect 408208 240363 408214 240375
rect 408266 240363 408272 240415
rect 237328 240289 237334 240341
rect 237386 240329 237392 240341
rect 262192 240329 262198 240341
rect 237386 240301 262198 240329
rect 237386 240289 237392 240301
rect 262192 240289 262198 240301
rect 262250 240289 262256 240341
rect 262288 240289 262294 240341
rect 262346 240329 262352 240341
rect 277936 240329 277942 240341
rect 262346 240301 277942 240329
rect 262346 240289 262352 240301
rect 277936 240289 277942 240301
rect 277994 240289 278000 240341
rect 278032 240289 278038 240341
rect 278090 240329 278096 240341
rect 288400 240329 288406 240341
rect 278090 240301 288406 240329
rect 278090 240289 278096 240301
rect 288400 240289 288406 240301
rect 288458 240289 288464 240341
rect 289168 240289 289174 240341
rect 289226 240329 289232 240341
rect 306928 240329 306934 240341
rect 289226 240301 306934 240329
rect 289226 240289 289232 240301
rect 306928 240289 306934 240301
rect 306986 240289 306992 240341
rect 314608 240289 314614 240341
rect 314666 240329 314672 240341
rect 373264 240329 373270 240341
rect 314666 240301 373270 240329
rect 314666 240289 314672 240301
rect 373264 240289 373270 240301
rect 373322 240289 373328 240341
rect 377872 240289 377878 240341
rect 377930 240329 377936 240341
rect 407536 240329 407542 240341
rect 377930 240301 407542 240329
rect 377930 240289 377936 240301
rect 407536 240289 407542 240301
rect 407594 240289 407600 240341
rect 225424 240215 225430 240267
rect 225482 240255 225488 240267
rect 230896 240255 230902 240267
rect 225482 240227 230902 240255
rect 225482 240215 225488 240227
rect 230896 240215 230902 240227
rect 230954 240215 230960 240267
rect 238768 240215 238774 240267
rect 238826 240255 238832 240267
rect 259408 240255 259414 240267
rect 238826 240227 259414 240255
rect 238826 240215 238832 240227
rect 259408 240215 259414 240227
rect 259466 240215 259472 240267
rect 276784 240215 276790 240267
rect 276842 240255 276848 240267
rect 283888 240255 283894 240267
rect 276842 240227 283894 240255
rect 276842 240215 276848 240227
rect 283888 240215 283894 240227
rect 283946 240215 283952 240267
rect 296560 240255 296566 240267
rect 288034 240227 296566 240255
rect 218416 240141 218422 240193
rect 218474 240181 218480 240193
rect 237904 240181 237910 240193
rect 218474 240153 237910 240181
rect 218474 240141 218480 240153
rect 237904 240141 237910 240153
rect 237962 240141 237968 240193
rect 244144 240141 244150 240193
rect 244202 240181 244208 240193
rect 246352 240181 246358 240193
rect 244202 240153 246358 240181
rect 244202 240141 244208 240153
rect 246352 240141 246358 240153
rect 246410 240141 246416 240193
rect 257200 240141 257206 240193
rect 257258 240181 257264 240193
rect 277840 240181 277846 240193
rect 257258 240153 277846 240181
rect 257258 240141 257264 240153
rect 277840 240141 277846 240153
rect 277898 240141 277904 240193
rect 277936 240141 277942 240193
rect 277994 240181 278000 240193
rect 286768 240181 286774 240193
rect 277994 240153 286774 240181
rect 277994 240141 278000 240153
rect 286768 240141 286774 240153
rect 286826 240141 286832 240193
rect 288034 240181 288062 240227
rect 296560 240215 296566 240227
rect 296618 240215 296624 240267
rect 298096 240215 298102 240267
rect 298154 240255 298160 240267
rect 311632 240255 311638 240267
rect 298154 240227 311638 240255
rect 298154 240215 298160 240227
rect 311632 240215 311638 240227
rect 311690 240215 311696 240267
rect 314224 240215 314230 240267
rect 314282 240255 314288 240267
rect 372400 240255 372406 240267
rect 314282 240227 372406 240255
rect 314282 240215 314288 240227
rect 372400 240215 372406 240227
rect 372458 240215 372464 240267
rect 376432 240215 376438 240267
rect 376490 240255 376496 240267
rect 376490 240227 386942 240255
rect 376490 240215 376496 240227
rect 295792 240181 295798 240193
rect 287938 240153 288062 240181
rect 288130 240153 295798 240181
rect 226288 240067 226294 240119
rect 226346 240107 226352 240119
rect 230704 240107 230710 240119
rect 226346 240079 230710 240107
rect 226346 240067 226352 240079
rect 230704 240067 230710 240079
rect 230762 240067 230768 240119
rect 236464 240067 236470 240119
rect 236522 240107 236528 240119
rect 264400 240107 264406 240119
rect 236522 240079 264406 240107
rect 236522 240067 236528 240079
rect 264400 240067 264406 240079
rect 264458 240067 264464 240119
rect 277648 240067 277654 240119
rect 277706 240107 277712 240119
rect 277706 240079 279422 240107
rect 277706 240067 277712 240079
rect 236272 239993 236278 240045
rect 236330 240033 236336 240045
rect 241648 240033 241654 240045
rect 236330 240005 241654 240033
rect 236330 239993 236336 240005
rect 241648 239993 241654 240005
rect 241706 239993 241712 240045
rect 256432 239993 256438 240045
rect 256490 240033 256496 240045
rect 277744 240033 277750 240045
rect 256490 240005 277750 240033
rect 256490 239993 256496 240005
rect 277744 239993 277750 240005
rect 277802 239993 277808 240045
rect 279394 240033 279422 240079
rect 279472 240067 279478 240119
rect 279530 240107 279536 240119
rect 287938 240107 287966 240153
rect 279530 240079 287966 240107
rect 279530 240067 279536 240079
rect 288130 240033 288158 240153
rect 295792 240141 295798 240153
rect 295850 240141 295856 240193
rect 295888 240141 295894 240193
rect 295946 240181 295952 240193
rect 313168 240181 313174 240193
rect 295946 240153 313174 240181
rect 295946 240141 295952 240153
rect 313168 240141 313174 240153
rect 313226 240141 313232 240193
rect 313456 240141 313462 240193
rect 313514 240181 313520 240193
rect 371344 240181 371350 240193
rect 313514 240153 371350 240181
rect 313514 240141 313520 240153
rect 371344 240141 371350 240153
rect 371402 240141 371408 240193
rect 373072 240141 373078 240193
rect 373130 240181 373136 240193
rect 386800 240181 386806 240193
rect 373130 240153 386806 240181
rect 373130 240141 373136 240153
rect 386800 240141 386806 240153
rect 386858 240141 386864 240193
rect 386914 240181 386942 240227
rect 386992 240215 386998 240267
rect 387050 240255 387056 240267
rect 403216 240255 403222 240267
rect 387050 240227 403222 240255
rect 387050 240215 387056 240227
rect 403216 240215 403222 240227
rect 403274 240215 403280 240267
rect 404080 240181 404086 240193
rect 386914 240153 404086 240181
rect 404080 240141 404086 240153
rect 404138 240141 404144 240193
rect 288208 240067 288214 240119
rect 288266 240107 288272 240119
rect 300592 240107 300598 240119
rect 288266 240079 300598 240107
rect 288266 240067 288272 240079
rect 300592 240067 300598 240079
rect 300650 240067 300656 240119
rect 316816 240067 316822 240119
rect 316874 240107 316880 240119
rect 326992 240107 326998 240119
rect 316874 240079 326998 240107
rect 316874 240067 316880 240079
rect 326992 240067 326998 240079
rect 327050 240067 327056 240119
rect 329296 240067 329302 240119
rect 329354 240107 329360 240119
rect 354544 240107 354550 240119
rect 329354 240079 354550 240107
rect 329354 240067 329360 240079
rect 354544 240067 354550 240079
rect 354602 240067 354608 240119
rect 360592 240067 360598 240119
rect 360650 240107 360656 240119
rect 378736 240107 378742 240119
rect 360650 240079 378742 240107
rect 360650 240067 360656 240079
rect 378736 240067 378742 240079
rect 378794 240067 378800 240119
rect 381808 240067 381814 240119
rect 381866 240107 381872 240119
rect 383056 240107 383062 240119
rect 381866 240079 383062 240107
rect 381866 240067 381872 240079
rect 383056 240067 383062 240079
rect 383114 240067 383120 240119
rect 279394 240005 288158 240033
rect 289072 239993 289078 240045
rect 289130 240033 289136 240045
rect 292624 240033 292630 240045
rect 289130 240005 292630 240033
rect 289130 239993 289136 240005
rect 292624 239993 292630 240005
rect 292682 239993 292688 240045
rect 294256 239993 294262 240045
rect 294314 240033 294320 240045
rect 303568 240033 303574 240045
rect 294314 240005 303574 240033
rect 294314 239993 294320 240005
rect 303568 239993 303574 240005
rect 303626 239993 303632 240045
rect 304720 239993 304726 240045
rect 304778 240033 304784 240045
rect 308176 240033 308182 240045
rect 304778 240005 308182 240033
rect 304778 239993 304784 240005
rect 308176 239993 308182 240005
rect 308234 239993 308240 240045
rect 310480 239993 310486 240045
rect 310538 240033 310544 240045
rect 334384 240033 334390 240045
rect 310538 240005 325406 240033
rect 310538 239993 310544 240005
rect 221488 239919 221494 239971
rect 221546 239959 221552 239971
rect 232912 239959 232918 239971
rect 221546 239931 232918 239959
rect 221546 239919 221552 239931
rect 232912 239919 232918 239931
rect 232970 239919 232976 239971
rect 238288 239919 238294 239971
rect 238346 239959 238352 239971
rect 260656 239959 260662 239971
rect 238346 239931 260662 239959
rect 238346 239919 238352 239931
rect 260656 239919 260662 239931
rect 260714 239919 260720 239971
rect 268720 239919 268726 239971
rect 268778 239959 268784 239971
rect 280336 239959 280342 239971
rect 268778 239931 280342 239959
rect 268778 239919 268784 239931
rect 280336 239919 280342 239931
rect 280394 239919 280400 239971
rect 286960 239919 286966 239971
rect 287018 239959 287024 239971
rect 297616 239959 297622 239971
rect 287018 239931 297622 239959
rect 287018 239919 287024 239931
rect 297616 239919 297622 239931
rect 297674 239919 297680 239971
rect 298192 239919 298198 239971
rect 298250 239959 298256 239971
rect 312784 239959 312790 239971
rect 298250 239931 312790 239959
rect 298250 239919 298256 239931
rect 312784 239919 312790 239931
rect 312842 239919 312848 239971
rect 313744 239919 313750 239971
rect 313802 239959 313808 239971
rect 325264 239959 325270 239971
rect 313802 239931 325270 239959
rect 313802 239919 313808 239931
rect 325264 239919 325270 239931
rect 325322 239919 325328 239971
rect 325378 239959 325406 240005
rect 327202 240005 334390 240033
rect 327202 239959 327230 240005
rect 334384 239993 334390 240005
rect 334442 239993 334448 240045
rect 334480 239993 334486 240045
rect 334538 240033 334544 240045
rect 365872 240033 365878 240045
rect 334538 240005 365878 240033
rect 334538 239993 334544 240005
rect 365872 239993 365878 240005
rect 365930 239993 365936 240045
rect 377200 239993 377206 240045
rect 377258 240033 377264 240045
rect 405520 240033 405526 240045
rect 377258 240005 405526 240033
rect 377258 239993 377264 240005
rect 405520 239993 405526 240005
rect 405578 239993 405584 240045
rect 325378 239931 327230 239959
rect 327856 239919 327862 239971
rect 327914 239959 327920 239971
rect 351760 239959 351766 239971
rect 327914 239931 351766 239959
rect 327914 239919 327920 239931
rect 351760 239919 351766 239931
rect 351818 239919 351824 239971
rect 360208 239919 360214 239971
rect 360266 239959 360272 239971
rect 378640 239959 378646 239971
rect 360266 239931 378646 239959
rect 360266 239919 360272 239931
rect 378640 239919 378646 239931
rect 378698 239919 378704 239971
rect 383056 239959 383062 239971
rect 378754 239931 383062 239959
rect 234544 239845 234550 239897
rect 234602 239885 234608 239897
rect 238576 239885 238582 239897
rect 234602 239857 238582 239885
rect 234602 239845 234608 239857
rect 238576 239845 238582 239857
rect 238634 239845 238640 239897
rect 277072 239845 277078 239897
rect 277130 239885 277136 239897
rect 283792 239885 283798 239897
rect 277130 239857 283798 239885
rect 277130 239845 277136 239857
rect 283792 239845 283798 239857
rect 283850 239845 283856 239897
rect 283888 239845 283894 239897
rect 283946 239885 283952 239897
rect 295216 239885 295222 239897
rect 283946 239857 295222 239885
rect 283946 239845 283952 239857
rect 295216 239845 295222 239857
rect 295274 239845 295280 239897
rect 295696 239845 295702 239897
rect 295754 239885 295760 239897
rect 295754 239857 308030 239885
rect 295754 239845 295760 239857
rect 218704 239771 218710 239823
rect 218762 239811 218768 239823
rect 234352 239811 234358 239823
rect 218762 239783 234358 239811
rect 218762 239771 218768 239783
rect 234352 239771 234358 239783
rect 234410 239771 234416 239823
rect 274864 239771 274870 239823
rect 274922 239811 274928 239823
rect 274922 239783 276446 239811
rect 274922 239771 274928 239783
rect 228016 239697 228022 239749
rect 228074 239737 228080 239749
rect 229936 239737 229942 239749
rect 228074 239709 229942 239737
rect 228074 239697 228080 239709
rect 229936 239697 229942 239709
rect 229994 239697 230000 239749
rect 241072 239697 241078 239749
rect 241130 239737 241136 239749
rect 244624 239737 244630 239749
rect 241130 239709 244630 239737
rect 241130 239697 241136 239709
rect 244624 239697 244630 239709
rect 244682 239697 244688 239749
rect 269392 239697 269398 239749
rect 269450 239737 269456 239749
rect 276304 239737 276310 239749
rect 269450 239709 276310 239737
rect 269450 239697 269456 239709
rect 276304 239697 276310 239709
rect 276362 239697 276368 239749
rect 276418 239737 276446 239783
rect 277648 239771 277654 239823
rect 277706 239811 277712 239823
rect 282928 239811 282934 239823
rect 277706 239783 282934 239811
rect 277706 239771 277712 239783
rect 282928 239771 282934 239783
rect 282986 239771 282992 239823
rect 283024 239771 283030 239823
rect 283082 239811 283088 239823
rect 294736 239811 294742 239823
rect 283082 239783 294742 239811
rect 283082 239771 283088 239783
rect 294736 239771 294742 239783
rect 294794 239771 294800 239823
rect 299056 239771 299062 239823
rect 299114 239811 299120 239823
rect 305776 239811 305782 239823
rect 299114 239783 305782 239811
rect 299114 239771 299120 239783
rect 305776 239771 305782 239783
rect 305834 239771 305840 239823
rect 278032 239737 278038 239749
rect 276418 239709 278038 239737
rect 278032 239697 278038 239709
rect 278090 239697 278096 239749
rect 278224 239697 278230 239749
rect 278282 239737 278288 239749
rect 281776 239737 281782 239749
rect 278282 239709 281782 239737
rect 278282 239697 278288 239709
rect 281776 239697 281782 239709
rect 281834 239697 281840 239749
rect 281872 239697 281878 239749
rect 281930 239737 281936 239749
rect 292144 239737 292150 239749
rect 281930 239709 292150 239737
rect 281930 239697 281936 239709
rect 292144 239697 292150 239709
rect 292202 239697 292208 239749
rect 292240 239697 292246 239749
rect 292298 239737 292304 239749
rect 297904 239737 297910 239749
rect 292298 239709 297910 239737
rect 292298 239697 292304 239709
rect 297904 239697 297910 239709
rect 297962 239697 297968 239749
rect 302992 239697 302998 239749
rect 303050 239737 303056 239749
rect 307600 239737 307606 239749
rect 303050 239709 307606 239737
rect 303050 239697 303056 239709
rect 307600 239697 307606 239709
rect 307658 239697 307664 239749
rect 308002 239737 308030 239857
rect 326608 239845 326614 239897
rect 326666 239885 326672 239897
rect 348688 239885 348694 239897
rect 326666 239857 348694 239885
rect 326666 239845 326672 239857
rect 348688 239845 348694 239857
rect 348746 239845 348752 239897
rect 375664 239845 375670 239897
rect 375722 239885 375728 239897
rect 378754 239885 378782 239931
rect 383056 239919 383062 239931
rect 383114 239919 383120 239971
rect 375722 239857 378782 239885
rect 375722 239845 375728 239857
rect 380848 239845 380854 239897
rect 380906 239885 380912 239897
rect 388144 239885 388150 239897
rect 380906 239857 388150 239885
rect 380906 239845 380912 239857
rect 388144 239845 388150 239857
rect 388202 239845 388208 239897
rect 314800 239811 314806 239823
rect 308290 239783 314806 239811
rect 308290 239737 308318 239783
rect 314800 239771 314806 239783
rect 314858 239771 314864 239823
rect 327088 239771 327094 239823
rect 327146 239811 327152 239823
rect 350032 239811 350038 239823
rect 327146 239783 350038 239811
rect 327146 239771 327152 239783
rect 350032 239771 350038 239783
rect 350090 239771 350096 239823
rect 380560 239771 380566 239823
rect 380618 239811 380624 239823
rect 384880 239811 384886 239823
rect 380618 239783 384886 239811
rect 380618 239771 380624 239783
rect 384880 239771 384886 239783
rect 384938 239771 384944 239823
rect 308002 239709 308318 239737
rect 308848 239697 308854 239749
rect 308906 239737 308912 239749
rect 310192 239737 310198 239749
rect 308906 239709 310198 239737
rect 308906 239697 308912 239709
rect 310192 239697 310198 239709
rect 310250 239697 310256 239749
rect 311632 239697 311638 239749
rect 311690 239737 311696 239749
rect 323632 239737 323638 239749
rect 311690 239709 323638 239737
rect 311690 239697 311696 239709
rect 323632 239697 323638 239709
rect 323690 239697 323696 239749
rect 328816 239737 328822 239749
rect 323746 239709 328822 239737
rect 214480 239623 214486 239675
rect 214538 239663 214544 239675
rect 225136 239663 225142 239675
rect 214538 239635 225142 239663
rect 214538 239623 214544 239635
rect 225136 239623 225142 239635
rect 225194 239623 225200 239675
rect 229072 239623 229078 239675
rect 229130 239663 229136 239675
rect 230224 239663 230230 239675
rect 229130 239635 230230 239663
rect 229130 239623 229136 239635
rect 230224 239623 230230 239635
rect 230282 239623 230288 239675
rect 238192 239623 238198 239675
rect 238250 239663 238256 239675
rect 241840 239663 241846 239675
rect 238250 239635 241846 239663
rect 238250 239623 238256 239635
rect 241840 239623 241846 239635
rect 241898 239623 241904 239675
rect 265648 239623 265654 239675
rect 265706 239663 265712 239675
rect 270160 239663 270166 239675
rect 265706 239635 270166 239663
rect 265706 239623 265712 239635
rect 270160 239623 270166 239635
rect 270218 239623 270224 239675
rect 270256 239623 270262 239675
rect 270314 239663 270320 239675
rect 272272 239663 272278 239675
rect 270314 239635 272278 239663
rect 270314 239623 270320 239635
rect 272272 239623 272278 239635
rect 272330 239623 272336 239675
rect 277936 239663 277942 239675
rect 272386 239635 277942 239663
rect 226288 239549 226294 239601
rect 226346 239589 226352 239601
rect 235792 239589 235798 239601
rect 226346 239561 235798 239589
rect 226346 239549 226352 239561
rect 235792 239549 235798 239561
rect 235850 239549 235856 239601
rect 271408 239549 271414 239601
rect 271466 239589 271472 239601
rect 272386 239589 272414 239635
rect 277936 239623 277942 239635
rect 277994 239623 278000 239675
rect 278896 239623 278902 239675
rect 278954 239663 278960 239675
rect 279664 239663 279670 239675
rect 278954 239635 279670 239663
rect 278954 239623 278960 239635
rect 279664 239623 279670 239635
rect 279722 239623 279728 239675
rect 280528 239623 280534 239675
rect 280586 239663 280592 239675
rect 280586 239635 286622 239663
rect 280586 239623 280592 239635
rect 271466 239561 272414 239589
rect 271466 239549 271472 239561
rect 275344 239549 275350 239601
rect 275402 239589 275408 239601
rect 281104 239589 281110 239601
rect 275402 239561 281110 239589
rect 275402 239549 275408 239561
rect 281104 239549 281110 239561
rect 281162 239549 281168 239601
rect 273520 239475 273526 239527
rect 273578 239515 273584 239527
rect 281584 239515 281590 239527
rect 273578 239487 281590 239515
rect 273578 239475 273584 239487
rect 281584 239475 281590 239487
rect 281642 239475 281648 239527
rect 285040 239475 285046 239527
rect 285098 239515 285104 239527
rect 286594 239515 286622 239635
rect 287056 239623 287062 239675
rect 287114 239663 287120 239675
rect 290800 239663 290806 239675
rect 287114 239635 290806 239663
rect 287114 239623 287120 239635
rect 290800 239623 290806 239635
rect 290858 239623 290864 239675
rect 304048 239623 304054 239675
rect 304106 239663 304112 239675
rect 307984 239663 307990 239675
rect 304106 239635 307990 239663
rect 304106 239623 304112 239635
rect 307984 239623 307990 239635
rect 308042 239623 308048 239675
rect 309520 239623 309526 239675
rect 309578 239663 309584 239675
rect 310288 239663 310294 239675
rect 309578 239635 310294 239663
rect 309578 239623 309584 239635
rect 310288 239623 310294 239635
rect 310346 239623 310352 239675
rect 315664 239623 315670 239675
rect 315722 239663 315728 239675
rect 323746 239663 323774 239709
rect 328816 239697 328822 239709
rect 328874 239697 328880 239749
rect 330064 239697 330070 239749
rect 330122 239737 330128 239749
rect 339184 239737 339190 239749
rect 330122 239709 339190 239737
rect 330122 239697 330128 239709
rect 339184 239697 339190 239709
rect 339242 239697 339248 239749
rect 376048 239697 376054 239749
rect 376106 239737 376112 239749
rect 386992 239737 386998 239749
rect 376106 239709 386998 239737
rect 376106 239697 376112 239709
rect 386992 239697 386998 239709
rect 387050 239697 387056 239749
rect 315722 239635 323774 239663
rect 315722 239623 315728 239635
rect 325648 239623 325654 239675
rect 325706 239663 325712 239675
rect 328624 239663 328630 239675
rect 325706 239635 328630 239663
rect 325706 239623 325712 239635
rect 328624 239623 328630 239635
rect 328682 239623 328688 239675
rect 328720 239623 328726 239675
rect 328778 239663 328784 239675
rect 353488 239663 353494 239675
rect 328778 239635 353494 239663
rect 328778 239623 328784 239635
rect 353488 239623 353494 239635
rect 353546 239623 353552 239675
rect 374800 239623 374806 239675
rect 374858 239663 374864 239675
rect 382672 239663 382678 239675
rect 374858 239635 382678 239663
rect 374858 239623 374864 239635
rect 382672 239623 382678 239635
rect 382730 239623 382736 239675
rect 383248 239623 383254 239675
rect 383306 239663 383312 239675
rect 396400 239663 396406 239675
rect 383306 239635 396406 239663
rect 383306 239623 383312 239635
rect 396400 239623 396406 239635
rect 396458 239623 396464 239675
rect 286672 239549 286678 239601
rect 286730 239589 286736 239601
rect 292528 239589 292534 239601
rect 286730 239561 292534 239589
rect 286730 239549 286736 239561
rect 292528 239549 292534 239561
rect 292586 239549 292592 239601
rect 292624 239549 292630 239601
rect 292682 239589 292688 239601
rect 298000 239589 298006 239601
rect 292682 239561 298006 239589
rect 292682 239549 292688 239561
rect 298000 239549 298006 239561
rect 298058 239549 298064 239601
rect 301840 239549 301846 239601
rect 301898 239589 301904 239601
rect 306832 239589 306838 239601
rect 301898 239561 306838 239589
rect 301898 239549 301904 239561
rect 306832 239549 306838 239561
rect 306890 239549 306896 239601
rect 306928 239549 306934 239601
rect 306986 239589 306992 239601
rect 313840 239589 313846 239601
rect 306986 239561 313846 239589
rect 306986 239549 306992 239561
rect 313840 239549 313846 239561
rect 313898 239549 313904 239601
rect 324400 239549 324406 239601
rect 324458 239589 324464 239601
rect 343696 239589 343702 239601
rect 324458 239561 343702 239589
rect 324458 239549 324464 239561
rect 343696 239549 343702 239561
rect 343754 239549 343760 239601
rect 373840 239549 373846 239601
rect 373898 239589 373904 239601
rect 398608 239589 398614 239601
rect 373898 239561 398614 239589
rect 373898 239549 373904 239561
rect 398608 239549 398614 239561
rect 398666 239549 398672 239601
rect 296944 239515 296950 239527
rect 285098 239487 286526 239515
rect 286594 239487 296950 239515
rect 285098 239475 285104 239487
rect 275920 239401 275926 239453
rect 275978 239441 275984 239453
rect 286000 239441 286006 239453
rect 275978 239413 286006 239441
rect 275978 239401 275984 239413
rect 286000 239401 286006 239413
rect 286058 239401 286064 239453
rect 286498 239441 286526 239487
rect 296944 239475 296950 239487
rect 297002 239475 297008 239527
rect 297616 239475 297622 239527
rect 297674 239515 297680 239527
rect 312592 239515 312598 239527
rect 297674 239487 312598 239515
rect 297674 239475 297680 239487
rect 312592 239475 312598 239487
rect 312650 239475 312656 239527
rect 321616 239475 321622 239527
rect 321674 239515 321680 239527
rect 338896 239515 338902 239527
rect 321674 239487 338902 239515
rect 321674 239475 321680 239487
rect 338896 239475 338902 239487
rect 338954 239475 338960 239527
rect 383056 239515 383062 239527
rect 368770 239487 383062 239515
rect 291856 239441 291862 239453
rect 286498 239413 291862 239441
rect 291856 239401 291862 239413
rect 291914 239401 291920 239453
rect 297520 239441 297526 239453
rect 291970 239413 297526 239441
rect 42544 239367 42550 239379
rect 42370 239339 42550 239367
rect 42370 239305 42398 239339
rect 42544 239327 42550 239339
rect 42602 239327 42608 239379
rect 275440 239327 275446 239379
rect 275498 239367 275504 239379
rect 287728 239367 287734 239379
rect 275498 239339 287734 239367
rect 275498 239327 275504 239339
rect 287728 239327 287734 239339
rect 287786 239327 287792 239379
rect 287824 239327 287830 239379
rect 287882 239367 287888 239379
rect 288976 239367 288982 239379
rect 287882 239339 288982 239367
rect 287882 239327 287888 239339
rect 288976 239327 288982 239339
rect 289034 239327 289040 239379
rect 42352 239253 42358 239305
rect 42410 239253 42416 239305
rect 215920 239253 215926 239305
rect 215978 239293 215984 239305
rect 218896 239293 218902 239305
rect 215978 239265 218902 239293
rect 215978 239253 215984 239265
rect 218896 239253 218902 239265
rect 218954 239253 218960 239305
rect 272464 239253 272470 239305
rect 272522 239293 272528 239305
rect 285520 239293 285526 239305
rect 272522 239265 285526 239293
rect 272522 239253 272528 239265
rect 285520 239253 285526 239265
rect 285578 239253 285584 239305
rect 287248 239253 287254 239305
rect 287306 239293 287312 239305
rect 291970 239293 291998 239413
rect 297520 239401 297526 239413
rect 297578 239401 297584 239453
rect 297808 239401 297814 239453
rect 297866 239441 297872 239453
rect 305008 239441 305014 239453
rect 297866 239413 305014 239441
rect 297866 239401 297872 239413
rect 305008 239401 305014 239413
rect 305066 239401 305072 239453
rect 323056 239401 323062 239453
rect 323114 239441 323120 239453
rect 323114 239413 324830 239441
rect 323114 239401 323120 239413
rect 292048 239327 292054 239379
rect 292106 239367 292112 239379
rect 302416 239367 302422 239379
rect 292106 239339 302422 239367
rect 292106 239327 292112 239339
rect 302416 239327 302422 239339
rect 302474 239327 302480 239379
rect 302512 239327 302518 239379
rect 302570 239367 302576 239379
rect 307216 239367 307222 239379
rect 302570 239339 307222 239367
rect 302570 239327 302576 239339
rect 307216 239327 307222 239339
rect 307274 239327 307280 239379
rect 320848 239327 320854 239379
rect 320906 239367 320912 239379
rect 324688 239367 324694 239379
rect 320906 239339 324694 239367
rect 320906 239327 320912 239339
rect 324688 239327 324694 239339
rect 324746 239327 324752 239379
rect 324802 239367 324830 239413
rect 324880 239401 324886 239453
rect 324938 239441 324944 239453
rect 331312 239441 331318 239453
rect 324938 239413 331318 239441
rect 324938 239401 324944 239413
rect 331312 239401 331318 239413
rect 331370 239401 331376 239453
rect 361552 239401 361558 239453
rect 361610 239441 361616 239453
rect 368770 239441 368798 239487
rect 383056 239475 383062 239487
rect 383114 239475 383120 239527
rect 361610 239413 368798 239441
rect 361610 239401 361616 239413
rect 378640 239401 378646 239453
rect 378698 239441 378704 239453
rect 392080 239441 392086 239453
rect 378698 239413 392086 239441
rect 378698 239401 378704 239413
rect 392080 239401 392086 239413
rect 392138 239401 392144 239453
rect 341296 239367 341302 239379
rect 324802 239339 341302 239367
rect 341296 239327 341302 239339
rect 341354 239327 341360 239379
rect 380080 239327 380086 239379
rect 380138 239367 380144 239379
rect 386608 239367 386614 239379
rect 380138 239339 386614 239367
rect 380138 239327 380144 239339
rect 386608 239327 386614 239339
rect 386666 239327 386672 239379
rect 386704 239327 386710 239379
rect 386762 239367 386768 239379
rect 406672 239367 406678 239379
rect 386762 239339 406678 239367
rect 386762 239327 386768 239339
rect 406672 239327 406678 239339
rect 406730 239327 406736 239379
rect 287306 239265 291998 239293
rect 287306 239253 287312 239265
rect 293200 239253 293206 239305
rect 293258 239293 293264 239305
rect 302800 239293 302806 239305
rect 293258 239265 302806 239293
rect 293258 239253 293264 239265
rect 302800 239253 302806 239265
rect 302858 239253 302864 239305
rect 323440 239253 323446 239305
rect 323498 239293 323504 239305
rect 341968 239293 341974 239305
rect 323498 239265 341974 239293
rect 323498 239253 323504 239265
rect 341968 239253 341974 239265
rect 342026 239253 342032 239305
rect 378736 239253 378742 239305
rect 378794 239293 378800 239305
rect 394096 239293 394102 239305
rect 378794 239265 394102 239293
rect 378794 239253 378800 239265
rect 394096 239253 394102 239265
rect 394154 239253 394160 239305
rect 42544 239179 42550 239231
rect 42602 239219 42608 239231
rect 43216 239219 43222 239231
rect 42602 239191 43222 239219
rect 42602 239179 42608 239191
rect 43216 239179 43222 239191
rect 43274 239179 43280 239231
rect 240496 239179 240502 239231
rect 240554 239219 240560 239231
rect 255664 239219 255670 239231
rect 240554 239191 255670 239219
rect 240554 239179 240560 239191
rect 255664 239179 255670 239191
rect 255722 239179 255728 239231
rect 276208 239179 276214 239231
rect 276266 239219 276272 239231
rect 280432 239219 280438 239231
rect 276266 239191 280438 239219
rect 276266 239179 276272 239191
rect 280432 239179 280438 239191
rect 280490 239179 280496 239231
rect 291472 239179 291478 239231
rect 291530 239219 291536 239231
rect 301840 239219 301846 239231
rect 291530 239191 301846 239219
rect 291530 239179 291536 239191
rect 301840 239179 301846 239191
rect 301898 239179 301904 239231
rect 318256 239179 318262 239231
rect 318314 239219 318320 239231
rect 324880 239219 324886 239231
rect 318314 239191 324886 239219
rect 318314 239179 318320 239191
rect 324880 239179 324886 239191
rect 324938 239179 324944 239231
rect 328624 239179 328630 239231
rect 328682 239219 328688 239231
rect 346960 239219 346966 239231
rect 328682 239191 346966 239219
rect 328682 239179 328688 239191
rect 346960 239179 346966 239191
rect 347018 239179 347024 239231
rect 378640 239179 378646 239231
rect 378698 239219 378704 239231
rect 383824 239219 383830 239231
rect 378698 239191 383830 239219
rect 378698 239179 378704 239191
rect 383824 239179 383830 239191
rect 383882 239179 383888 239231
rect 386800 239179 386806 239231
rect 386858 239219 386864 239231
rect 396880 239219 396886 239231
rect 386858 239191 396886 239219
rect 386858 239179 386864 239191
rect 396880 239179 396886 239191
rect 396938 239179 396944 239231
rect 273232 239105 273238 239157
rect 273290 239145 273296 239157
rect 286672 239145 286678 239157
rect 273290 239117 286678 239145
rect 273290 239105 273296 239117
rect 286672 239105 286678 239117
rect 286730 239105 286736 239157
rect 286768 239105 286774 239157
rect 286826 239145 286832 239157
rect 289360 239145 289366 239157
rect 286826 239117 289366 239145
rect 286826 239105 286832 239117
rect 289360 239105 289366 239117
rect 289418 239105 289424 239157
rect 291856 239105 291862 239157
rect 291914 239145 291920 239157
rect 299152 239145 299158 239157
rect 291914 239117 299158 239145
rect 291914 239105 291920 239117
rect 299152 239105 299158 239117
rect 299210 239105 299216 239157
rect 322672 239105 322678 239157
rect 322730 239145 322736 239157
rect 340912 239145 340918 239157
rect 322730 239117 340918 239145
rect 322730 239105 322736 239117
rect 340912 239105 340918 239117
rect 340970 239105 340976 239157
rect 377488 239105 377494 239157
rect 377546 239145 377552 239157
rect 386704 239145 386710 239157
rect 377546 239117 386710 239145
rect 377546 239105 377552 239117
rect 386704 239105 386710 239117
rect 386762 239105 386768 239157
rect 236176 239031 236182 239083
rect 236234 239071 236240 239083
rect 238384 239071 238390 239083
rect 236234 239043 238390 239071
rect 236234 239031 236240 239043
rect 238384 239031 238390 239043
rect 238442 239031 238448 239083
rect 271888 239031 271894 239083
rect 271946 239071 271952 239083
rect 287824 239071 287830 239083
rect 271946 239043 287830 239071
rect 271946 239031 271952 239043
rect 287824 239031 287830 239043
rect 287882 239031 287888 239083
rect 288976 239031 288982 239083
rect 289034 239071 289040 239083
rect 294448 239071 294454 239083
rect 289034 239043 294454 239071
rect 289034 239031 289040 239043
rect 294448 239031 294454 239043
rect 294506 239031 294512 239083
rect 295984 239031 295990 239083
rect 296042 239071 296048 239083
rect 304048 239071 304054 239083
rect 296042 239043 304054 239071
rect 296042 239031 296048 239043
rect 304048 239031 304054 239043
rect 304106 239031 304112 239083
rect 321232 239031 321238 239083
rect 321290 239071 321296 239083
rect 337168 239071 337174 239083
rect 321290 239043 337174 239071
rect 321290 239031 321296 239043
rect 337168 239031 337174 239043
rect 337226 239031 337232 239083
rect 339856 239031 339862 239083
rect 339914 239071 339920 239083
rect 340240 239071 340246 239083
rect 339914 239043 340246 239071
rect 339914 239031 339920 239043
rect 340240 239031 340246 239043
rect 340298 239031 340304 239083
rect 375184 239031 375190 239083
rect 375242 239071 375248 239083
rect 400624 239071 400630 239083
rect 375242 239043 400630 239071
rect 375242 239031 375248 239043
rect 400624 239031 400630 239043
rect 400682 239031 400688 239083
rect 142960 238957 142966 239009
rect 143018 238997 143024 239009
rect 211024 238997 211030 239009
rect 143018 238969 211030 238997
rect 143018 238957 143024 238969
rect 211024 238957 211030 238969
rect 211082 238997 211088 239009
rect 216688 238997 216694 239009
rect 211082 238969 216694 238997
rect 211082 238957 211088 238969
rect 216688 238957 216694 238969
rect 216746 238957 216752 239009
rect 228112 238957 228118 239009
rect 228170 238997 228176 239009
rect 231952 238997 231958 239009
rect 228170 238969 231958 238997
rect 228170 238957 228176 238969
rect 231952 238957 231958 238969
rect 232010 238957 232016 239009
rect 237520 238957 237526 239009
rect 237578 238997 237584 239009
rect 268144 238997 268150 239009
rect 237578 238969 268150 238997
rect 237578 238957 237584 238969
rect 268144 238957 268150 238969
rect 268202 238957 268208 239009
rect 268240 238957 268246 239009
rect 268298 238997 268304 239009
rect 270928 238997 270934 239009
rect 268298 238969 270934 238997
rect 268298 238957 268304 238969
rect 270928 238957 270934 238969
rect 270986 238957 270992 239009
rect 278512 238957 278518 239009
rect 278570 238997 278576 239009
rect 280720 238997 280726 239009
rect 278570 238969 280726 238997
rect 278570 238957 278576 238969
rect 280720 238957 280726 238969
rect 280778 238957 280784 239009
rect 290896 238957 290902 239009
rect 290954 238997 290960 239009
rect 293296 238997 293302 239009
rect 290954 238969 293302 238997
rect 290954 238957 290960 238969
rect 293296 238957 293302 238969
rect 293354 238957 293360 239009
rect 294064 238957 294070 239009
rect 294122 238997 294128 239009
rect 303184 238997 303190 239009
rect 294122 238969 303190 238997
rect 294122 238957 294128 238969
rect 303184 238957 303190 238969
rect 303242 238957 303248 239009
rect 316432 238957 316438 239009
rect 316490 238997 316496 239009
rect 377296 238997 377302 239009
rect 316490 238969 377302 238997
rect 316490 238957 316496 238969
rect 377296 238957 377302 238969
rect 377354 238957 377360 239009
rect 380464 238957 380470 239009
rect 380522 238997 380528 239009
rect 387568 238997 387574 239009
rect 380522 238969 387574 238997
rect 380522 238957 380528 238969
rect 387568 238957 387574 238969
rect 387626 238957 387632 239009
rect 240112 238883 240118 238935
rect 240170 238923 240176 238935
rect 256816 238923 256822 238935
rect 240170 238895 256822 238923
rect 240170 238883 240176 238895
rect 256816 238883 256822 238895
rect 256874 238883 256880 238935
rect 258256 238883 258262 238935
rect 258314 238923 258320 238935
rect 258314 238895 309182 238923
rect 258314 238883 258320 238895
rect 226864 238809 226870 238861
rect 226922 238849 226928 238861
rect 235024 238849 235030 238861
rect 226922 238821 235030 238849
rect 226922 238809 226928 238821
rect 235024 238809 235030 238821
rect 235082 238809 235088 238861
rect 239152 238809 239158 238861
rect 239210 238849 239216 238861
rect 258544 238849 258550 238861
rect 239210 238821 258550 238849
rect 239210 238809 239216 238821
rect 258544 238809 258550 238821
rect 258602 238809 258608 238861
rect 309154 238849 309182 238895
rect 317680 238883 317686 238935
rect 317738 238923 317744 238935
rect 325936 238923 325942 238935
rect 317738 238895 325942 238923
rect 317738 238883 317744 238895
rect 325936 238883 325942 238895
rect 325994 238883 326000 238935
rect 326704 238883 326710 238935
rect 326762 238923 326768 238935
rect 328912 238923 328918 238935
rect 326762 238895 328918 238923
rect 326762 238883 326768 238895
rect 328912 238883 328918 238895
rect 328970 238883 328976 238935
rect 331888 238883 331894 238935
rect 331946 238923 331952 238935
rect 360496 238923 360502 238935
rect 331946 238895 360502 238923
rect 331946 238883 331952 238895
rect 360496 238883 360502 238895
rect 360554 238883 360560 238935
rect 366832 238883 366838 238935
rect 366890 238923 366896 238935
rect 366890 238895 376094 238923
rect 366890 238883 366896 238895
rect 329104 238849 329110 238861
rect 258658 238821 309086 238849
rect 309154 238821 329110 238849
rect 224560 238735 224566 238787
rect 224618 238775 224624 238787
rect 239536 238775 239542 238787
rect 224618 238747 239542 238775
rect 224618 238735 224624 238747
rect 239536 238735 239542 238747
rect 239594 238735 239600 238787
rect 257776 238735 257782 238787
rect 257834 238775 257840 238787
rect 258658 238775 258686 238821
rect 308944 238775 308950 238787
rect 257834 238747 258686 238775
rect 258754 238747 308950 238775
rect 257834 238735 257840 238747
rect 256048 238661 256054 238713
rect 256106 238701 256112 238713
rect 258754 238701 258782 238747
rect 308944 238735 308950 238747
rect 309002 238735 309008 238787
rect 309058 238775 309086 238821
rect 329104 238809 329110 238821
rect 329162 238809 329168 238861
rect 330640 238809 330646 238861
rect 330698 238849 330704 238861
rect 357232 238849 357238 238861
rect 330698 238821 357238 238849
rect 330698 238809 330704 238821
rect 357232 238809 357238 238821
rect 357290 238809 357296 238861
rect 368176 238809 368182 238861
rect 368234 238849 368240 238861
rect 375952 238849 375958 238861
rect 368234 238821 375958 238849
rect 368234 238809 368240 238821
rect 375952 238809 375958 238821
rect 376010 238809 376016 238861
rect 376066 238849 376094 238895
rect 381424 238883 381430 238935
rect 381482 238923 381488 238935
rect 389200 238923 389206 238935
rect 381482 238895 389206 238923
rect 381482 238883 381488 238895
rect 389200 238883 389206 238895
rect 389258 238883 389264 238935
rect 383344 238849 383350 238861
rect 376066 238821 383350 238849
rect 383344 238809 383350 238821
rect 383402 238809 383408 238861
rect 318160 238775 318166 238787
rect 309058 238747 318166 238775
rect 318160 238735 318166 238747
rect 318218 238735 318224 238787
rect 318640 238735 318646 238787
rect 318698 238775 318704 238787
rect 332176 238775 332182 238787
rect 318698 238747 332182 238775
rect 318698 238735 318704 238747
rect 332176 238735 332182 238747
rect 332234 238735 332240 238787
rect 332272 238735 332278 238787
rect 332330 238775 332336 238787
rect 345904 238775 345910 238787
rect 332330 238747 345910 238775
rect 332330 238735 332336 238747
rect 345904 238735 345910 238747
rect 345962 238735 345968 238787
rect 358768 238775 358774 238787
rect 351298 238747 358774 238775
rect 256106 238673 258782 238701
rect 256106 238661 256112 238673
rect 258832 238661 258838 238713
rect 258890 238701 258896 238713
rect 325840 238701 325846 238713
rect 258890 238673 325846 238701
rect 258890 238661 258896 238673
rect 325840 238661 325846 238673
rect 325898 238661 325904 238713
rect 325936 238661 325942 238713
rect 325994 238701 326000 238713
rect 327568 238701 327574 238713
rect 325994 238673 327574 238701
rect 325994 238661 326000 238673
rect 327568 238661 327574 238673
rect 327626 238661 327632 238713
rect 331120 238661 331126 238713
rect 331178 238701 331184 238713
rect 351298 238701 351326 238747
rect 358768 238735 358774 238747
rect 358826 238735 358832 238787
rect 368560 238735 368566 238787
rect 368618 238775 368624 238787
rect 379024 238775 379030 238787
rect 368618 238747 379030 238775
rect 368618 238735 368624 238747
rect 379024 238735 379030 238747
rect 379082 238735 379088 238787
rect 379696 238735 379702 238787
rect 379754 238775 379760 238787
rect 385360 238775 385366 238787
rect 379754 238747 385366 238775
rect 379754 238735 379760 238747
rect 385360 238735 385366 238747
rect 385418 238735 385424 238787
rect 331178 238673 332222 238701
rect 331178 238661 331184 238673
rect 217072 238587 217078 238639
rect 217130 238627 217136 238639
rect 255184 238627 255190 238639
rect 217130 238599 255190 238627
rect 217130 238587 217136 238599
rect 255184 238587 255190 238599
rect 255242 238587 255248 238639
rect 255568 238587 255574 238639
rect 255626 238627 255632 238639
rect 317968 238627 317974 238639
rect 255626 238599 317974 238627
rect 255626 238587 255632 238599
rect 317968 238587 317974 238599
rect 318026 238587 318032 238639
rect 320080 238587 320086 238639
rect 320138 238627 320144 238639
rect 322096 238627 322102 238639
rect 320138 238599 322102 238627
rect 320138 238587 320144 238599
rect 322096 238587 322102 238599
rect 322154 238587 322160 238639
rect 322288 238587 322294 238639
rect 322346 238627 322352 238639
rect 322346 238599 331742 238627
rect 322346 238587 322352 238599
rect 42160 238513 42166 238565
rect 42218 238553 42224 238565
rect 42352 238553 42358 238565
rect 42218 238525 42358 238553
rect 42218 238513 42224 238525
rect 42352 238513 42358 238525
rect 42410 238513 42416 238565
rect 253840 238513 253846 238565
rect 253898 238553 253904 238565
rect 318064 238553 318070 238565
rect 253898 238525 318070 238553
rect 253898 238513 253904 238525
rect 318064 238513 318070 238525
rect 318122 238513 318128 238565
rect 318160 238513 318166 238565
rect 318218 238553 318224 238565
rect 322384 238553 322390 238565
rect 318218 238525 322390 238553
rect 318218 238513 318224 238525
rect 322384 238513 322390 238525
rect 322442 238513 322448 238565
rect 322480 238513 322486 238565
rect 322538 238553 322544 238565
rect 331600 238553 331606 238565
rect 322538 238525 331606 238553
rect 322538 238513 322544 238525
rect 331600 238513 331606 238525
rect 331658 238513 331664 238565
rect 331714 238553 331742 238599
rect 331792 238587 331798 238639
rect 331850 238627 331856 238639
rect 332080 238627 332086 238639
rect 331850 238599 332086 238627
rect 331850 238587 331856 238599
rect 332080 238587 332086 238599
rect 332138 238587 332144 238639
rect 332194 238627 332222 238673
rect 332386 238673 351326 238701
rect 332386 238627 332414 238673
rect 351376 238661 351382 238713
rect 351434 238701 351440 238713
rect 358864 238701 358870 238713
rect 351434 238673 358870 238701
rect 351434 238661 351440 238673
rect 358864 238661 358870 238673
rect 358922 238661 358928 238713
rect 372592 238661 372598 238713
rect 372650 238701 372656 238713
rect 383056 238701 383062 238713
rect 372650 238673 383062 238701
rect 372650 238661 372656 238673
rect 383056 238661 383062 238673
rect 383114 238661 383120 238713
rect 332194 238599 332414 238627
rect 334096 238587 334102 238639
rect 334154 238627 334160 238639
rect 365296 238627 365302 238639
rect 334154 238599 365302 238627
rect 334154 238587 334160 238599
rect 365296 238587 365302 238599
rect 365354 238587 365360 238639
rect 368656 238587 368662 238639
rect 368714 238627 368720 238639
rect 387088 238627 387094 238639
rect 368714 238599 387094 238627
rect 368714 238587 368720 238599
rect 387088 238587 387094 238599
rect 387146 238587 387152 238639
rect 334960 238553 334966 238565
rect 331714 238525 334966 238553
rect 334960 238513 334966 238525
rect 335018 238513 335024 238565
rect 335074 238525 335294 238553
rect 218032 238439 218038 238491
rect 218090 238479 218096 238491
rect 253456 238479 253462 238491
rect 218090 238451 253462 238479
rect 218090 238439 218096 238451
rect 253456 238439 253462 238451
rect 253514 238439 253520 238491
rect 254608 238439 254614 238491
rect 254666 238479 254672 238491
rect 335074 238479 335102 238525
rect 254666 238451 335102 238479
rect 335266 238479 335294 238525
rect 335344 238513 335350 238565
rect 335402 238553 335408 238565
rect 348016 238553 348022 238565
rect 335402 238525 348022 238553
rect 335402 238513 335408 238525
rect 348016 238513 348022 238525
rect 348074 238513 348080 238565
rect 375952 238513 375958 238565
rect 376010 238553 376016 238565
rect 384592 238553 384598 238565
rect 376010 238525 384598 238553
rect 376010 238513 376016 238525
rect 384592 238513 384598 238525
rect 384650 238513 384656 238565
rect 336976 238479 336982 238491
rect 335266 238451 336982 238479
rect 254666 238439 254672 238451
rect 336976 238439 336982 238451
rect 337034 238439 337040 238491
rect 369424 238439 369430 238491
rect 369482 238479 369488 238491
rect 388816 238479 388822 238491
rect 369482 238451 388822 238479
rect 369482 238439 369488 238451
rect 388816 238439 388822 238451
rect 388874 238439 388880 238491
rect 216304 238365 216310 238417
rect 216362 238405 216368 238417
rect 237520 238405 237526 238417
rect 216362 238377 237526 238405
rect 216362 238365 216368 238377
rect 237520 238365 237526 238377
rect 237578 238365 237584 238417
rect 240592 238365 240598 238417
rect 240650 238405 240656 238417
rect 317680 238405 317686 238417
rect 240650 238377 317686 238405
rect 240650 238365 240656 238377
rect 317680 238365 317686 238377
rect 317738 238365 317744 238417
rect 318064 238365 318070 238417
rect 318122 238405 318128 238417
rect 318122 238377 322430 238405
rect 318122 238365 318128 238377
rect 253360 238291 253366 238343
rect 253418 238331 253424 238343
rect 322402 238331 322430 238377
rect 322480 238365 322486 238417
rect 322538 238405 322544 238417
rect 330736 238405 330742 238417
rect 322538 238377 330742 238405
rect 322538 238365 322544 238377
rect 330736 238365 330742 238377
rect 330794 238365 330800 238417
rect 335248 238365 335254 238417
rect 335306 238405 335312 238417
rect 367024 238405 367030 238417
rect 335306 238377 367030 238405
rect 335306 238365 335312 238377
rect 367024 238365 367030 238377
rect 367082 238365 367088 238417
rect 371632 238365 371638 238417
rect 371690 238405 371696 238417
rect 393616 238405 393622 238417
rect 371690 238377 393622 238405
rect 371690 238365 371696 238377
rect 393616 238365 393622 238377
rect 393674 238365 393680 238417
rect 338704 238331 338710 238343
rect 253418 238303 322142 238331
rect 322402 238303 338710 238331
rect 253418 238291 253424 238303
rect 252400 238217 252406 238269
rect 252458 238257 252464 238269
rect 321904 238257 321910 238269
rect 252458 238229 321910 238257
rect 252458 238217 252464 238229
rect 321904 238217 321910 238229
rect 321962 238217 321968 238269
rect 322114 238257 322142 238303
rect 338704 238291 338710 238303
rect 338762 238291 338768 238343
rect 370384 238291 370390 238343
rect 370442 238331 370448 238343
rect 390352 238331 390358 238343
rect 370442 238303 390358 238331
rect 370442 238291 370448 238303
rect 390352 238291 390358 238303
rect 390410 238291 390416 238343
rect 639760 238291 639766 238343
rect 639818 238331 639824 238343
rect 649936 238331 649942 238343
rect 639818 238303 649942 238331
rect 639818 238291 639824 238303
rect 649936 238291 649942 238303
rect 649994 238291 650000 238343
rect 322114 238229 331550 238257
rect 251632 238143 251638 238195
rect 251690 238183 251696 238195
rect 331522 238183 331550 238229
rect 331600 238217 331606 238269
rect 331658 238257 331664 238269
rect 341488 238257 341494 238269
rect 331658 238229 341494 238257
rect 331658 238217 331664 238229
rect 341488 238217 341494 238229
rect 341546 238217 341552 238269
rect 369808 238217 369814 238269
rect 369866 238257 369872 238269
rect 389680 238257 389686 238269
rect 369866 238229 389686 238257
rect 369866 238217 369872 238229
rect 389680 238217 389686 238229
rect 389738 238217 389744 238269
rect 340432 238183 340438 238195
rect 251690 238155 331454 238183
rect 331522 238155 340438 238183
rect 251690 238143 251696 238155
rect 228208 238069 228214 238121
rect 228266 238109 228272 238121
rect 245872 238109 245878 238121
rect 228266 238081 245878 238109
rect 228266 238069 228272 238081
rect 245872 238069 245878 238081
rect 245930 238069 245936 238121
rect 251152 238069 251158 238121
rect 251210 238109 251216 238121
rect 331426 238109 331454 238155
rect 340432 238143 340438 238155
rect 340490 238143 340496 238195
rect 370864 238143 370870 238195
rect 370922 238183 370928 238195
rect 391888 238183 391894 238195
rect 370922 238155 391894 238183
rect 370922 238143 370928 238155
rect 391888 238143 391894 238155
rect 391946 238143 391952 238195
rect 343504 238109 343510 238121
rect 251210 238081 331358 238109
rect 331426 238081 343510 238109
rect 251210 238069 251216 238081
rect 222832 237995 222838 238047
rect 222890 238035 222896 238047
rect 243760 238035 243766 238047
rect 222890 238007 243766 238035
rect 222890 237995 222896 238007
rect 243760 237995 243766 238007
rect 243818 237995 243824 238047
rect 249424 237995 249430 238047
rect 249482 238035 249488 238047
rect 321904 238035 321910 238047
rect 249482 238007 321910 238035
rect 249482 237995 249488 238007
rect 321904 237995 321910 238007
rect 321962 237995 321968 238047
rect 322096 237995 322102 238047
rect 322154 238035 322160 238047
rect 322154 238007 322430 238035
rect 322154 237995 322160 238007
rect 223312 237921 223318 237973
rect 223370 237961 223376 237973
rect 242416 237961 242422 237973
rect 223370 237933 242422 237961
rect 223370 237921 223376 237933
rect 242416 237921 242422 237933
rect 242474 237921 242480 237973
rect 250192 237921 250198 237973
rect 250250 237961 250256 237973
rect 315856 237961 315862 237973
rect 250250 237933 315862 237961
rect 250250 237921 250256 237933
rect 315856 237921 315862 237933
rect 315914 237921 315920 237973
rect 322288 237961 322294 237973
rect 315970 237933 322294 237961
rect 42160 237847 42166 237899
rect 42218 237887 42224 237899
rect 47536 237887 47542 237899
rect 42218 237859 47542 237887
rect 42218 237847 42224 237859
rect 47536 237847 47542 237859
rect 47594 237847 47600 237899
rect 222928 237847 222934 237899
rect 222986 237887 222992 237899
rect 222986 237859 228446 237887
rect 222986 237847 222992 237859
rect 221872 237773 221878 237825
rect 221930 237813 221936 237825
rect 228418 237813 228446 237859
rect 228496 237847 228502 237899
rect 228554 237887 228560 237899
rect 230800 237887 230806 237899
rect 228554 237859 230806 237887
rect 228554 237847 228560 237859
rect 230800 237847 230806 237859
rect 230858 237847 230864 237899
rect 247984 237847 247990 237899
rect 248042 237887 248048 237899
rect 315970 237887 315998 237933
rect 322288 237921 322294 237933
rect 322346 237921 322352 237973
rect 322402 237961 322430 238007
rect 322480 237995 322486 238047
rect 322538 238035 322544 238047
rect 326800 238035 326806 238047
rect 322538 238007 326806 238035
rect 322538 237995 322544 238007
rect 326800 237995 326806 238007
rect 326858 237995 326864 238047
rect 331330 238035 331358 238081
rect 343504 238069 343510 238081
rect 343562 238069 343568 238121
rect 372016 238069 372022 238121
rect 372074 238109 372080 238121
rect 394192 238109 394198 238121
rect 372074 238081 394198 238109
rect 372074 238069 372080 238081
rect 394192 238069 394198 238081
rect 394250 238069 394256 238121
rect 345232 238035 345238 238047
rect 331330 238007 345238 238035
rect 345232 237995 345238 238007
rect 345290 237995 345296 238047
rect 371248 237995 371254 238047
rect 371306 238035 371312 238047
rect 392464 238035 392470 238047
rect 371306 238007 392470 238035
rect 371306 237995 371312 238007
rect 392464 237995 392470 238007
rect 392522 237995 392528 238047
rect 346288 237961 346294 237973
rect 322402 237933 346294 237961
rect 346288 237921 346294 237933
rect 346346 237921 346352 237973
rect 375280 237921 375286 237973
rect 375338 237961 375344 237973
rect 401200 237961 401206 237973
rect 375338 237933 401206 237961
rect 375338 237921 375344 237933
rect 401200 237921 401206 237933
rect 401258 237921 401264 237973
rect 639376 237921 639382 237973
rect 639434 237961 639440 237973
rect 649744 237961 649750 237973
rect 639434 237933 649750 237961
rect 639434 237921 639440 237933
rect 649744 237921 649750 237933
rect 649802 237921 649808 237973
rect 248042 237859 315998 237887
rect 248042 237847 248048 237859
rect 316048 237847 316054 237899
rect 316106 237887 316112 237899
rect 316106 237859 322526 237887
rect 316106 237847 316112 237859
rect 242608 237813 242614 237825
rect 221930 237785 228350 237813
rect 228418 237785 242614 237813
rect 221930 237773 221936 237785
rect 221488 237699 221494 237751
rect 221546 237739 221552 237751
rect 228208 237739 228214 237751
rect 221546 237711 228214 237739
rect 221546 237699 221552 237711
rect 228208 237699 228214 237711
rect 228266 237699 228272 237751
rect 228322 237739 228350 237785
rect 242608 237773 242614 237785
rect 242666 237773 242672 237825
rect 247216 237773 247222 237825
rect 247274 237813 247280 237825
rect 315760 237813 315766 237825
rect 247274 237785 315766 237813
rect 247274 237773 247280 237785
rect 315760 237773 315766 237785
rect 315818 237773 315824 237825
rect 315856 237773 315862 237825
rect 315914 237813 315920 237825
rect 322000 237813 322006 237825
rect 315914 237785 322006 237813
rect 315914 237773 315920 237785
rect 322000 237773 322006 237785
rect 322058 237773 322064 237825
rect 322498 237813 322526 237859
rect 326800 237847 326806 237899
rect 326858 237887 326864 237899
rect 351280 237887 351286 237899
rect 326858 237859 351286 237887
rect 326858 237847 326864 237859
rect 351280 237847 351286 237859
rect 351338 237847 351344 237899
rect 362800 237847 362806 237899
rect 362858 237887 362864 237899
rect 382288 237887 382294 237899
rect 362858 237859 382294 237887
rect 362858 237847 362864 237859
rect 382288 237847 382294 237859
rect 382346 237847 382352 237899
rect 384112 237847 384118 237899
rect 384170 237887 384176 237899
rect 410416 237887 410422 237899
rect 384170 237859 410422 237887
rect 384170 237847 384176 237859
rect 410416 237847 410422 237859
rect 410474 237847 410480 237899
rect 637936 237847 637942 237899
rect 637994 237887 638000 237899
rect 650416 237887 650422 237899
rect 637994 237859 650422 237887
rect 637994 237847 638000 237859
rect 650416 237847 650422 237859
rect 650474 237847 650480 237899
rect 353008 237813 353014 237825
rect 322498 237785 353014 237813
rect 353008 237773 353014 237785
rect 353066 237773 353072 237825
rect 359824 237773 359830 237825
rect 359882 237813 359888 237825
rect 380944 237813 380950 237825
rect 359882 237785 380950 237813
rect 359882 237773 359888 237785
rect 380944 237773 380950 237785
rect 381002 237773 381008 237825
rect 384496 237773 384502 237825
rect 384554 237813 384560 237825
rect 410992 237813 410998 237825
rect 384554 237785 410998 237813
rect 384554 237773 384560 237785
rect 410992 237773 410998 237785
rect 411050 237773 411056 237825
rect 638896 237773 638902 237825
rect 638954 237813 638960 237825
rect 649552 237813 649558 237825
rect 638954 237785 649558 237813
rect 638954 237773 638960 237785
rect 649552 237773 649558 237785
rect 649610 237773 649616 237825
rect 244816 237739 244822 237751
rect 228322 237711 244822 237739
rect 244816 237699 244822 237711
rect 244874 237699 244880 237751
rect 245776 237699 245782 237751
rect 245834 237739 245840 237751
rect 356176 237739 356182 237751
rect 245834 237711 356182 237739
rect 245834 237699 245840 237711
rect 356176 237699 356182 237711
rect 356234 237699 356240 237751
rect 637360 237699 637366 237751
rect 637418 237739 637424 237751
rect 650128 237739 650134 237751
rect 637418 237711 650134 237739
rect 637418 237699 637424 237711
rect 650128 237699 650134 237711
rect 650186 237699 650192 237751
rect 224080 237625 224086 237677
rect 224138 237665 224144 237677
rect 240688 237665 240694 237677
rect 224138 237637 240694 237665
rect 224138 237625 224144 237637
rect 240688 237625 240694 237637
rect 240746 237625 240752 237677
rect 246736 237625 246742 237677
rect 246794 237665 246800 237677
rect 315568 237665 315574 237677
rect 246794 237637 315574 237665
rect 246794 237625 246800 237637
rect 315568 237625 315574 237637
rect 315626 237625 315632 237677
rect 322384 237625 322390 237677
rect 322442 237665 322448 237677
rect 354448 237665 354454 237677
rect 322442 237637 354454 237665
rect 322442 237625 322448 237637
rect 354448 237625 354454 237637
rect 354506 237625 354512 237677
rect 549232 237625 549238 237677
rect 549290 237665 549296 237677
rect 650992 237665 650998 237677
rect 549290 237637 650998 237665
rect 549290 237625 549296 237637
rect 650992 237625 650998 237637
rect 651050 237625 651056 237677
rect 148336 237551 148342 237603
rect 148394 237591 148400 237603
rect 207088 237591 207094 237603
rect 148394 237563 207094 237591
rect 148394 237551 148400 237563
rect 207088 237551 207094 237563
rect 207146 237591 207152 237603
rect 221968 237591 221974 237603
rect 207146 237563 221974 237591
rect 207146 237551 207152 237563
rect 221968 237551 221974 237563
rect 222026 237551 222032 237603
rect 223696 237551 223702 237603
rect 223754 237591 223760 237603
rect 241552 237591 241558 237603
rect 223754 237563 241558 237591
rect 223754 237551 223760 237563
rect 241552 237551 241558 237563
rect 241610 237551 241616 237603
rect 245008 237551 245014 237603
rect 245066 237591 245072 237603
rect 357808 237591 357814 237603
rect 245066 237563 357814 237591
rect 245066 237551 245072 237563
rect 357808 237551 357814 237563
rect 357866 237551 357872 237603
rect 374224 237551 374230 237603
rect 374282 237591 374288 237603
rect 399664 237591 399670 237603
rect 374282 237563 399670 237591
rect 374282 237551 374288 237563
rect 399664 237551 399670 237563
rect 399722 237551 399728 237603
rect 420592 237551 420598 237603
rect 420650 237591 420656 237603
rect 608176 237591 608182 237603
rect 420650 237563 608182 237591
rect 420650 237551 420656 237563
rect 608176 237551 608182 237563
rect 608234 237551 608240 237603
rect 637840 237551 637846 237603
rect 637898 237591 637904 237603
rect 650224 237591 650230 237603
rect 637898 237563 650230 237591
rect 637898 237551 637904 237563
rect 650224 237551 650230 237563
rect 650282 237551 650288 237603
rect 256816 237477 256822 237529
rect 256874 237517 256880 237529
rect 310000 237517 310006 237529
rect 256874 237489 310006 237517
rect 256874 237477 256880 237489
rect 310000 237477 310006 237489
rect 310058 237477 310064 237529
rect 317584 237517 317590 237529
rect 315490 237489 317590 237517
rect 248944 237403 248950 237455
rect 249002 237443 249008 237455
rect 258832 237443 258838 237455
rect 249002 237415 258838 237443
rect 249002 237403 249008 237415
rect 258832 237403 258838 237415
rect 258890 237403 258896 237455
rect 268144 237403 268150 237455
rect 268202 237443 268208 237455
rect 282256 237443 282262 237455
rect 268202 237415 282262 237443
rect 268202 237403 268208 237415
rect 282256 237403 282262 237415
rect 282314 237403 282320 237455
rect 286480 237403 286486 237455
rect 286538 237443 286544 237455
rect 287152 237443 287158 237455
rect 286538 237415 287158 237443
rect 286538 237403 286544 237415
rect 287152 237403 287158 237415
rect 287210 237403 287216 237455
rect 292528 237403 292534 237455
rect 292586 237443 292592 237455
rect 293680 237443 293686 237455
rect 292586 237415 293686 237443
rect 292586 237403 292592 237415
rect 293680 237403 293686 237415
rect 293738 237403 293744 237455
rect 293776 237403 293782 237455
rect 293834 237443 293840 237455
rect 295408 237443 295414 237455
rect 293834 237415 295414 237443
rect 293834 237403 293840 237415
rect 295408 237403 295414 237415
rect 295466 237403 295472 237455
rect 304720 237403 304726 237455
rect 304778 237443 304784 237455
rect 315376 237443 315382 237455
rect 304778 237415 315382 237443
rect 304778 237403 304784 237415
rect 315376 237403 315382 237415
rect 315434 237403 315440 237455
rect 239536 237329 239542 237381
rect 239594 237369 239600 237381
rect 257392 237369 257398 237381
rect 239594 237341 257398 237369
rect 239594 237329 239600 237341
rect 257392 237329 257398 237341
rect 257450 237329 257456 237381
rect 274192 237329 274198 237381
rect 274250 237369 274256 237381
rect 281488 237369 281494 237381
rect 274250 237341 281494 237369
rect 274250 237329 274256 237341
rect 281488 237329 281494 237341
rect 281546 237329 281552 237381
rect 281680 237329 281686 237381
rect 281738 237369 281744 237381
rect 286768 237369 286774 237381
rect 281738 237341 286774 237369
rect 281738 237329 281744 237341
rect 286768 237329 286774 237341
rect 286826 237329 286832 237381
rect 291280 237329 291286 237381
rect 291338 237369 291344 237381
rect 315490 237369 315518 237489
rect 317584 237477 317590 237489
rect 317642 237477 317648 237529
rect 319024 237477 319030 237529
rect 319082 237517 319088 237529
rect 332368 237517 332374 237529
rect 319082 237489 332374 237517
rect 319082 237477 319088 237489
rect 332368 237477 332374 237489
rect 332426 237477 332432 237529
rect 332752 237477 332758 237529
rect 332810 237517 332816 237529
rect 347920 237517 347926 237529
rect 332810 237489 347926 237517
rect 332810 237477 332816 237489
rect 347920 237477 347926 237489
rect 347978 237477 347984 237529
rect 373456 237477 373462 237529
rect 373514 237517 373520 237529
rect 397936 237517 397942 237529
rect 373514 237489 397942 237517
rect 373514 237477 373520 237489
rect 397936 237477 397942 237489
rect 397994 237477 398000 237529
rect 315568 237403 315574 237455
rect 315626 237443 315632 237455
rect 322384 237443 322390 237455
rect 315626 237415 322390 237443
rect 315626 237403 315632 237415
rect 322384 237403 322390 237415
rect 322442 237403 322448 237455
rect 322480 237403 322486 237455
rect 322538 237443 322544 237455
rect 322538 237415 368702 237443
rect 322538 237403 322544 237415
rect 291338 237341 315518 237369
rect 291338 237329 291344 237341
rect 317392 237329 317398 237381
rect 317450 237369 317456 237381
rect 368560 237369 368566 237381
rect 317450 237341 368566 237369
rect 317450 237329 317456 237341
rect 368560 237329 368566 237341
rect 368618 237329 368624 237381
rect 368674 237369 368702 237415
rect 372976 237403 372982 237455
rect 373034 237443 373040 237455
rect 396208 237443 396214 237455
rect 373034 237415 396214 237443
rect 373034 237403 373040 237415
rect 396208 237403 396214 237415
rect 396266 237403 396272 237455
rect 376624 237369 376630 237381
rect 368674 237341 376630 237369
rect 376624 237329 376630 237341
rect 376682 237329 376688 237381
rect 225520 237255 225526 237307
rect 225578 237295 225584 237307
rect 237424 237295 237430 237307
rect 225578 237267 237430 237295
rect 225578 237255 225584 237267
rect 237424 237255 237430 237267
rect 237482 237255 237488 237307
rect 276688 237255 276694 237307
rect 276746 237295 276752 237307
rect 284464 237295 284470 237307
rect 276746 237267 284470 237295
rect 276746 237255 276752 237267
rect 284464 237255 284470 237267
rect 284522 237255 284528 237307
rect 287152 237255 287158 237307
rect 287210 237295 287216 237307
rect 299632 237295 299638 237307
rect 287210 237267 299638 237295
rect 287210 237255 287216 237267
rect 299632 237255 299638 237267
rect 299690 237255 299696 237307
rect 299728 237255 299734 237307
rect 299786 237295 299792 237307
rect 322288 237295 322294 237307
rect 299786 237267 322294 237295
rect 299786 237255 299792 237267
rect 322288 237255 322294 237267
rect 322346 237255 322352 237307
rect 322768 237255 322774 237307
rect 322826 237295 322832 237307
rect 358384 237295 358390 237307
rect 322826 237267 358390 237295
rect 322826 237255 322832 237267
rect 358384 237255 358390 237267
rect 358442 237255 358448 237307
rect 369040 237255 369046 237307
rect 369098 237295 369104 237307
rect 369098 237267 380126 237295
rect 369098 237255 369104 237267
rect 227344 237181 227350 237233
rect 227402 237221 227408 237233
rect 233488 237221 233494 237233
rect 227402 237193 233494 237221
rect 227402 237181 227408 237193
rect 233488 237181 233494 237193
rect 233546 237181 233552 237233
rect 275824 237181 275830 237233
rect 275882 237221 275888 237233
rect 286576 237221 286582 237233
rect 275882 237193 286582 237221
rect 275882 237181 275888 237193
rect 286576 237181 286582 237193
rect 286634 237181 286640 237233
rect 291664 237221 291670 237233
rect 286978 237193 291670 237221
rect 273520 237107 273526 237159
rect 273578 237147 273584 237159
rect 286978 237147 287006 237193
rect 291664 237181 291670 237193
rect 291722 237181 291728 237233
rect 291778 237193 310430 237221
rect 273578 237119 287006 237147
rect 273578 237107 273584 237119
rect 291376 237107 291382 237159
rect 291434 237147 291440 237159
rect 291778 237147 291806 237193
rect 291434 237119 291806 237147
rect 291434 237107 291440 237119
rect 302320 237107 302326 237159
rect 302378 237147 302384 237159
rect 305872 237147 305878 237159
rect 302378 237119 305878 237147
rect 302378 237107 302384 237119
rect 305872 237107 305878 237119
rect 305930 237107 305936 237159
rect 310402 237147 310430 237193
rect 315568 237181 315574 237233
rect 315626 237221 315632 237233
rect 316624 237221 316630 237233
rect 315626 237193 316630 237221
rect 315626 237181 315632 237193
rect 316624 237181 316630 237193
rect 316682 237181 316688 237233
rect 339856 237221 339862 237233
rect 322498 237193 339862 237221
rect 322498 237159 322526 237193
rect 339856 237181 339862 237193
rect 339914 237181 339920 237233
rect 380098 237221 380126 237267
rect 380176 237255 380182 237307
rect 380234 237295 380240 237307
rect 385936 237295 385942 237307
rect 380234 237267 385942 237295
rect 380234 237255 380240 237267
rect 385936 237255 385942 237267
rect 385994 237255 386000 237307
rect 387664 237221 387670 237233
rect 380098 237193 387670 237221
rect 387664 237181 387670 237193
rect 387722 237181 387728 237233
rect 318448 237147 318454 237159
rect 310402 237119 318454 237147
rect 318448 237107 318454 237119
rect 318506 237107 318512 237159
rect 322480 237107 322486 237159
rect 322538 237107 322544 237159
rect 329680 237107 329686 237159
rect 329738 237147 329744 237159
rect 355696 237147 355702 237159
rect 329738 237119 355702 237147
rect 329738 237107 329744 237119
rect 355696 237107 355702 237119
rect 355754 237107 355760 237159
rect 379984 237107 379990 237159
rect 380042 237147 380048 237159
rect 380176 237147 380182 237159
rect 380042 237119 380182 237147
rect 380042 237107 380048 237119
rect 380176 237107 380182 237119
rect 380234 237107 380240 237159
rect 221104 237033 221110 237085
rect 221162 237073 221168 237085
rect 246544 237073 246550 237085
rect 221162 237045 246550 237073
rect 221162 237033 221168 237045
rect 246544 237033 246550 237045
rect 246602 237033 246608 237085
rect 282736 237033 282742 237085
rect 282794 237073 282800 237085
rect 282794 237045 289214 237073
rect 282794 237033 282800 237045
rect 227248 236959 227254 237011
rect 227306 236999 227312 237011
rect 234064 236999 234070 237011
rect 227306 236971 234070 236999
rect 227306 236959 227312 236971
rect 234064 236959 234070 236971
rect 234122 236959 234128 237011
rect 277264 236959 277270 237011
rect 277322 236999 277328 237011
rect 279760 236999 279766 237011
rect 277322 236971 279766 236999
rect 277322 236959 277328 236971
rect 279760 236959 279766 236971
rect 279818 236959 279824 237011
rect 288976 236999 288982 237011
rect 279874 236971 288982 236999
rect 220720 236885 220726 236937
rect 220778 236925 220784 236937
rect 246928 236925 246934 236937
rect 220778 236897 246934 236925
rect 220778 236885 220784 236897
rect 246928 236885 246934 236897
rect 246986 236885 246992 236937
rect 271024 236885 271030 236937
rect 271082 236925 271088 236937
rect 279874 236925 279902 236971
rect 288976 236959 288982 236971
rect 289034 236959 289040 237011
rect 289186 236999 289214 237045
rect 289264 237033 289270 237085
rect 289322 237073 289328 237085
rect 300976 237073 300982 237085
rect 289322 237045 300982 237073
rect 289322 237033 289328 237045
rect 300976 237033 300982 237045
rect 301034 237033 301040 237085
rect 310000 237033 310006 237085
rect 310058 237073 310064 237085
rect 324112 237073 324118 237085
rect 310058 237045 324118 237073
rect 310058 237033 310064 237045
rect 324112 237033 324118 237045
rect 324170 237033 324176 237085
rect 327472 237033 327478 237085
rect 327530 237073 327536 237085
rect 350704 237073 350710 237085
rect 327530 237045 350710 237073
rect 327530 237033 327536 237045
rect 350704 237033 350710 237045
rect 350762 237033 350768 237085
rect 298000 236999 298006 237011
rect 289186 236971 298006 236999
rect 298000 236959 298006 236971
rect 298058 236959 298064 237011
rect 300784 236959 300790 237011
rect 300842 236999 300848 237011
rect 306256 236999 306262 237011
rect 300842 236971 306262 236999
rect 300842 236959 300848 236971
rect 306256 236959 306262 236971
rect 306314 236959 306320 237011
rect 326704 236959 326710 237011
rect 326762 236999 326768 237011
rect 349552 236999 349558 237011
rect 326762 236971 349558 236999
rect 326762 236959 326768 236971
rect 349552 236959 349558 236971
rect 349610 236959 349616 237011
rect 271082 236897 279902 236925
rect 271082 236885 271088 236897
rect 284368 236885 284374 236937
rect 284426 236925 284432 236937
rect 298768 236925 298774 236937
rect 284426 236897 298774 236925
rect 284426 236885 284432 236897
rect 298768 236885 298774 236897
rect 298826 236885 298832 236937
rect 326224 236885 326230 236937
rect 326282 236925 326288 236937
rect 332752 236925 332758 236937
rect 326282 236897 332758 236925
rect 326282 236885 326288 236897
rect 332752 236885 332758 236897
rect 332810 236885 332816 236937
rect 332848 236885 332854 236937
rect 332906 236925 332912 236937
rect 339472 236925 339478 236937
rect 332906 236897 339478 236925
rect 332906 236885 332912 236897
rect 339472 236885 339478 236897
rect 339530 236885 339536 236937
rect 217456 236811 217462 236863
rect 217514 236851 217520 236863
rect 254320 236851 254326 236863
rect 217514 236823 254326 236851
rect 217514 236811 217520 236823
rect 254320 236811 254326 236823
rect 254378 236811 254384 236863
rect 278800 236811 278806 236863
rect 278858 236851 278864 236863
rect 278858 236823 295262 236851
rect 278858 236811 278864 236823
rect 274672 236737 274678 236789
rect 274730 236777 274736 236789
rect 294352 236777 294358 236789
rect 274730 236749 294358 236777
rect 274730 236737 274736 236749
rect 294352 236737 294358 236749
rect 294410 236737 294416 236789
rect 295234 236777 295262 236823
rect 295312 236811 295318 236863
rect 295370 236851 295376 236863
rect 303664 236851 303670 236863
rect 295370 236823 303670 236851
rect 295370 236811 295376 236823
rect 303664 236811 303670 236823
rect 303722 236811 303728 236863
rect 308944 236811 308950 236863
rect 309002 236851 309008 236863
rect 333904 236851 333910 236863
rect 309002 236823 333910 236851
rect 309002 236811 309008 236823
rect 333904 236811 333910 236823
rect 333962 236811 333968 236863
rect 370768 236811 370774 236863
rect 370826 236851 370832 236863
rect 381136 236851 381142 236863
rect 370826 236823 381142 236851
rect 370826 236811 370832 236823
rect 381136 236811 381142 236823
rect 381194 236811 381200 236863
rect 296176 236777 296182 236789
rect 295234 236749 296182 236777
rect 296176 236737 296182 236749
rect 296234 236737 296240 236789
rect 328240 236737 328246 236789
rect 328298 236777 328304 236789
rect 352432 236777 352438 236789
rect 328298 236749 352438 236777
rect 328298 236737 328304 236749
rect 352432 236737 352438 236749
rect 352490 236737 352496 236789
rect 42160 236663 42166 236715
rect 42218 236703 42224 236715
rect 42928 236703 42934 236715
rect 42218 236675 42934 236703
rect 42218 236663 42224 236675
rect 42928 236663 42934 236675
rect 42986 236663 42992 236715
rect 278416 236663 278422 236715
rect 278474 236703 278480 236715
rect 279376 236703 279382 236715
rect 278474 236675 279382 236703
rect 278474 236663 278480 236675
rect 279376 236663 279382 236675
rect 279434 236663 279440 236715
rect 285808 236663 285814 236715
rect 285866 236703 285872 236715
rect 299248 236703 299254 236715
rect 285866 236675 299254 236703
rect 285866 236663 285872 236675
rect 299248 236663 299254 236675
rect 299306 236663 299312 236715
rect 324496 236663 324502 236715
rect 324554 236703 324560 236715
rect 344752 236703 344758 236715
rect 324554 236675 344758 236703
rect 324554 236663 324560 236675
rect 344752 236663 344758 236675
rect 344810 236663 344816 236715
rect 381904 236663 381910 236715
rect 381962 236703 381968 236715
rect 390928 236703 390934 236715
rect 381962 236675 390934 236703
rect 381962 236663 381968 236675
rect 390928 236663 390934 236675
rect 390986 236663 390992 236715
rect 258160 236589 258166 236641
rect 258218 236629 258224 236641
rect 262288 236629 262294 236641
rect 258218 236601 262294 236629
rect 258218 236589 258224 236601
rect 262288 236589 262294 236601
rect 262346 236589 262352 236641
rect 268336 236589 268342 236641
rect 268394 236629 268400 236641
rect 281392 236629 281398 236641
rect 268394 236601 281398 236629
rect 268394 236589 268400 236601
rect 281392 236589 281398 236601
rect 281450 236589 281456 236641
rect 288688 236589 288694 236641
rect 288746 236629 288752 236641
rect 312112 236629 312118 236641
rect 288746 236601 312118 236629
rect 288746 236589 288752 236601
rect 312112 236589 312118 236601
rect 312170 236589 312176 236641
rect 325264 236589 325270 236641
rect 325322 236629 325328 236641
rect 331696 236629 331702 236641
rect 325322 236601 331702 236629
rect 325322 236589 325328 236601
rect 331696 236589 331702 236601
rect 331754 236589 331760 236641
rect 343024 236629 343030 236641
rect 331810 236601 343030 236629
rect 274096 236515 274102 236567
rect 274154 236555 274160 236567
rect 289648 236555 289654 236567
rect 274154 236527 289654 236555
rect 274154 236515 274160 236527
rect 289648 236515 289654 236527
rect 289706 236515 289712 236567
rect 289936 236515 289942 236567
rect 289994 236555 290000 236567
rect 304720 236555 304726 236567
rect 289994 236527 304726 236555
rect 289994 236515 290000 236527
rect 304720 236515 304726 236527
rect 304778 236515 304784 236567
rect 324016 236515 324022 236567
rect 324074 236555 324080 236567
rect 331810 236555 331838 236601
rect 343024 236589 343030 236601
rect 343082 236589 343088 236641
rect 338224 236555 338230 236567
rect 324074 236527 331838 236555
rect 331906 236527 338230 236555
rect 324074 236515 324080 236527
rect 225040 236441 225046 236493
rect 225098 236481 225104 236493
rect 238864 236481 238870 236493
rect 225098 236453 238870 236481
rect 225098 236441 225104 236453
rect 238864 236441 238870 236453
rect 238922 236441 238928 236493
rect 276400 236441 276406 236493
rect 276458 236481 276464 236493
rect 294832 236481 294838 236493
rect 276458 236453 294838 236481
rect 276458 236441 276464 236453
rect 294832 236441 294838 236453
rect 294890 236441 294896 236493
rect 321808 236441 321814 236493
rect 321866 236481 321872 236493
rect 331906 236481 331934 236527
rect 338224 236515 338230 236527
rect 338282 236515 338288 236567
rect 321866 236453 331934 236481
rect 321866 236441 321872 236453
rect 205936 236367 205942 236419
rect 205994 236367 206000 236419
rect 272656 236367 272662 236419
rect 272714 236407 272720 236419
rect 272714 236379 288926 236407
rect 272714 236367 272720 236379
rect 146800 236219 146806 236271
rect 146858 236259 146864 236271
rect 168400 236259 168406 236271
rect 146858 236231 168406 236259
rect 146858 236219 146864 236231
rect 168400 236219 168406 236231
rect 168458 236219 168464 236271
rect 205954 236197 205982 236367
rect 271504 236293 271510 236345
rect 271562 236333 271568 236345
rect 271562 236305 281342 236333
rect 271562 236293 271568 236305
rect 227728 236219 227734 236271
rect 227786 236259 227792 236271
rect 232816 236259 232822 236271
rect 227786 236231 232822 236259
rect 227786 236219 227792 236231
rect 232816 236219 232822 236231
rect 232874 236219 232880 236271
rect 236560 236219 236566 236271
rect 236618 236259 236624 236271
rect 238960 236259 238966 236271
rect 236618 236231 238966 236259
rect 236618 236219 236624 236231
rect 238960 236219 238966 236231
rect 239018 236219 239024 236271
rect 278128 236219 278134 236271
rect 278186 236259 278192 236271
rect 281200 236259 281206 236271
rect 278186 236231 281206 236259
rect 278186 236219 278192 236231
rect 281200 236219 281206 236231
rect 281258 236219 281264 236271
rect 281314 236259 281342 236305
rect 281392 236293 281398 236345
rect 281450 236333 281456 236345
rect 288112 236333 288118 236345
rect 281450 236305 288118 236333
rect 281450 236293 281456 236305
rect 288112 236293 288118 236305
rect 288170 236293 288176 236345
rect 288898 236333 288926 236379
rect 288976 236367 288982 236419
rect 289034 236407 289040 236419
rect 297328 236407 297334 236419
rect 289034 236379 297334 236407
rect 289034 236367 289040 236379
rect 297328 236367 297334 236379
rect 297386 236367 297392 236419
rect 288898 236305 289694 236333
rect 289360 236259 289366 236271
rect 281314 236231 289366 236259
rect 289360 236219 289366 236231
rect 289418 236219 289424 236271
rect 145552 236145 145558 236197
rect 145610 236185 145616 236197
rect 146416 236185 146422 236197
rect 145610 236157 146422 236185
rect 145610 236145 145616 236157
rect 146416 236145 146422 236157
rect 146474 236145 146480 236197
rect 146704 236145 146710 236197
rect 146762 236185 146768 236197
rect 174160 236185 174166 236197
rect 146762 236157 174166 236185
rect 146762 236145 146768 236157
rect 174160 236145 174166 236157
rect 174218 236145 174224 236197
rect 205936 236145 205942 236197
rect 205994 236145 206000 236197
rect 210256 236145 210262 236197
rect 210314 236185 210320 236197
rect 210640 236185 210646 236197
rect 210314 236157 210646 236185
rect 210314 236145 210320 236157
rect 210640 236145 210646 236157
rect 210698 236185 210704 236197
rect 213040 236185 213046 236197
rect 210698 236157 213046 236185
rect 210698 236145 210704 236157
rect 213040 236145 213046 236157
rect 213098 236145 213104 236197
rect 225904 236145 225910 236197
rect 225962 236185 225968 236197
rect 236752 236185 236758 236197
rect 225962 236157 236758 236185
rect 225962 236145 225968 236157
rect 236752 236145 236758 236157
rect 236810 236145 236816 236197
rect 289666 236185 289694 236305
rect 290320 236293 290326 236345
rect 290378 236333 290384 236345
rect 301456 236333 301462 236345
rect 290378 236305 301462 236333
rect 290378 236293 290384 236305
rect 301456 236293 301462 236305
rect 301514 236293 301520 236345
rect 332272 236293 332278 236345
rect 332330 236333 332336 236345
rect 361072 236333 361078 236345
rect 332330 236305 361078 236333
rect 332330 236293 332336 236305
rect 361072 236293 361078 236305
rect 361130 236293 361136 236345
rect 290800 236219 290806 236271
rect 290858 236259 290864 236271
rect 293968 236259 293974 236271
rect 290858 236231 293974 236259
rect 290858 236219 290864 236231
rect 293968 236219 293974 236231
rect 294026 236219 294032 236271
rect 297520 236219 297526 236271
rect 297578 236259 297584 236271
rect 300208 236259 300214 236271
rect 297578 236231 300214 236259
rect 297578 236219 297584 236231
rect 300208 236219 300214 236231
rect 300266 236219 300272 236271
rect 319984 236219 319990 236271
rect 320042 236259 320048 236271
rect 334192 236259 334198 236271
rect 320042 236231 334198 236259
rect 320042 236219 320048 236231
rect 334192 236219 334198 236231
rect 334250 236219 334256 236271
rect 335056 236219 335062 236271
rect 335114 236259 335120 236271
rect 335248 236259 335254 236271
rect 335114 236231 335254 236259
rect 335114 236219 335120 236231
rect 335248 236219 335254 236231
rect 335306 236219 335312 236271
rect 290896 236185 290902 236197
rect 289666 236157 290902 236185
rect 290896 236145 290902 236157
rect 290954 236145 290960 236197
rect 291760 236145 291766 236197
rect 291818 236185 291824 236197
rect 319312 236185 319318 236197
rect 291818 236157 319318 236185
rect 291818 236145 291824 236157
rect 319312 236145 319318 236157
rect 319370 236145 319376 236197
rect 320464 236145 320470 236197
rect 320522 236185 320528 236197
rect 336112 236185 336118 236197
rect 320522 236157 336118 236185
rect 320522 236145 320528 236157
rect 336112 236145 336118 236157
rect 336170 236145 336176 236197
rect 541456 236145 541462 236197
rect 541514 236185 541520 236197
rect 549232 236185 549238 236197
rect 541514 236157 549238 236185
rect 541514 236145 541520 236157
rect 549232 236145 549238 236157
rect 549290 236145 549296 236197
rect 638704 236145 638710 236197
rect 638762 236185 638768 236197
rect 639184 236185 639190 236197
rect 638762 236157 639190 236185
rect 638762 236145 638768 236157
rect 639184 236145 639190 236157
rect 639242 236145 639248 236197
rect 265936 236071 265942 236123
rect 265994 236111 266000 236123
rect 339952 236111 339958 236123
rect 265994 236083 339958 236111
rect 265994 236071 266000 236083
rect 339952 236071 339958 236083
rect 340010 236071 340016 236123
rect 264784 235997 264790 236049
rect 264842 236037 264848 236049
rect 310768 236037 310774 236049
rect 264842 236009 310774 236037
rect 264842 235997 264848 236009
rect 310768 235997 310774 236009
rect 310826 235997 310832 236049
rect 312976 235997 312982 236049
rect 313034 236037 313040 236049
rect 369616 236037 369622 236049
rect 313034 236009 369622 236037
rect 313034 235997 313040 236009
rect 369616 235997 369622 236009
rect 369674 235997 369680 236049
rect 267664 235923 267670 235975
rect 267722 235963 267728 235975
rect 340720 235963 340726 235975
rect 267722 235935 340726 235963
rect 267722 235923 267728 235935
rect 340720 235923 340726 235935
rect 340778 235923 340784 235975
rect 262864 235849 262870 235901
rect 262922 235889 262928 235901
rect 338512 235889 338518 235901
rect 262922 235861 338518 235889
rect 262922 235849 262928 235861
rect 338512 235849 338518 235861
rect 338570 235849 338576 235901
rect 258352 235775 258358 235827
rect 258410 235815 258416 235827
rect 336304 235815 336310 235827
rect 258410 235787 336310 235815
rect 258410 235775 258416 235787
rect 336304 235775 336310 235787
rect 336362 235775 336368 235827
rect 261136 235701 261142 235753
rect 261194 235741 261200 235753
rect 337744 235741 337750 235753
rect 261194 235713 337750 235741
rect 261194 235701 261200 235713
rect 337744 235701 337750 235713
rect 337802 235701 337808 235753
rect 256336 235627 256342 235679
rect 256394 235667 256400 235679
rect 335536 235667 335542 235679
rect 256394 235639 335542 235667
rect 256394 235627 256400 235639
rect 335536 235627 335542 235639
rect 335594 235627 335600 235679
rect 260080 235553 260086 235605
rect 260138 235593 260144 235605
rect 336976 235593 336982 235605
rect 260138 235565 336982 235593
rect 260138 235553 260144 235565
rect 336976 235553 336982 235565
rect 337034 235553 337040 235605
rect 273904 235479 273910 235531
rect 273962 235519 273968 235531
rect 355408 235519 355414 235531
rect 273962 235491 355414 235519
rect 273962 235479 273968 235491
rect 355408 235479 355414 235491
rect 355466 235479 355472 235531
rect 42160 235405 42166 235457
rect 42218 235445 42224 235457
rect 43024 235445 43030 235457
rect 42218 235417 43030 235445
rect 42218 235405 42224 235417
rect 43024 235405 43030 235417
rect 43082 235405 43088 235457
rect 236080 235405 236086 235457
rect 236138 235445 236144 235457
rect 265456 235445 265462 235457
rect 236138 235417 265462 235445
rect 236138 235405 236144 235417
rect 265456 235405 265462 235417
rect 265514 235405 265520 235457
rect 273808 235405 273814 235457
rect 273866 235445 273872 235457
rect 356176 235445 356182 235457
rect 273866 235417 356182 235445
rect 273866 235405 273872 235417
rect 356176 235405 356182 235417
rect 356234 235405 356240 235457
rect 245680 235331 245686 235383
rect 245738 235371 245744 235383
rect 353968 235371 353974 235383
rect 245738 235343 353974 235371
rect 245738 235331 245744 235343
rect 353968 235331 353974 235343
rect 354026 235331 354032 235383
rect 239344 235257 239350 235309
rect 239402 235297 239408 235309
rect 350992 235297 350998 235309
rect 239402 235269 350998 235297
rect 239402 235257 239408 235269
rect 350992 235257 350998 235269
rect 351050 235257 351056 235309
rect 146128 235183 146134 235235
rect 146186 235223 146192 235235
rect 146416 235223 146422 235235
rect 146186 235195 146422 235223
rect 146186 235183 146192 235195
rect 146416 235183 146422 235195
rect 146474 235183 146480 235235
rect 246352 235183 246358 235235
rect 246410 235223 246416 235235
rect 353200 235223 353206 235235
rect 246410 235195 353206 235223
rect 246410 235183 246416 235195
rect 353200 235183 353206 235195
rect 353258 235183 353264 235235
rect 241840 235109 241846 235161
rect 241898 235149 241904 235161
rect 350032 235149 350038 235161
rect 241898 235121 350038 235149
rect 241898 235109 241904 235121
rect 350032 235109 350038 235121
rect 350090 235109 350096 235161
rect 238672 235035 238678 235087
rect 238730 235075 238736 235087
rect 347824 235075 347830 235087
rect 238730 235047 347830 235075
rect 238730 235035 238736 235047
rect 347824 235035 347830 235047
rect 347882 235035 347888 235087
rect 241648 234961 241654 235013
rect 241706 235001 241712 235013
rect 349552 235001 349558 235013
rect 241706 234973 349558 235001
rect 241706 234961 241712 234973
rect 349552 234961 349558 234973
rect 349610 234961 349616 235013
rect 244624 234887 244630 234939
rect 244682 234927 244688 234939
rect 351760 234927 351766 234939
rect 244682 234899 351766 234927
rect 244682 234887 244688 234899
rect 351760 234887 351766 234899
rect 351818 234887 351824 234939
rect 42160 234813 42166 234865
rect 42218 234853 42224 234865
rect 42352 234853 42358 234865
rect 42218 234825 42358 234853
rect 42218 234813 42224 234825
rect 42352 234813 42358 234825
rect 42410 234813 42416 234865
rect 238576 234813 238582 234865
rect 238634 234853 238640 234865
rect 348784 234853 348790 234865
rect 238634 234825 348790 234853
rect 238634 234813 238640 234825
rect 348784 234813 348790 234825
rect 348842 234813 348848 234865
rect 231664 234739 231670 234791
rect 231722 234779 231728 234791
rect 347344 234779 347350 234791
rect 231722 234751 347350 234779
rect 231722 234739 231728 234751
rect 347344 234739 347350 234751
rect 347402 234739 347408 234791
rect 226960 234665 226966 234717
rect 227018 234705 227024 234717
rect 345136 234705 345142 234717
rect 227018 234677 345142 234705
rect 227018 234665 227024 234677
rect 345136 234665 345142 234677
rect 345194 234665 345200 234717
rect 265264 234591 265270 234643
rect 265322 234631 265328 234643
rect 308848 234631 308854 234643
rect 265322 234603 308854 234631
rect 265322 234591 265328 234603
rect 308848 234591 308854 234603
rect 308906 234591 308912 234643
rect 312016 234591 312022 234643
rect 312074 234631 312080 234643
rect 367696 234631 367702 234643
rect 312074 234603 367702 234631
rect 312074 234591 312080 234603
rect 367696 234591 367702 234603
rect 367754 234591 367760 234643
rect 266608 234517 266614 234569
rect 266666 234557 266672 234569
rect 306736 234557 306742 234569
rect 266666 234529 306742 234557
rect 266666 234517 266672 234529
rect 306736 234517 306742 234529
rect 306794 234517 306800 234569
rect 316048 234517 316054 234569
rect 316106 234557 316112 234569
rect 322384 234557 322390 234569
rect 316106 234529 322390 234557
rect 316106 234517 316112 234529
rect 322384 234517 322390 234529
rect 322442 234517 322448 234569
rect 266032 234443 266038 234495
rect 266090 234483 266096 234495
rect 307312 234483 307318 234495
rect 266090 234455 307318 234483
rect 266090 234443 266096 234455
rect 307312 234443 307318 234455
rect 307370 234443 307376 234495
rect 368560 234443 368566 234495
rect 368618 234483 368624 234495
rect 379984 234483 379990 234495
rect 368618 234455 379990 234483
rect 368618 234443 368624 234455
rect 379984 234443 379990 234455
rect 380042 234443 380048 234495
rect 283312 234369 283318 234421
rect 283370 234409 283376 234421
rect 320368 234409 320374 234421
rect 283370 234381 320374 234409
rect 283370 234369 283376 234381
rect 320368 234369 320374 234381
rect 320426 234369 320432 234421
rect 283696 234295 283702 234347
rect 283754 234335 283760 234347
rect 319696 234335 319702 234347
rect 283754 234307 319702 234335
rect 283754 234295 283760 234307
rect 319696 234295 319702 234307
rect 319754 234295 319760 234347
rect 383056 234295 383062 234347
rect 383114 234335 383120 234347
rect 384400 234335 384406 234347
rect 383114 234307 384406 234335
rect 383114 234295 383120 234307
rect 384400 234295 384406 234307
rect 384458 234295 384464 234347
rect 267088 234221 267094 234273
rect 267146 234261 267152 234273
rect 305104 234261 305110 234273
rect 267146 234233 305110 234261
rect 267146 234221 267152 234233
rect 305104 234221 305110 234233
rect 305162 234221 305168 234273
rect 42064 234147 42070 234199
rect 42122 234187 42128 234199
rect 43120 234187 43126 234199
rect 42122 234159 43126 234187
rect 42122 234147 42128 234159
rect 43120 234147 43126 234159
rect 43178 234147 43184 234199
rect 267856 234147 267862 234199
rect 267914 234187 267920 234199
rect 303376 234187 303382 234199
rect 267914 234159 303382 234187
rect 267914 234147 267920 234159
rect 303376 234147 303382 234159
rect 303434 234147 303440 234199
rect 268816 234073 268822 234125
rect 268874 234113 268880 234125
rect 301936 234113 301942 234125
rect 268874 234085 301942 234113
rect 268874 234073 268880 234085
rect 301936 234073 301942 234085
rect 301994 234073 302000 234125
rect 269296 233999 269302 234051
rect 269354 234039 269360 234051
rect 300304 234039 300310 234051
rect 269354 234011 300310 234039
rect 269354 233999 269360 234011
rect 300304 233999 300310 234011
rect 300362 233999 300368 234051
rect 293488 233925 293494 233977
rect 293546 233965 293552 233977
rect 322576 233965 322582 233977
rect 293546 233937 322582 233965
rect 293546 233925 293552 233937
rect 322576 233925 322582 233937
rect 322634 233925 322640 233977
rect 269872 233851 269878 233903
rect 269930 233891 269936 233903
rect 301360 233891 301366 233903
rect 269930 233863 301366 233891
rect 269930 233851 269936 233863
rect 301360 233851 301366 233863
rect 301418 233851 301424 233903
rect 286480 233777 286486 233829
rect 286538 233817 286544 233829
rect 314320 233817 314326 233829
rect 286538 233789 314326 233817
rect 286538 233777 286544 233789
rect 314320 233777 314326 233789
rect 314378 233777 314384 233829
rect 292864 233703 292870 233755
rect 292922 233743 292928 233755
rect 321424 233743 321430 233755
rect 292922 233715 321430 233743
rect 292922 233703 292928 233715
rect 321424 233703 321430 233715
rect 321482 233703 321488 233755
rect 210352 233629 210358 233681
rect 210410 233669 210416 233681
rect 212368 233669 212374 233681
rect 210410 233641 212374 233669
rect 210410 233629 210416 233641
rect 212368 233629 212374 233641
rect 212426 233629 212432 233681
rect 286096 233629 286102 233681
rect 286154 233669 286160 233681
rect 315088 233669 315094 233681
rect 286154 233641 315094 233669
rect 286154 233629 286160 233641
rect 315088 233629 315094 233641
rect 315146 233629 315152 233681
rect 208048 233555 208054 233607
rect 208106 233595 208112 233607
rect 213520 233595 213526 233607
rect 208106 233567 213526 233595
rect 208106 233555 208112 233567
rect 213520 233555 213526 233567
rect 213578 233555 213584 233607
rect 269104 233555 269110 233607
rect 269162 233555 269168 233607
rect 270256 233555 270262 233607
rect 270314 233595 270320 233607
rect 298576 233595 298582 233607
rect 270314 233567 298582 233595
rect 270314 233555 270320 233567
rect 298576 233555 298582 233567
rect 298634 233555 298640 233607
rect 210064 233481 210070 233533
rect 210122 233521 210128 233533
rect 213136 233521 213142 233533
rect 210122 233493 213142 233521
rect 210122 233481 210128 233493
rect 213136 233481 213142 233493
rect 213194 233481 213200 233533
rect 213904 233481 213910 233533
rect 213962 233481 213968 233533
rect 209968 233407 209974 233459
rect 210026 233447 210032 233459
rect 213922 233447 213950 233481
rect 210026 233419 213950 233447
rect 269122 233447 269150 233555
rect 289840 233481 289846 233533
rect 289898 233521 289904 233533
rect 295696 233521 295702 233533
rect 289898 233493 295702 233521
rect 289898 233481 289904 233493
rect 295696 233481 295702 233493
rect 295754 233481 295760 233533
rect 297040 233481 297046 233533
rect 297098 233481 297104 233533
rect 297058 233447 297086 233481
rect 269122 233419 297086 233447
rect 210026 233407 210032 233419
rect 146800 233259 146806 233311
rect 146858 233299 146864 233311
rect 171280 233299 171286 233311
rect 146858 233271 171286 233299
rect 146858 233259 146864 233271
rect 171280 233259 171286 233271
rect 171338 233259 171344 233311
rect 645712 232889 645718 232941
rect 645770 232929 645776 232941
rect 649840 232929 649846 232941
rect 645770 232901 649846 232929
rect 645770 232889 645776 232901
rect 649840 232889 649846 232901
rect 649898 232889 649904 232941
rect 42256 232519 42262 232571
rect 42314 232559 42320 232571
rect 43216 232559 43222 232571
rect 42314 232531 43222 232559
rect 42314 232519 42320 232531
rect 43216 232519 43222 232531
rect 43274 232519 43280 232571
rect 645136 232297 645142 232349
rect 645194 232337 645200 232349
rect 645520 232337 645526 232349
rect 645194 232309 645526 232337
rect 645194 232297 645200 232309
rect 645520 232297 645526 232309
rect 645578 232337 645584 232349
rect 649648 232337 649654 232349
rect 645578 232309 649654 232337
rect 645578 232297 645584 232309
rect 649648 232297 649654 232309
rect 649706 232297 649712 232349
rect 204976 232075 204982 232127
rect 205034 232115 205040 232127
rect 205552 232115 205558 232127
rect 205034 232087 205558 232115
rect 205034 232075 205040 232087
rect 205552 232075 205558 232087
rect 205610 232075 205616 232127
rect 645136 231557 645142 231609
rect 645194 231597 645200 231609
rect 650512 231597 650518 231609
rect 645194 231569 650518 231597
rect 645194 231557 645200 231569
rect 650512 231557 650518 231569
rect 650570 231557 650576 231609
rect 645136 231113 645142 231165
rect 645194 231153 645200 231165
rect 645328 231153 645334 231165
rect 645194 231125 645334 231153
rect 645194 231113 645200 231125
rect 645328 231113 645334 231125
rect 645386 231153 645392 231165
rect 650320 231153 650326 231165
rect 645386 231125 650326 231153
rect 645386 231113 645392 231125
rect 650320 231113 650326 231125
rect 650378 231113 650384 231165
rect 645136 230669 645142 230721
rect 645194 230709 645200 230721
rect 650032 230709 650038 230721
rect 645194 230681 650038 230709
rect 645194 230669 645200 230681
rect 650032 230669 650038 230681
rect 650090 230669 650096 230721
rect 146800 230521 146806 230573
rect 146858 230561 146864 230573
rect 151120 230561 151126 230573
rect 146858 230533 151126 230561
rect 146858 230521 146864 230533
rect 151120 230521 151126 230533
rect 151178 230521 151184 230573
rect 144400 230447 144406 230499
rect 144458 230487 144464 230499
rect 165520 230487 165526 230499
rect 144458 230459 165526 230487
rect 144458 230447 144464 230459
rect 165520 230447 165526 230459
rect 165578 230447 165584 230499
rect 666640 229485 666646 229537
rect 666698 229525 666704 229537
rect 674416 229525 674422 229537
rect 666698 229497 674422 229525
rect 666698 229485 666704 229497
rect 674416 229485 674422 229497
rect 674474 229485 674480 229537
rect 669616 228893 669622 228945
rect 669674 228933 669680 228945
rect 674704 228933 674710 228945
rect 669674 228905 674710 228933
rect 669674 228893 669680 228905
rect 674704 228893 674710 228905
rect 674762 228893 674768 228945
rect 146800 228745 146806 228797
rect 146858 228785 146864 228797
rect 159760 228785 159766 228797
rect 146858 228757 159766 228785
rect 146858 228745 146864 228757
rect 159760 228745 159766 228757
rect 159818 228745 159824 228797
rect 669712 227857 669718 227909
rect 669770 227897 669776 227909
rect 674416 227897 674422 227909
rect 669770 227869 674422 227897
rect 669770 227857 669776 227869
rect 674416 227857 674422 227869
rect 674474 227857 674480 227909
rect 146704 227635 146710 227687
rect 146762 227675 146768 227687
rect 162640 227675 162646 227687
rect 146762 227647 162646 227675
rect 146762 227635 146768 227647
rect 162640 227635 162646 227647
rect 162698 227635 162704 227687
rect 43216 227561 43222 227613
rect 43274 227601 43280 227613
rect 43504 227601 43510 227613
rect 43274 227573 43510 227601
rect 43274 227561 43280 227573
rect 43504 227561 43510 227573
rect 43562 227561 43568 227613
rect 146800 227561 146806 227613
rect 146858 227601 146864 227613
rect 202960 227601 202966 227613
rect 146858 227573 202966 227601
rect 146858 227561 146864 227573
rect 202960 227561 202966 227573
rect 203018 227561 203024 227613
rect 146320 227487 146326 227539
rect 146378 227527 146384 227539
rect 146512 227527 146518 227539
rect 146378 227499 146518 227527
rect 146378 227487 146384 227499
rect 146512 227487 146518 227499
rect 146570 227487 146576 227539
rect 205072 227413 205078 227465
rect 205130 227453 205136 227465
rect 207376 227453 207382 227465
rect 205130 227425 207382 227453
rect 205130 227413 205136 227425
rect 207376 227413 207382 227425
rect 207434 227413 207440 227465
rect 144016 226377 144022 226429
rect 144074 226417 144080 226429
rect 156880 226417 156886 226429
rect 144074 226389 156886 226417
rect 144074 226377 144080 226389
rect 156880 226377 156886 226389
rect 156938 226377 156944 226429
rect 673360 225785 673366 225837
rect 673418 225825 673424 225837
rect 674704 225825 674710 225837
rect 673418 225797 674710 225825
rect 673418 225785 673424 225797
rect 674704 225785 674710 225797
rect 674762 225825 674768 225837
rect 679792 225825 679798 225837
rect 674762 225797 679798 225825
rect 674762 225785 674768 225797
rect 679792 225785 679798 225797
rect 679850 225785 679856 225837
rect 206128 224823 206134 224875
rect 206186 224823 206192 224875
rect 144016 224675 144022 224727
rect 144074 224715 144080 224727
rect 200080 224715 200086 224727
rect 144074 224687 200086 224715
rect 144074 224675 144080 224687
rect 200080 224675 200086 224687
rect 200138 224675 200144 224727
rect 206146 224653 206174 224823
rect 673840 224675 673846 224727
rect 673898 224715 673904 224727
rect 679984 224715 679990 224727
rect 673898 224687 679990 224715
rect 673898 224675 673904 224687
rect 679984 224675 679990 224687
rect 680042 224675 680048 224727
rect 141040 224601 141046 224653
rect 141098 224641 141104 224653
rect 204496 224641 204502 224653
rect 141098 224613 204502 224641
rect 141098 224601 141104 224613
rect 204496 224601 204502 224613
rect 204554 224601 204560 224653
rect 206128 224601 206134 224653
rect 206186 224601 206192 224653
rect 146608 224527 146614 224579
rect 146666 224567 146672 224579
rect 205456 224567 205462 224579
rect 146666 224539 205462 224567
rect 146666 224527 146672 224539
rect 205456 224527 205462 224539
rect 205514 224527 205520 224579
rect 206416 224527 206422 224579
rect 206474 224567 206480 224579
rect 206800 224567 206806 224579
rect 206474 224539 206806 224567
rect 206474 224527 206480 224539
rect 206800 224527 206806 224539
rect 206858 224527 206864 224579
rect 149680 224453 149686 224505
rect 149738 224493 149744 224505
rect 204592 224493 204598 224505
rect 149738 224465 204598 224493
rect 149738 224453 149744 224465
rect 204592 224453 204598 224465
rect 204650 224453 204656 224505
rect 152560 224379 152566 224431
rect 152618 224419 152624 224431
rect 206416 224419 206422 224431
rect 152618 224391 206422 224419
rect 152618 224379 152624 224391
rect 206416 224379 206422 224391
rect 206474 224379 206480 224431
rect 144016 221863 144022 221915
rect 144074 221903 144080 221915
rect 179920 221903 179926 221915
rect 144074 221875 179926 221903
rect 144074 221863 144080 221875
rect 179920 221863 179926 221875
rect 179978 221863 179984 221915
rect 144112 221789 144118 221841
rect 144170 221829 144176 221841
rect 182800 221829 182806 221841
rect 144170 221801 182806 221829
rect 144170 221789 144176 221801
rect 182800 221789 182806 221801
rect 182858 221789 182864 221841
rect 146128 221715 146134 221767
rect 146186 221755 146192 221767
rect 146224 221755 146230 221767
rect 146186 221727 146230 221755
rect 146186 221715 146192 221727
rect 146224 221715 146230 221727
rect 146282 221715 146288 221767
rect 155440 221715 155446 221767
rect 155498 221755 155504 221767
rect 204496 221755 204502 221767
rect 155498 221727 204502 221755
rect 155498 221715 155504 221727
rect 204496 221715 204502 221727
rect 204554 221715 204560 221767
rect 161200 221641 161206 221693
rect 161258 221681 161264 221693
rect 204976 221681 204982 221693
rect 161258 221653 204982 221681
rect 161258 221641 161264 221653
rect 204976 221641 204982 221653
rect 205034 221641 205040 221693
rect 164080 221567 164086 221619
rect 164138 221607 164144 221619
rect 205360 221607 205366 221619
rect 164138 221579 205366 221607
rect 164138 221567 164144 221579
rect 205360 221567 205366 221579
rect 205418 221567 205424 221619
rect 166960 221493 166966 221545
rect 167018 221533 167024 221545
rect 206896 221533 206902 221545
rect 167018 221505 206902 221533
rect 167018 221493 167024 221505
rect 206896 221493 206902 221505
rect 206954 221493 206960 221545
rect 169840 221419 169846 221471
rect 169898 221459 169904 221471
rect 204592 221459 204598 221471
rect 169898 221431 204598 221459
rect 169898 221419 169904 221431
rect 204592 221419 204598 221431
rect 204650 221419 204656 221471
rect 42352 221049 42358 221101
rect 42410 221089 42416 221101
rect 44944 221089 44950 221101
rect 42410 221061 44950 221089
rect 42410 221049 42416 221061
rect 44944 221049 44950 221061
rect 45002 221049 45008 221101
rect 42352 220309 42358 220361
rect 42410 220349 42416 220361
rect 45136 220349 45142 220361
rect 42410 220321 45142 220349
rect 42410 220309 42416 220321
rect 45136 220309 45142 220321
rect 45194 220309 45200 220361
rect 42352 219421 42358 219473
rect 42410 219461 42416 219473
rect 44848 219461 44854 219473
rect 42410 219433 44854 219461
rect 42410 219421 42416 219433
rect 44848 219421 44854 219433
rect 44906 219421 44912 219473
rect 144016 218903 144022 218955
rect 144074 218943 144080 218955
rect 177136 218943 177142 218955
rect 144074 218915 177142 218943
rect 144074 218903 144080 218915
rect 177136 218903 177142 218915
rect 177194 218903 177200 218955
rect 175600 218829 175606 218881
rect 175658 218869 175664 218881
rect 204496 218869 204502 218881
rect 175658 218841 204502 218869
rect 175658 218829 175664 218841
rect 204496 218829 204502 218841
rect 204554 218829 204560 218881
rect 178480 218755 178486 218807
rect 178538 218795 178544 218807
rect 204592 218795 204598 218807
rect 178538 218767 204598 218795
rect 178538 218755 178544 218767
rect 204592 218755 204598 218767
rect 204650 218755 204656 218807
rect 181360 218681 181366 218733
rect 181418 218721 181424 218733
rect 204688 218721 204694 218733
rect 181418 218693 204694 218721
rect 181418 218681 181424 218693
rect 204688 218681 204694 218693
rect 204746 218681 204752 218733
rect 184240 218607 184246 218659
rect 184298 218647 184304 218659
rect 205360 218647 205366 218659
rect 184298 218619 205366 218647
rect 184298 218607 184304 218619
rect 205360 218607 205366 218619
rect 205418 218607 205424 218659
rect 146512 217719 146518 217771
rect 146570 217719 146576 217771
rect 146530 217623 146558 217719
rect 146512 217571 146518 217623
rect 146570 217571 146576 217623
rect 144016 216017 144022 216069
rect 144074 216057 144080 216069
rect 174256 216057 174262 216069
rect 144074 216029 174262 216057
rect 144074 216017 144080 216029
rect 174256 216017 174262 216029
rect 174314 216017 174320 216069
rect 187120 215943 187126 215995
rect 187178 215983 187184 215995
rect 204784 215983 204790 215995
rect 187178 215955 204790 215983
rect 187178 215943 187184 215955
rect 204784 215943 204790 215955
rect 204842 215943 204848 215995
rect 192880 215869 192886 215921
rect 192938 215909 192944 215921
rect 204496 215909 204502 215921
rect 192938 215881 204502 215909
rect 192938 215869 192944 215881
rect 204496 215869 204502 215881
rect 204554 215869 204560 215921
rect 146416 213427 146422 213479
rect 146474 213467 146480 213479
rect 146704 213467 146710 213479
rect 146474 213439 146710 213467
rect 146474 213427 146480 213439
rect 146704 213427 146710 213439
rect 146762 213427 146768 213479
rect 146416 213279 146422 213331
rect 146474 213319 146480 213331
rect 171376 213319 171382 213331
rect 146474 213291 171382 213319
rect 146474 213279 146480 213291
rect 171376 213279 171382 213291
rect 171434 213279 171440 213331
rect 144112 213205 144118 213257
rect 144170 213245 144176 213257
rect 154000 213245 154006 213257
rect 144170 213217 154006 213245
rect 144170 213205 144176 213217
rect 154000 213205 154006 213217
rect 154058 213205 154064 213257
rect 144016 213131 144022 213183
rect 144074 213171 144080 213183
rect 148240 213171 148246 213183
rect 144074 213143 148246 213171
rect 144074 213131 144080 213143
rect 148240 213131 148246 213143
rect 148298 213131 148304 213183
rect 205552 213131 205558 213183
rect 205610 213171 205616 213183
rect 207184 213171 207190 213183
rect 205610 213143 207190 213171
rect 205610 213131 205616 213143
rect 207184 213131 207190 213143
rect 207242 213131 207248 213183
rect 679792 212243 679798 212295
rect 679850 212283 679856 212295
rect 680080 212283 680086 212295
rect 679850 212255 680086 212283
rect 679850 212243 679856 212255
rect 680080 212243 680086 212255
rect 680138 212243 680144 212295
rect 146224 211577 146230 211629
rect 146282 211617 146288 211629
rect 146512 211617 146518 211629
rect 146282 211589 146518 211617
rect 146282 211577 146288 211589
rect 146512 211577 146518 211589
rect 146570 211577 146576 211629
rect 647920 210245 647926 210297
rect 647978 210285 647984 210297
rect 679792 210285 679798 210297
rect 647978 210257 679798 210285
rect 647978 210245 647984 210257
rect 679792 210245 679798 210257
rect 679850 210245 679856 210297
rect 144016 207433 144022 207485
rect 144074 207473 144080 207485
rect 165616 207473 165622 207485
rect 144074 207445 165622 207473
rect 144074 207433 144080 207445
rect 165616 207433 165622 207445
rect 165674 207433 165680 207485
rect 144112 207359 144118 207411
rect 144170 207399 144176 207411
rect 168496 207399 168502 207411
rect 144170 207371 168502 207399
rect 144170 207359 144176 207371
rect 168496 207359 168502 207371
rect 168554 207359 168560 207411
rect 674608 207359 674614 207411
rect 674666 207399 674672 207411
rect 676816 207399 676822 207411
rect 674666 207371 676822 207399
rect 674666 207359 674672 207371
rect 676816 207359 676822 207371
rect 676874 207359 676880 207411
rect 674416 205731 674422 205783
rect 674474 205771 674480 205783
rect 675472 205771 675478 205783
rect 674474 205743 675478 205771
rect 674474 205731 674480 205743
rect 675472 205731 675478 205743
rect 675530 205731 675536 205783
rect 675184 205139 675190 205191
rect 675242 205179 675248 205191
rect 675472 205179 675478 205191
rect 675242 205151 675478 205179
rect 675242 205139 675248 205151
rect 675472 205139 675478 205151
rect 675530 205139 675536 205191
rect 42352 204473 42358 204525
rect 42410 204513 42416 204525
rect 43024 204513 43030 204525
rect 42410 204485 43030 204513
rect 42410 204473 42416 204485
rect 43024 204473 43030 204485
rect 43082 204473 43088 204525
rect 144016 204473 144022 204525
rect 144074 204513 144080 204525
rect 148432 204513 148438 204525
rect 144074 204485 148438 204513
rect 144074 204473 144080 204485
rect 148432 204473 148438 204485
rect 148490 204473 148496 204525
rect 673936 204399 673942 204451
rect 673994 204439 674000 204451
rect 675376 204439 675382 204451
rect 673994 204411 675382 204439
rect 673994 204399 674000 204411
rect 675376 204399 675382 204411
rect 675434 204399 675440 204451
rect 42352 204325 42358 204377
rect 42410 204365 42416 204377
rect 44560 204365 44566 204377
rect 42410 204337 44566 204365
rect 42410 204325 42416 204337
rect 44560 204325 44566 204337
rect 44618 204325 44624 204377
rect 674992 202179 674998 202231
rect 675050 202219 675056 202231
rect 675280 202219 675286 202231
rect 675050 202191 675286 202219
rect 675050 202179 675056 202191
rect 675280 202179 675286 202191
rect 675338 202179 675344 202231
rect 675088 202031 675094 202083
rect 675146 202071 675152 202083
rect 675280 202071 675286 202083
rect 675146 202043 675286 202071
rect 675146 202031 675152 202043
rect 675280 202031 675286 202043
rect 675338 202031 675344 202083
rect 144016 201587 144022 201639
rect 144074 201627 144080 201639
rect 197200 201627 197206 201639
rect 144074 201599 197206 201627
rect 144074 201587 144080 201599
rect 197200 201587 197206 201599
rect 197258 201587 197264 201639
rect 40240 201513 40246 201565
rect 40298 201553 40304 201565
rect 41776 201553 41782 201565
rect 40298 201525 41782 201553
rect 40298 201513 40304 201525
rect 41776 201513 41782 201525
rect 41834 201513 41840 201565
rect 40048 201439 40054 201491
rect 40106 201479 40112 201491
rect 42160 201479 42166 201491
rect 40106 201451 42166 201479
rect 40106 201439 40112 201451
rect 42160 201439 42166 201451
rect 42218 201439 42224 201491
rect 674032 201291 674038 201343
rect 674090 201331 674096 201343
rect 675376 201331 675382 201343
rect 674090 201303 675382 201331
rect 674090 201291 674096 201303
rect 675376 201291 675382 201303
rect 675434 201291 675440 201343
rect 41968 201069 41974 201121
rect 42026 201109 42032 201121
rect 42352 201109 42358 201121
rect 42026 201081 42358 201109
rect 42026 201069 42032 201081
rect 42352 201069 42358 201081
rect 42410 201069 42416 201121
rect 674896 200847 674902 200899
rect 674954 200887 674960 200899
rect 675376 200887 675382 200899
rect 674954 200859 675382 200887
rect 674954 200847 674960 200859
rect 675376 200847 675382 200859
rect 675434 200847 675440 200899
rect 144112 198849 144118 198901
rect 144170 198889 144176 198901
rect 188560 198889 188566 198901
rect 144170 198861 188566 198889
rect 144170 198849 144176 198861
rect 188560 198849 188566 198861
rect 188618 198849 188624 198901
rect 37360 198775 37366 198827
rect 37418 198815 37424 198827
rect 43216 198815 43222 198827
rect 37418 198787 43222 198815
rect 37418 198775 37424 198787
rect 43216 198775 43222 198787
rect 43274 198775 43280 198827
rect 144016 198775 144022 198827
rect 144074 198815 144080 198827
rect 191440 198815 191446 198827
rect 144074 198787 191446 198815
rect 144074 198775 144080 198787
rect 191440 198775 191446 198787
rect 191498 198775 191504 198827
rect 40144 198701 40150 198753
rect 40202 198741 40208 198753
rect 40912 198741 40918 198753
rect 40202 198713 40918 198741
rect 40202 198701 40208 198713
rect 40912 198701 40918 198713
rect 40970 198701 40976 198753
rect 146224 198701 146230 198753
rect 146282 198741 146288 198753
rect 194320 198741 194326 198753
rect 146282 198713 194326 198741
rect 146282 198701 146288 198713
rect 194320 198701 194326 198713
rect 194378 198701 194384 198753
rect 674800 197591 674806 197643
rect 674858 197631 674864 197643
rect 675376 197631 675382 197643
rect 674858 197603 675382 197631
rect 674858 197591 674864 197603
rect 675376 197591 675382 197603
rect 675434 197591 675440 197643
rect 42064 197443 42070 197495
rect 42122 197483 42128 197495
rect 42928 197483 42934 197495
rect 42122 197455 42934 197483
rect 42122 197443 42128 197455
rect 42928 197443 42934 197455
rect 42986 197443 42992 197495
rect 41776 197369 41782 197421
rect 41834 197369 41840 197421
rect 41794 197199 41822 197369
rect 41776 197147 41782 197199
rect 41834 197147 41840 197199
rect 674608 196999 674614 197051
rect 674666 197039 674672 197051
rect 675472 197039 675478 197051
rect 674666 197011 675478 197039
rect 674666 196999 674672 197011
rect 675472 196999 675478 197011
rect 675530 196999 675536 197051
rect 674704 196555 674710 196607
rect 674762 196595 674768 196607
rect 675376 196595 675382 196607
rect 674762 196567 675382 196595
rect 674762 196555 674768 196567
rect 675376 196555 675382 196567
rect 675434 196555 675440 196607
rect 144016 195815 144022 195867
rect 144074 195855 144080 195867
rect 185680 195855 185686 195867
rect 144074 195827 185686 195855
rect 144074 195815 144080 195827
rect 185680 195815 185686 195827
rect 185738 195815 185744 195867
rect 42544 195741 42550 195793
rect 42602 195781 42608 195793
rect 42832 195781 42838 195793
rect 42602 195753 42838 195781
rect 42602 195741 42608 195753
rect 42832 195741 42838 195753
rect 42890 195741 42896 195793
rect 42832 195593 42838 195645
rect 42890 195633 42896 195645
rect 43216 195633 43222 195645
rect 42890 195605 43222 195633
rect 42890 195593 42896 195605
rect 43216 195593 43222 195605
rect 43274 195593 43280 195645
rect 42160 195297 42166 195349
rect 42218 195337 42224 195349
rect 42352 195337 42358 195349
rect 42218 195309 42358 195337
rect 42218 195297 42224 195309
rect 42352 195297 42358 195309
rect 42410 195297 42416 195349
rect 42064 194483 42070 194535
rect 42122 194523 42128 194535
rect 50416 194523 50422 194535
rect 42122 194495 50422 194523
rect 42122 194483 42128 194495
rect 50416 194483 50422 194495
rect 50474 194483 50480 194535
rect 42064 193447 42070 193499
rect 42122 193487 42128 193499
rect 43024 193487 43030 193499
rect 42122 193459 43030 193487
rect 42122 193447 42128 193459
rect 43024 193447 43030 193459
rect 43082 193447 43088 193499
rect 42160 192189 42166 192241
rect 42218 192229 42224 192241
rect 43120 192229 43126 192241
rect 42218 192201 43126 192229
rect 42218 192189 42224 192201
rect 43120 192189 43126 192201
rect 43178 192189 43184 192241
rect 42064 191449 42070 191501
rect 42122 191489 42128 191501
rect 42352 191489 42358 191501
rect 42122 191461 42358 191489
rect 42122 191449 42128 191461
rect 42352 191449 42358 191461
rect 42410 191449 42416 191501
rect 144016 190117 144022 190169
rect 144074 190157 144080 190169
rect 151216 190157 151222 190169
rect 144074 190129 151222 190157
rect 144074 190117 144080 190129
rect 151216 190117 151222 190129
rect 151274 190117 151280 190169
rect 204880 190117 204886 190169
rect 204938 190157 204944 190169
rect 205072 190157 205078 190169
rect 204938 190129 205078 190157
rect 204938 190117 204944 190129
rect 205072 190117 205078 190129
rect 205130 190117 205136 190169
rect 42160 187675 42166 187727
rect 42218 187715 42224 187727
rect 42832 187715 42838 187727
rect 42218 187687 42838 187715
rect 42218 187675 42224 187687
rect 42832 187675 42838 187687
rect 42890 187675 42896 187727
rect 42928 187271 42934 187283
rect 42370 187243 42934 187271
rect 42256 187157 42262 187209
rect 42314 187197 42320 187209
rect 42370 187197 42398 187243
rect 42928 187231 42934 187243
rect 42986 187231 42992 187283
rect 146416 187231 146422 187283
rect 146474 187271 146480 187283
rect 197296 187271 197302 187283
rect 146474 187243 197302 187271
rect 146474 187231 146480 187243
rect 197296 187231 197302 187243
rect 197354 187231 197360 187283
rect 42314 187169 42398 187197
rect 42314 187157 42320 187169
rect 204880 187157 204886 187209
rect 204938 187197 204944 187209
rect 205072 187197 205078 187209
rect 204938 187169 205078 187197
rect 204938 187157 204944 187169
rect 205072 187157 205078 187169
rect 205130 187157 205136 187209
rect 206992 187157 206998 187209
rect 207050 187197 207056 187209
rect 207280 187197 207286 187209
rect 207050 187169 207286 187197
rect 207050 187157 207056 187169
rect 207280 187157 207286 187169
rect 207338 187157 207344 187209
rect 42160 187083 42166 187135
rect 42218 187123 42224 187135
rect 42544 187123 42550 187135
rect 42218 187095 42550 187123
rect 42218 187083 42224 187095
rect 42544 187083 42550 187095
rect 42602 187083 42608 187135
rect 144496 184419 144502 184471
rect 144554 184459 144560 184471
rect 148528 184459 148534 184471
rect 144554 184431 148534 184459
rect 144554 184419 144560 184431
rect 148528 184419 148534 184431
rect 148586 184419 148592 184471
rect 146800 184345 146806 184397
rect 146858 184385 146864 184397
rect 194416 184385 194422 184397
rect 146858 184357 194422 184385
rect 146858 184345 146864 184357
rect 194416 184345 194422 184357
rect 194474 184345 194480 184397
rect 655312 184345 655318 184397
rect 655370 184385 655376 184397
rect 674416 184385 674422 184397
rect 655370 184357 674422 184385
rect 655370 184345 655376 184357
rect 674416 184345 674422 184357
rect 674474 184345 674480 184397
rect 660976 183901 660982 183953
rect 661034 183941 661040 183953
rect 674704 183941 674710 183953
rect 661034 183913 674710 183941
rect 661034 183901 661040 183913
rect 674704 183901 674710 183913
rect 674762 183901 674768 183953
rect 666736 182865 666742 182917
rect 666794 182905 666800 182917
rect 674416 182905 674422 182917
rect 666794 182877 674422 182905
rect 666794 182865 666800 182877
rect 674416 182865 674422 182877
rect 674474 182865 674480 182917
rect 146800 181459 146806 181511
rect 146858 181499 146864 181511
rect 188656 181499 188662 181511
rect 146858 181471 188662 181499
rect 146858 181459 146864 181471
rect 188656 181459 188662 181471
rect 188714 181459 188720 181511
rect 145264 178647 145270 178699
rect 145322 178687 145328 178699
rect 148624 178687 148630 178699
rect 145322 178659 148630 178687
rect 145322 178647 145328 178659
rect 148624 178647 148630 178659
rect 148682 178647 148688 178699
rect 146800 178573 146806 178625
rect 146858 178613 146864 178625
rect 191536 178613 191542 178625
rect 146858 178585 191542 178613
rect 146858 178573 146864 178585
rect 191536 178573 191542 178585
rect 191594 178573 191600 178625
rect 146800 175687 146806 175739
rect 146858 175727 146864 175739
rect 185776 175727 185782 175739
rect 146858 175699 185782 175727
rect 146858 175687 146864 175699
rect 185776 175687 185782 175699
rect 185834 175687 185840 175739
rect 144016 175613 144022 175665
rect 144074 175653 144080 175665
rect 146512 175653 146518 175665
rect 144074 175625 146518 175653
rect 144074 175613 144080 175625
rect 146512 175613 146518 175625
rect 146570 175613 146576 175665
rect 146800 172801 146806 172853
rect 146858 172841 146864 172853
rect 162736 172841 162742 172853
rect 146858 172813 162742 172841
rect 146858 172801 146864 172813
rect 162736 172801 162742 172813
rect 162794 172801 162800 172853
rect 146800 171247 146806 171299
rect 146858 171287 146864 171299
rect 159856 171287 159862 171299
rect 146858 171259 159862 171287
rect 146858 171247 146864 171259
rect 159856 171247 159862 171259
rect 159914 171247 159920 171299
rect 146800 167251 146806 167303
rect 146858 167291 146864 167303
rect 156976 167291 156982 167303
rect 146858 167263 156982 167291
rect 146858 167251 146864 167263
rect 156976 167251 156982 167263
rect 157034 167251 157040 167303
rect 647056 167177 647062 167229
rect 647114 167217 647120 167229
rect 674704 167217 674710 167229
rect 647114 167189 674710 167217
rect 647114 167177 647120 167189
rect 674704 167177 674710 167189
rect 674762 167177 674768 167229
rect 144016 166659 144022 166711
rect 144074 166699 144080 166711
rect 146512 166699 146518 166711
rect 144074 166671 146518 166699
rect 144074 166659 144080 166671
rect 146512 166659 146518 166671
rect 146570 166659 146576 166711
rect 646288 164217 646294 164269
rect 646346 164257 646352 164269
rect 674608 164257 674614 164269
rect 646346 164229 674614 164257
rect 646346 164217 646352 164229
rect 674608 164217 674614 164229
rect 674666 164217 674672 164269
rect 144016 164143 144022 164195
rect 144074 164183 144080 164195
rect 208720 164183 208726 164195
rect 144074 164155 208726 164183
rect 144074 164143 144080 164155
rect 208720 164143 208726 164155
rect 208778 164143 208784 164195
rect 647920 164143 647926 164195
rect 647978 164183 647984 164195
rect 674704 164183 674710 164195
rect 647978 164155 674710 164183
rect 647978 164143 647984 164155
rect 674704 164143 674710 164155
rect 674762 164143 674768 164195
rect 144688 163699 144694 163751
rect 144746 163739 144752 163751
rect 146800 163739 146806 163751
rect 144746 163711 146806 163739
rect 144746 163699 144752 163711
rect 146800 163699 146806 163711
rect 146858 163699 146864 163751
rect 674704 163625 674710 163677
rect 674762 163665 674768 163677
rect 677104 163665 677110 163677
rect 674762 163637 677110 163665
rect 674762 163625 674768 163637
rect 677104 163625 677110 163637
rect 677162 163625 677168 163677
rect 674800 163255 674806 163307
rect 674858 163295 674864 163307
rect 676816 163295 676822 163307
rect 674858 163267 676822 163295
rect 674858 163255 674864 163267
rect 676816 163255 676822 163267
rect 676874 163255 676880 163307
rect 206992 162885 206998 162937
rect 207050 162925 207056 162937
rect 207376 162925 207382 162937
rect 207050 162897 207382 162925
rect 207050 162885 207056 162897
rect 207376 162885 207382 162897
rect 207434 162885 207440 162937
rect 144016 161257 144022 161309
rect 144074 161297 144080 161309
rect 148720 161297 148726 161309
rect 144074 161269 148726 161297
rect 144074 161257 144080 161269
rect 148720 161257 148726 161269
rect 148778 161257 148784 161309
rect 674896 160739 674902 160791
rect 674954 160779 674960 160791
rect 675376 160779 675382 160791
rect 674954 160751 675382 160779
rect 674954 160739 674960 160751
rect 675376 160739 675382 160751
rect 675434 160739 675440 160791
rect 674992 159999 674998 160051
rect 675050 160039 675056 160051
rect 675472 160039 675478 160051
rect 675050 160011 675478 160039
rect 675050 159999 675056 160011
rect 675472 159999 675478 160011
rect 675530 159999 675536 160051
rect 144016 158445 144022 158497
rect 144074 158485 144080 158497
rect 148816 158485 148822 158497
rect 144074 158457 148822 158485
rect 144074 158445 144080 158457
rect 148816 158445 148822 158457
rect 148874 158445 148880 158497
rect 674512 157705 674518 157757
rect 674570 157745 674576 157757
rect 675184 157745 675190 157757
rect 674570 157717 675190 157745
rect 674570 157705 674576 157717
rect 675184 157705 675190 157717
rect 675242 157705 675248 157757
rect 674608 156891 674614 156943
rect 674666 156931 674672 156943
rect 675472 156931 675478 156943
rect 674666 156903 675478 156931
rect 674666 156891 674672 156903
rect 675472 156891 675478 156903
rect 675530 156891 675536 156943
rect 144016 155707 144022 155759
rect 144074 155747 144080 155759
rect 148912 155747 148918 155759
rect 144074 155719 148918 155747
rect 144074 155707 144080 155719
rect 148912 155707 148918 155719
rect 148970 155707 148976 155759
rect 144112 155633 144118 155685
rect 144170 155673 144176 155685
rect 200176 155673 200182 155685
rect 144170 155645 200182 155673
rect 144170 155633 144176 155645
rect 200176 155633 200182 155645
rect 200234 155633 200240 155685
rect 144208 155559 144214 155611
rect 144266 155599 144272 155611
rect 203056 155599 203062 155611
rect 144266 155571 203062 155599
rect 144266 155559 144272 155571
rect 203056 155559 203062 155571
rect 203114 155559 203120 155611
rect 144016 152747 144022 152799
rect 144074 152787 144080 152799
rect 180016 152787 180022 152799
rect 144074 152759 180022 152787
rect 144074 152747 144080 152759
rect 180016 152747 180022 152759
rect 180074 152747 180080 152799
rect 144112 152673 144118 152725
rect 144170 152713 144176 152725
rect 182896 152713 182902 152725
rect 144170 152685 182902 152713
rect 144170 152673 144176 152685
rect 182896 152673 182902 152685
rect 182954 152673 182960 152725
rect 674224 152599 674230 152651
rect 674282 152639 674288 152651
rect 675376 152639 675382 152651
rect 674282 152611 675382 152639
rect 674282 152599 674288 152611
rect 675376 152599 675382 152611
rect 675434 152599 675440 152651
rect 674800 152155 674806 152207
rect 674858 152195 674864 152207
rect 675472 152195 675478 152207
rect 674858 152167 675478 152195
rect 674858 152155 674864 152167
rect 675472 152155 675478 152167
rect 675530 152155 675536 152207
rect 674128 151415 674134 151467
rect 674186 151455 674192 151467
rect 675376 151455 675382 151467
rect 674186 151427 675382 151455
rect 674186 151415 674192 151427
rect 675376 151415 675382 151427
rect 675434 151415 675440 151467
rect 674704 150305 674710 150357
rect 674762 150345 674768 150357
rect 675472 150345 675478 150357
rect 674762 150317 675478 150345
rect 674762 150305 674768 150317
rect 675472 150305 675478 150317
rect 675530 150305 675536 150357
rect 144112 149861 144118 149913
rect 144170 149901 144176 149913
rect 149008 149901 149014 149913
rect 144170 149873 149014 149901
rect 144170 149861 144176 149873
rect 149008 149861 149014 149873
rect 149066 149861 149072 149913
rect 144016 149787 144022 149839
rect 144074 149827 144080 149839
rect 177232 149827 177238 149839
rect 144074 149799 177238 149827
rect 144074 149787 144080 149799
rect 177232 149787 177238 149799
rect 177290 149787 177296 149839
rect 144016 149639 144022 149691
rect 144074 149679 144080 149691
rect 144496 149679 144502 149691
rect 144074 149651 144502 149679
rect 144074 149639 144080 149651
rect 144496 149639 144502 149651
rect 144554 149639 144560 149691
rect 144688 147237 144694 147249
rect 143938 147209 144694 147237
rect 143938 146941 143966 147209
rect 144688 147197 144694 147209
rect 144746 147197 144752 147249
rect 144016 147123 144022 147175
rect 144074 147163 144080 147175
rect 144074 147135 144734 147163
rect 144074 147123 144080 147135
rect 144706 147101 144734 147135
rect 144688 147049 144694 147101
rect 144746 147049 144752 147101
rect 144112 146941 144118 146953
rect 143938 146913 144118 146941
rect 144112 146901 144118 146913
rect 144170 146901 144176 146953
rect 144496 146901 144502 146953
rect 144554 146941 144560 146953
rect 174352 146941 174358 146953
rect 144554 146913 174358 146941
rect 144554 146901 144560 146913
rect 174352 146901 174358 146913
rect 174410 146901 174416 146953
rect 144496 146235 144502 146287
rect 144554 146275 144560 146287
rect 146320 146275 146326 146287
rect 144554 146247 146326 146275
rect 144554 146235 144560 146247
rect 146320 146235 146326 146247
rect 146378 146235 146384 146287
rect 144208 146087 144214 146139
rect 144266 146127 144272 146139
rect 146320 146127 146326 146139
rect 144266 146099 146326 146127
rect 144266 146087 144272 146099
rect 146320 146087 146326 146099
rect 146378 146087 146384 146139
rect 144208 144311 144214 144363
rect 144266 144351 144272 144363
rect 154096 144351 154102 144363
rect 144266 144323 154102 144351
rect 144266 144311 144272 144323
rect 154096 144311 154102 144323
rect 154154 144311 154160 144363
rect 144208 144015 144214 144067
rect 144266 144055 144272 144067
rect 208816 144055 208822 144067
rect 144266 144027 208822 144055
rect 144266 144015 144272 144027
rect 208816 144015 208822 144027
rect 208874 144015 208880 144067
rect 144208 142535 144214 142587
rect 144266 142575 144272 142587
rect 149200 142575 149206 142587
rect 144266 142547 149206 142575
rect 144266 142535 144272 142547
rect 149200 142535 149206 142547
rect 149258 142535 149264 142587
rect 144208 141129 144214 141181
rect 144266 141169 144272 141181
rect 171472 141169 171478 141181
rect 144266 141141 171478 141169
rect 144266 141129 144272 141141
rect 171472 141129 171478 141141
rect 171530 141129 171536 141181
rect 144208 140833 144214 140885
rect 144266 140873 144272 140885
rect 144496 140873 144502 140885
rect 144266 140845 144502 140873
rect 144266 140833 144272 140845
rect 144496 140833 144502 140845
rect 144554 140833 144560 140885
rect 655216 138539 655222 138591
rect 655274 138579 655280 138591
rect 674704 138579 674710 138591
rect 655274 138551 674710 138579
rect 655274 138539 655280 138551
rect 674704 138539 674710 138551
rect 674762 138539 674768 138591
rect 655120 138391 655126 138443
rect 655178 138431 655184 138443
rect 674416 138431 674422 138443
rect 655178 138403 674422 138431
rect 655178 138391 655184 138403
rect 674416 138391 674422 138403
rect 674474 138391 674480 138443
rect 144496 138317 144502 138369
rect 144554 138357 144560 138369
rect 168592 138357 168598 138369
rect 144554 138329 168598 138357
rect 144554 138317 144560 138329
rect 168592 138317 168598 138329
rect 168650 138317 168656 138369
rect 143824 138243 143830 138295
rect 143882 138283 143888 138295
rect 208912 138283 208918 138295
rect 143882 138255 208918 138283
rect 143882 138243 143888 138255
rect 208912 138243 208918 138255
rect 208970 138243 208976 138295
rect 143920 138169 143926 138221
rect 143978 138209 143984 138221
rect 144496 138209 144502 138221
rect 143978 138181 144502 138209
rect 143978 138169 143984 138181
rect 144496 138169 144502 138181
rect 144554 138169 144560 138221
rect 144688 136911 144694 136963
rect 144746 136951 144752 136963
rect 144746 136923 144830 136951
rect 144746 136911 144752 136923
rect 144802 136741 144830 136923
rect 144784 136689 144790 136741
rect 144842 136689 144848 136741
rect 146896 136245 146902 136297
rect 146954 136285 146960 136297
rect 149296 136285 149302 136297
rect 146954 136257 149302 136285
rect 146954 136245 146960 136257
rect 149296 136245 149302 136257
rect 149354 136245 149360 136297
rect 146896 135949 146902 136001
rect 146954 135989 146960 136001
rect 149392 135989 149398 136001
rect 146954 135961 149398 135989
rect 146954 135949 146960 135961
rect 149392 135949 149398 135961
rect 149450 135949 149456 136001
rect 655408 135579 655414 135631
rect 655466 135619 655472 135631
rect 674608 135619 674614 135631
rect 655466 135591 674614 135619
rect 655466 135579 655472 135591
rect 674608 135579 674614 135591
rect 674666 135579 674672 135631
rect 646480 135357 646486 135409
rect 646538 135397 646544 135409
rect 674704 135397 674710 135409
rect 646538 135369 674710 135397
rect 646538 135357 646544 135369
rect 674704 135357 674710 135369
rect 674762 135357 674768 135409
rect 144208 134839 144214 134891
rect 144266 134879 144272 134891
rect 146992 134879 146998 134891
rect 144266 134851 146998 134879
rect 144266 134839 144272 134851
rect 146992 134839 146998 134851
rect 147050 134839 147056 134891
rect 146704 134543 146710 134595
rect 146762 134543 146768 134595
rect 146722 134361 146750 134543
rect 146800 134361 146806 134373
rect 146722 134333 146806 134361
rect 146800 134321 146806 134333
rect 146858 134321 146864 134373
rect 144208 134173 144214 134225
rect 144266 134213 144272 134225
rect 146800 134213 146806 134225
rect 144266 134185 146806 134213
rect 144266 134173 144272 134185
rect 146800 134173 146806 134185
rect 146858 134173 146864 134225
rect 144496 132915 144502 132967
rect 144554 132915 144560 132967
rect 144514 132807 144542 132915
rect 144130 132779 144542 132807
rect 144130 132585 144158 132779
rect 144208 132693 144214 132745
rect 144266 132733 144272 132745
rect 209104 132733 209110 132745
rect 144266 132705 209110 132733
rect 144266 132693 144272 132705
rect 209104 132693 209110 132705
rect 209162 132693 209168 132745
rect 146800 132619 146806 132671
rect 146858 132659 146864 132671
rect 165712 132659 165718 132671
rect 146858 132631 165718 132659
rect 146858 132619 146864 132631
rect 165712 132619 165718 132631
rect 165770 132619 165776 132671
rect 144208 132585 144214 132597
rect 144130 132557 144214 132585
rect 144208 132545 144214 132557
rect 144266 132545 144272 132597
rect 144496 132545 144502 132597
rect 144554 132585 144560 132597
rect 209008 132585 209014 132597
rect 144554 132557 209014 132585
rect 144554 132545 144560 132557
rect 209008 132545 209014 132557
rect 209066 132545 209072 132597
rect 143920 130103 143926 130155
rect 143978 130143 143984 130155
rect 144208 130143 144214 130155
rect 143978 130115 144214 130143
rect 143978 130103 143984 130115
rect 144208 130103 144214 130115
rect 144266 130103 144272 130155
rect 144496 129659 144502 129711
rect 144554 129699 144560 129711
rect 151408 129699 151414 129711
rect 144554 129671 151414 129699
rect 144554 129659 144560 129671
rect 151408 129659 151414 129671
rect 151466 129659 151472 129711
rect 144208 129585 144214 129637
rect 144266 129625 144272 129637
rect 209200 129625 209206 129637
rect 144266 129597 209206 129625
rect 144266 129585 144272 129597
rect 209200 129585 209206 129597
rect 209258 129585 209264 129637
rect 144496 129511 144502 129563
rect 144554 129551 144560 129563
rect 146320 129551 146326 129563
rect 144554 129523 146326 129551
rect 144554 129511 144560 129523
rect 146320 129511 146326 129523
rect 146378 129511 146384 129563
rect 147088 126847 147094 126899
rect 147146 126887 147152 126899
rect 149488 126887 149494 126899
rect 147146 126859 149494 126887
rect 147146 126847 147152 126859
rect 149488 126847 149494 126859
rect 149546 126847 149552 126899
rect 146704 126773 146710 126825
rect 146762 126813 146768 126825
rect 203152 126813 203158 126825
rect 146762 126785 203158 126813
rect 146762 126773 146768 126785
rect 203152 126773 203158 126785
rect 203210 126773 203216 126825
rect 143920 126699 143926 126751
rect 143978 126739 143984 126751
rect 144208 126739 144214 126751
rect 143978 126711 144214 126739
rect 143978 126699 143984 126711
rect 144208 126699 144214 126711
rect 144266 126699 144272 126751
rect 146320 126699 146326 126751
rect 146378 126739 146384 126751
rect 208624 126739 208630 126751
rect 146378 126711 208630 126739
rect 146378 126699 146384 126711
rect 208624 126699 208630 126711
rect 208682 126699 208688 126751
rect 204784 126625 204790 126677
rect 204842 126665 204848 126677
rect 204880 126665 204886 126677
rect 204842 126637 204886 126665
rect 204842 126625 204848 126637
rect 204880 126625 204886 126637
rect 204938 126625 204944 126677
rect 39856 125293 39862 125345
rect 39914 125333 39920 125345
rect 42448 125333 42454 125345
rect 39914 125305 42454 125333
rect 39914 125293 39920 125305
rect 42448 125293 42454 125305
rect 42506 125293 42512 125345
rect 146704 124035 146710 124087
rect 146762 124075 146768 124087
rect 197392 124075 197398 124087
rect 146762 124047 197398 124075
rect 146762 124035 146768 124047
rect 197392 124035 197398 124047
rect 197450 124035 197456 124087
rect 146320 123887 146326 123939
rect 146378 123927 146384 123939
rect 200272 123927 200278 123939
rect 146378 123899 200278 123927
rect 146378 123887 146384 123899
rect 200272 123887 200278 123899
rect 200330 123887 200336 123939
rect 146320 123739 146326 123791
rect 146378 123779 146384 123791
rect 146896 123779 146902 123791
rect 146378 123751 146902 123779
rect 146378 123739 146384 123751
rect 146896 123739 146902 123751
rect 146954 123739 146960 123791
rect 647824 121223 647830 121275
rect 647882 121263 647888 121275
rect 674704 121263 674710 121275
rect 647882 121235 674710 121263
rect 647882 121223 647888 121235
rect 674704 121223 674710 121235
rect 674762 121223 674768 121275
rect 647728 121149 647734 121201
rect 647786 121189 647792 121201
rect 674416 121189 674422 121201
rect 647786 121161 674422 121189
rect 647786 121149 647792 121161
rect 674416 121149 674422 121161
rect 674474 121149 674480 121201
rect 146896 121075 146902 121127
rect 146954 121115 146960 121127
rect 149584 121115 149590 121127
rect 146954 121087 149590 121115
rect 146954 121075 146960 121087
rect 149584 121075 149590 121087
rect 149642 121075 149648 121127
rect 647920 121075 647926 121127
rect 647978 121115 647984 121127
rect 674608 121115 674614 121127
rect 647978 121087 674614 121115
rect 647978 121075 647984 121087
rect 674608 121075 674614 121087
rect 674666 121075 674672 121127
rect 146704 121001 146710 121053
rect 146762 121041 146768 121053
rect 208528 121041 208534 121053
rect 146762 121013 208534 121041
rect 146762 121001 146768 121013
rect 208528 121001 208534 121013
rect 208586 121001 208592 121053
rect 146320 119151 146326 119203
rect 146378 119151 146384 119203
rect 146338 118229 146366 119151
rect 146704 118559 146710 118611
rect 146762 118599 146768 118611
rect 194512 118599 194518 118611
rect 146762 118571 194518 118599
rect 146762 118559 146768 118571
rect 194512 118559 194518 118571
rect 194570 118559 194576 118611
rect 146704 118263 146710 118315
rect 146762 118303 146768 118315
rect 188752 118303 188758 118315
rect 146762 118275 188758 118303
rect 146762 118263 146768 118275
rect 188752 118263 188758 118275
rect 188810 118263 188816 118315
rect 146242 118201 146366 118229
rect 146242 118007 146270 118201
rect 146320 118115 146326 118167
rect 146378 118155 146384 118167
rect 208432 118155 208438 118167
rect 146378 118127 208438 118155
rect 146378 118115 146384 118127
rect 208432 118115 208438 118127
rect 208490 118115 208496 118167
rect 674800 118041 674806 118093
rect 674858 118081 674864 118093
rect 676816 118081 676822 118093
rect 674858 118053 676822 118081
rect 674858 118041 674864 118053
rect 676816 118041 676822 118053
rect 676874 118041 676880 118093
rect 146320 118007 146326 118019
rect 146242 117979 146326 118007
rect 146320 117967 146326 117979
rect 146378 117967 146384 118019
rect 674704 117967 674710 118019
rect 674762 118007 674768 118019
rect 676912 118007 676918 118019
rect 674762 117979 676918 118007
rect 674762 117967 674768 117979
rect 676912 117967 676918 117979
rect 676970 117967 676976 118019
rect 675472 115747 675478 115799
rect 675530 115747 675536 115799
rect 675490 115577 675518 115747
rect 146896 115525 146902 115577
rect 146954 115565 146960 115577
rect 149680 115565 149686 115577
rect 146954 115537 149686 115565
rect 146954 115525 146960 115537
rect 149680 115525 149686 115537
rect 149738 115525 149744 115577
rect 675472 115525 675478 115577
rect 675530 115525 675536 115577
rect 146704 115229 146710 115281
rect 146762 115269 146768 115281
rect 208336 115269 208342 115281
rect 146762 115241 208342 115269
rect 146762 115229 146768 115241
rect 208336 115229 208342 115241
rect 208394 115229 208400 115281
rect 143824 115155 143830 115207
rect 143882 115195 143888 115207
rect 144304 115195 144310 115207
rect 143882 115167 144310 115195
rect 143882 115155 143888 115167
rect 144304 115155 144310 115167
rect 144362 115155 144368 115207
rect 144400 115155 144406 115207
rect 144458 115155 144464 115207
rect 144496 115155 144502 115207
rect 144554 115155 144560 115207
rect 146320 115195 146326 115207
rect 144610 115167 146326 115195
rect 143728 115081 143734 115133
rect 143786 115121 143792 115133
rect 144112 115121 144118 115133
rect 143786 115093 144118 115121
rect 143786 115081 143792 115093
rect 144112 115081 144118 115093
rect 144170 115081 144176 115133
rect 144112 114933 144118 114985
rect 144170 114973 144176 114985
rect 144418 114973 144446 115155
rect 144514 114985 144542 115155
rect 144610 114985 144638 115167
rect 146320 115155 146326 115167
rect 146378 115155 146384 115207
rect 146320 115007 146326 115059
rect 146378 115047 146384 115059
rect 146992 115047 146998 115059
rect 146378 115019 146998 115047
rect 146378 115007 146384 115019
rect 146992 115007 146998 115019
rect 147050 115007 147056 115059
rect 144170 114945 144446 114973
rect 144170 114933 144176 114945
rect 144496 114933 144502 114985
rect 144554 114933 144560 114985
rect 144592 114933 144598 114985
rect 144650 114933 144656 114985
rect 674608 114785 674614 114837
rect 674666 114825 674672 114837
rect 675376 114825 675382 114837
rect 674666 114797 675382 114825
rect 674666 114785 674672 114797
rect 675376 114785 675382 114797
rect 675434 114785 675440 114837
rect 146704 112639 146710 112691
rect 146762 112679 146768 112691
rect 191632 112679 191638 112691
rect 146762 112651 191638 112679
rect 146762 112639 146768 112651
rect 191632 112639 191638 112651
rect 191690 112639 191696 112691
rect 144400 112417 144406 112469
rect 144458 112457 144464 112469
rect 148144 112457 148150 112469
rect 144458 112429 148150 112457
rect 144458 112417 144464 112429
rect 148144 112417 148150 112429
rect 148202 112417 148208 112469
rect 146704 112343 146710 112395
rect 146762 112383 146768 112395
rect 148048 112383 148054 112395
rect 146762 112355 148054 112383
rect 146762 112343 146768 112355
rect 148048 112343 148054 112355
rect 148106 112343 148112 112395
rect 207184 112343 207190 112395
rect 207242 112383 207248 112395
rect 207376 112383 207382 112395
rect 207242 112355 207382 112383
rect 207242 112343 207248 112355
rect 207376 112343 207382 112355
rect 207434 112343 207440 112395
rect 674512 110937 674518 110989
rect 674570 110977 674576 110989
rect 675088 110977 675094 110989
rect 674570 110949 675094 110977
rect 674570 110937 674576 110949
rect 675088 110937 675094 110949
rect 675146 110937 675152 110989
rect 144400 109531 144406 109583
rect 144458 109571 144464 109583
rect 147952 109571 147958 109583
rect 144458 109543 147958 109571
rect 144458 109531 144464 109543
rect 147952 109531 147958 109543
rect 148010 109531 148016 109583
rect 146704 109457 146710 109509
rect 146762 109497 146768 109509
rect 185872 109497 185878 109509
rect 146762 109469 185878 109497
rect 146762 109457 146768 109469
rect 185872 109457 185878 109469
rect 185930 109457 185936 109509
rect 674320 107311 674326 107363
rect 674378 107351 674384 107363
rect 675376 107351 675382 107363
rect 674378 107323 675382 107351
rect 674378 107311 674384 107323
rect 675376 107311 675382 107323
rect 675434 107311 675440 107363
rect 674800 106941 674806 106993
rect 674858 106981 674864 106993
rect 675472 106981 675478 106993
rect 674858 106953 675478 106981
rect 674858 106941 674864 106953
rect 675472 106941 675478 106953
rect 675530 106941 675536 106993
rect 144400 106645 144406 106697
rect 144458 106685 144464 106697
rect 147856 106685 147862 106697
rect 144458 106657 147862 106685
rect 144458 106645 144464 106657
rect 147856 106645 147862 106657
rect 147914 106645 147920 106697
rect 146704 106571 146710 106623
rect 146762 106611 146768 106623
rect 162832 106611 162838 106623
rect 146762 106583 162838 106611
rect 146762 106571 146768 106583
rect 162832 106571 162838 106583
rect 162890 106571 162896 106623
rect 204784 106571 204790 106623
rect 204842 106611 204848 106623
rect 204976 106611 204982 106623
rect 204842 106583 204982 106611
rect 204842 106571 204848 106583
rect 204976 106571 204982 106583
rect 205034 106571 205040 106623
rect 143824 106497 143830 106549
rect 143882 106537 143888 106549
rect 143882 106509 146750 106537
rect 143882 106497 143888 106509
rect 146722 106475 146750 106509
rect 146704 106423 146710 106475
rect 146762 106423 146768 106475
rect 674128 106127 674134 106179
rect 674186 106167 674192 106179
rect 675376 106167 675382 106179
rect 674186 106139 675382 106167
rect 674186 106127 674192 106139
rect 675376 106127 675382 106139
rect 675434 106127 675440 106179
rect 674704 105165 674710 105217
rect 674762 105205 674768 105217
rect 675376 105205 675382 105217
rect 674762 105177 675382 105205
rect 674762 105165 674768 105177
rect 675376 105165 675382 105177
rect 675434 105165 675440 105217
rect 144016 104869 144022 104921
rect 144074 104869 144080 104921
rect 144034 104687 144062 104869
rect 146512 104795 146518 104847
rect 146570 104835 146576 104847
rect 146896 104835 146902 104847
rect 146570 104807 146902 104835
rect 146570 104795 146576 104807
rect 146896 104795 146902 104807
rect 146954 104795 146960 104847
rect 146512 104687 146518 104699
rect 144034 104659 146518 104687
rect 146512 104647 146518 104659
rect 146570 104647 146576 104699
rect 647920 104499 647926 104551
rect 647978 104539 647984 104551
rect 665200 104539 665206 104551
rect 647978 104511 665206 104539
rect 647978 104499 647984 104511
rect 665200 104499 665206 104511
rect 665258 104499 665264 104551
rect 144784 104203 144790 104255
rect 144842 104243 144848 104255
rect 159952 104243 159958 104255
rect 144842 104215 159958 104243
rect 144842 104203 144848 104215
rect 159952 104203 159958 104215
rect 160010 104203 160016 104255
rect 144304 103759 144310 103811
rect 144362 103799 144368 103811
rect 151312 103799 151318 103811
rect 144362 103771 151318 103799
rect 144362 103759 144368 103771
rect 151312 103759 151318 103771
rect 151370 103759 151376 103811
rect 144112 103685 144118 103737
rect 144170 103725 144176 103737
rect 208240 103725 208246 103737
rect 144170 103697 208246 103725
rect 144170 103685 144176 103697
rect 208240 103685 208246 103697
rect 208298 103685 208304 103737
rect 146896 103611 146902 103663
rect 146954 103651 146960 103663
rect 206704 103651 206710 103663
rect 146954 103623 206710 103651
rect 146954 103611 146960 103623
rect 206704 103611 206710 103623
rect 206762 103611 206768 103663
rect 146320 103537 146326 103589
rect 146378 103577 146384 103589
rect 204496 103577 204502 103589
rect 146378 103549 204502 103577
rect 146378 103537 146384 103549
rect 204496 103537 204502 103549
rect 204554 103537 204560 103589
rect 144592 103463 144598 103515
rect 144650 103503 144656 103515
rect 206224 103503 206230 103515
rect 144650 103475 206230 103503
rect 144650 103463 144656 103475
rect 206224 103463 206230 103475
rect 206282 103463 206288 103515
rect 143728 103315 143734 103367
rect 143786 103355 143792 103367
rect 144592 103355 144598 103367
rect 143786 103327 144598 103355
rect 143786 103315 143792 103327
rect 144592 103315 144598 103327
rect 144650 103315 144656 103367
rect 144016 101539 144022 101591
rect 144074 101579 144080 101591
rect 157072 101579 157078 101591
rect 144074 101551 157078 101579
rect 144074 101539 144080 101551
rect 157072 101539 157078 101551
rect 157130 101539 157136 101591
rect 144112 100799 144118 100851
rect 144170 100839 144176 100851
rect 147760 100839 147766 100851
rect 144170 100811 147766 100839
rect 144170 100799 144176 100811
rect 147760 100799 147766 100811
rect 147818 100799 147824 100851
rect 146704 100725 146710 100777
rect 146762 100765 146768 100777
rect 204688 100765 204694 100777
rect 146762 100737 204694 100765
rect 146762 100725 146768 100737
rect 204688 100725 204694 100737
rect 204746 100725 204752 100777
rect 144016 100651 144022 100703
rect 144074 100691 144080 100703
rect 206896 100691 206902 100703
rect 144074 100663 206902 100691
rect 144074 100651 144080 100663
rect 206896 100651 206902 100663
rect 206954 100651 206960 100703
rect 144400 100577 144406 100629
rect 144458 100617 144464 100629
rect 204592 100617 204598 100629
rect 144458 100589 204598 100617
rect 144458 100577 144464 100589
rect 204592 100577 204598 100589
rect 204650 100577 204656 100629
rect 151120 100503 151126 100555
rect 151178 100543 151184 100555
rect 204496 100543 204502 100555
rect 151178 100515 204502 100543
rect 151178 100503 151184 100515
rect 204496 100503 204502 100515
rect 204554 100503 204560 100555
rect 191440 100429 191446 100481
rect 191498 100469 191504 100481
rect 204784 100469 204790 100481
rect 191498 100441 204790 100469
rect 191498 100429 191504 100441
rect 204784 100429 204790 100441
rect 204842 100429 204848 100481
rect 143920 99985 143926 100037
rect 143978 100025 143984 100037
rect 144304 100025 144310 100037
rect 143978 99997 144310 100025
rect 143978 99985 143984 99997
rect 144304 99985 144310 99997
rect 144362 99985 144368 100037
rect 640720 99319 640726 99371
rect 640778 99359 640784 99371
rect 668176 99359 668182 99371
rect 640778 99331 668182 99359
rect 640778 99319 640784 99331
rect 668176 99319 668182 99331
rect 668234 99319 668240 99371
rect 144016 98061 144022 98113
rect 144074 98101 144080 98113
rect 180112 98101 180118 98113
rect 144074 98073 180118 98101
rect 144074 98061 144080 98073
rect 180112 98061 180118 98073
rect 180170 98061 180176 98113
rect 144112 97987 144118 98039
rect 144170 98027 144176 98039
rect 182992 98027 182998 98039
rect 144170 97999 182998 98027
rect 144170 97987 144176 97999
rect 182992 97987 182998 97999
rect 183050 97987 183056 98039
rect 144304 97913 144310 97965
rect 144362 97953 144368 97965
rect 208144 97953 208150 97965
rect 144362 97925 208150 97953
rect 144362 97913 144368 97925
rect 208144 97913 208150 97925
rect 208202 97913 208208 97965
rect 154000 97839 154006 97891
rect 154058 97879 154064 97891
rect 206512 97879 206518 97891
rect 154058 97851 206518 97879
rect 154058 97839 154064 97851
rect 206512 97839 206518 97851
rect 206570 97839 206576 97891
rect 156880 97765 156886 97817
rect 156938 97805 156944 97817
rect 204496 97805 204502 97817
rect 156938 97777 204502 97805
rect 156938 97765 156944 97777
rect 204496 97765 204502 97777
rect 204554 97765 204560 97817
rect 174256 97691 174262 97743
rect 174314 97731 174320 97743
rect 205264 97731 205270 97743
rect 174314 97703 205270 97731
rect 174314 97691 174320 97703
rect 205264 97691 205270 97703
rect 205322 97691 205328 97743
rect 177136 97617 177142 97669
rect 177194 97657 177200 97669
rect 206128 97657 206134 97669
rect 177194 97629 206134 97657
rect 177194 97617 177200 97629
rect 206128 97617 206134 97629
rect 206186 97617 206192 97669
rect 182800 97543 182806 97595
rect 182858 97583 182864 97595
rect 204496 97583 204502 97595
rect 182858 97555 204502 97583
rect 182858 97543 182864 97555
rect 204496 97543 204502 97555
rect 204554 97543 204560 97595
rect 144016 95101 144022 95153
rect 144074 95141 144080 95153
rect 174448 95141 174454 95153
rect 144074 95113 174454 95141
rect 144074 95101 144080 95113
rect 174448 95101 174454 95113
rect 174506 95101 174512 95153
rect 144112 95027 144118 95079
rect 144170 95067 144176 95079
rect 177328 95067 177334 95079
rect 144170 95039 177334 95067
rect 144170 95027 144176 95039
rect 177328 95027 177334 95039
rect 177386 95027 177392 95079
rect 146512 94953 146518 95005
rect 146570 94993 146576 95005
rect 206320 94993 206326 95005
rect 146570 94965 206326 94993
rect 146570 94953 146576 94965
rect 206320 94953 206326 94965
rect 206378 94953 206384 95005
rect 144592 94879 144598 94931
rect 144650 94919 144656 94931
rect 206896 94919 206902 94931
rect 144650 94891 206902 94919
rect 144650 94879 144656 94891
rect 206896 94879 206902 94891
rect 206954 94879 206960 94931
rect 151216 94805 151222 94857
rect 151274 94845 151280 94857
rect 204592 94845 204598 94857
rect 151274 94817 204598 94845
rect 151274 94805 151280 94817
rect 204592 94805 204598 94817
rect 204650 94805 204656 94857
rect 165616 94731 165622 94783
rect 165674 94771 165680 94783
rect 205840 94771 205846 94783
rect 165674 94743 205846 94771
rect 165674 94731 165680 94743
rect 205840 94731 205846 94743
rect 205898 94731 205904 94783
rect 168496 94657 168502 94709
rect 168554 94697 168560 94709
rect 205744 94697 205750 94709
rect 168554 94669 205750 94697
rect 168554 94657 168560 94669
rect 205744 94657 205750 94669
rect 205802 94657 205808 94709
rect 171376 94583 171382 94635
rect 171434 94623 171440 94635
rect 204496 94623 204502 94635
rect 171434 94595 204502 94623
rect 171434 94583 171440 94595
rect 204496 94583 204502 94595
rect 204554 94583 204560 94635
rect 647344 92733 647350 92785
rect 647402 92773 647408 92785
rect 660688 92773 660694 92785
rect 647402 92745 660694 92773
rect 647402 92733 647408 92745
rect 660688 92733 660694 92745
rect 660746 92733 660752 92785
rect 646672 92659 646678 92711
rect 646730 92699 646736 92711
rect 659824 92699 659830 92711
rect 646730 92671 659830 92699
rect 646730 92659 646736 92671
rect 659824 92659 659830 92671
rect 659882 92659 659888 92711
rect 647536 92585 647542 92637
rect 647594 92625 647600 92637
rect 661744 92625 661750 92637
rect 647594 92597 661750 92625
rect 647594 92585 647600 92597
rect 661744 92585 661750 92597
rect 661802 92585 661808 92637
rect 647248 92437 647254 92489
rect 647306 92477 647312 92489
rect 659728 92477 659734 92489
rect 647306 92449 659734 92477
rect 647306 92437 647312 92449
rect 659728 92437 659734 92449
rect 659786 92437 659792 92489
rect 647824 92363 647830 92415
rect 647882 92403 647888 92415
rect 663088 92403 663094 92415
rect 647882 92375 663094 92403
rect 647882 92363 647888 92375
rect 663088 92363 663094 92375
rect 663146 92363 663152 92415
rect 647728 92289 647734 92341
rect 647786 92329 647792 92341
rect 662512 92329 662518 92341
rect 647786 92301 662518 92329
rect 647786 92289 647792 92301
rect 662512 92289 662518 92301
rect 662570 92289 662576 92341
rect 144112 92215 144118 92267
rect 144170 92255 144176 92267
rect 154000 92255 154006 92267
rect 144170 92227 154006 92255
rect 144170 92215 144176 92227
rect 154000 92215 154006 92227
rect 154058 92215 154064 92267
rect 646192 92215 646198 92267
rect 646250 92255 646256 92267
rect 661168 92255 661174 92267
rect 646250 92227 661174 92255
rect 646250 92215 646256 92227
rect 661168 92215 661174 92227
rect 661226 92215 661232 92267
rect 144016 92141 144022 92193
rect 144074 92181 144080 92193
rect 171568 92181 171574 92193
rect 144074 92153 171574 92181
rect 144074 92141 144080 92153
rect 171568 92141 171574 92153
rect 171626 92141 171632 92193
rect 646576 92141 646582 92193
rect 646634 92181 646640 92193
rect 658864 92181 658870 92193
rect 646634 92153 658870 92181
rect 646634 92141 646640 92153
rect 658864 92141 658870 92153
rect 658922 92141 658928 92193
rect 203056 92067 203062 92119
rect 203114 92107 203120 92119
rect 204592 92107 204598 92119
rect 203114 92079 204598 92107
rect 203114 92067 203120 92079
rect 204592 92067 204598 92079
rect 204650 92067 204656 92119
rect 200176 91993 200182 92045
rect 200234 92033 200240 92045
rect 204496 92033 204502 92045
rect 200234 92005 204502 92033
rect 200234 91993 200240 92005
rect 204496 91993 204502 92005
rect 204554 91993 204560 92045
rect 197296 91919 197302 91971
rect 197354 91959 197360 91971
rect 204688 91959 204694 91971
rect 197354 91931 204694 91959
rect 197354 91919 197360 91931
rect 204688 91919 204694 91931
rect 204746 91919 204752 91971
rect 194416 91845 194422 91897
rect 194474 91885 194480 91897
rect 204592 91885 204598 91897
rect 194474 91857 204598 91885
rect 194474 91845 194480 91857
rect 204592 91845 204598 91857
rect 204650 91845 204656 91897
rect 188656 91771 188662 91823
rect 188714 91811 188720 91823
rect 204784 91811 204790 91823
rect 188714 91783 204790 91811
rect 188714 91771 188720 91783
rect 204784 91771 204790 91783
rect 204842 91771 204848 91823
rect 144016 89403 144022 89455
rect 144074 89443 144080 89455
rect 151216 89443 151222 89455
rect 144074 89415 151222 89443
rect 144074 89403 144080 89415
rect 151216 89403 151222 89415
rect 151274 89403 151280 89455
rect 144304 89329 144310 89381
rect 144362 89369 144368 89381
rect 165616 89369 165622 89381
rect 144362 89341 165622 89369
rect 144362 89329 144368 89341
rect 165616 89329 165622 89341
rect 165674 89329 165680 89381
rect 204976 89329 204982 89381
rect 205034 89329 205040 89381
rect 144112 89255 144118 89307
rect 144170 89295 144176 89307
rect 168496 89295 168502 89307
rect 144170 89267 168502 89295
rect 144170 89255 144176 89267
rect 168496 89255 168502 89267
rect 168554 89255 168560 89307
rect 204994 89295 205022 89329
rect 205072 89295 205078 89307
rect 204994 89267 205078 89295
rect 205072 89255 205078 89267
rect 205130 89255 205136 89307
rect 156976 89181 156982 89233
rect 157034 89221 157040 89233
rect 204688 89221 204694 89233
rect 157034 89193 204694 89221
rect 157034 89181 157040 89193
rect 204688 89181 204694 89193
rect 204746 89181 204752 89233
rect 206992 89181 206998 89233
rect 207050 89221 207056 89233
rect 207184 89221 207190 89233
rect 207050 89193 207190 89221
rect 207050 89181 207056 89193
rect 207184 89181 207190 89193
rect 207242 89181 207248 89233
rect 159856 89107 159862 89159
rect 159914 89147 159920 89159
rect 205264 89147 205270 89159
rect 159914 89119 205270 89147
rect 159914 89107 159920 89119
rect 205264 89107 205270 89119
rect 205322 89107 205328 89159
rect 162736 89033 162742 89085
rect 162794 89073 162800 89085
rect 204592 89073 204598 89085
rect 162794 89045 204598 89073
rect 162794 89033 162800 89045
rect 204592 89033 204598 89045
rect 204650 89033 204656 89085
rect 185776 88959 185782 89011
rect 185834 88999 185840 89011
rect 204496 88999 204502 89011
rect 185834 88971 204502 88999
rect 185834 88959 185840 88971
rect 204496 88959 204502 88971
rect 204554 88959 204560 89011
rect 191536 88885 191542 88937
rect 191594 88925 191600 88937
rect 204784 88925 204790 88937
rect 191594 88897 204790 88925
rect 191594 88885 191600 88897
rect 204784 88885 204790 88897
rect 204842 88885 204848 88937
rect 646864 87997 646870 88049
rect 646922 88037 646928 88049
rect 650896 88037 650902 88049
rect 646922 88009 650902 88037
rect 646922 87997 646928 88009
rect 650896 87997 650902 88009
rect 650954 87997 650960 88049
rect 658000 87297 658006 87309
rect 657058 87269 658006 87297
rect 657058 87161 657086 87269
rect 658000 87257 658006 87269
rect 658058 87257 658064 87309
rect 657040 87109 657046 87161
rect 657098 87109 657104 87161
rect 647920 87035 647926 87087
rect 647978 87075 647984 87087
rect 663280 87075 663286 87087
rect 647978 87047 663286 87075
rect 647978 87035 647984 87047
rect 663280 87035 663286 87047
rect 663338 87035 663344 87087
rect 144496 86443 144502 86495
rect 144554 86443 144560 86495
rect 647920 86443 647926 86495
rect 647978 86483 647984 86495
rect 651088 86483 651094 86495
rect 647978 86455 651094 86483
rect 647978 86443 647984 86455
rect 651088 86443 651094 86455
rect 651146 86443 651152 86495
rect 144514 86347 144542 86443
rect 154096 86369 154102 86421
rect 154154 86409 154160 86421
rect 204688 86409 204694 86421
rect 154154 86381 204694 86409
rect 154154 86369 154160 86381
rect 204688 86369 204694 86381
rect 204746 86369 204752 86421
rect 144496 86295 144502 86347
rect 144554 86295 144560 86347
rect 174352 86295 174358 86347
rect 174410 86335 174416 86347
rect 206608 86335 206614 86347
rect 174410 86307 206614 86335
rect 174410 86295 174416 86307
rect 206608 86295 206614 86307
rect 206666 86295 206672 86347
rect 177232 86221 177238 86273
rect 177290 86261 177296 86273
rect 204592 86261 204598 86273
rect 177290 86233 204598 86261
rect 177290 86221 177296 86233
rect 204592 86221 204598 86233
rect 204650 86221 204656 86273
rect 180016 86147 180022 86199
rect 180074 86187 180080 86199
rect 205552 86187 205558 86199
rect 180074 86159 205558 86187
rect 180074 86147 180080 86159
rect 205552 86147 205558 86159
rect 205610 86147 205616 86199
rect 182896 86073 182902 86125
rect 182954 86113 182960 86125
rect 204496 86113 204502 86125
rect 182954 86085 204502 86113
rect 182954 86073 182960 86085
rect 204496 86073 204502 86085
rect 204554 86073 204560 86125
rect 646864 85111 646870 85163
rect 646922 85151 646928 85163
rect 650992 85151 650998 85163
rect 646922 85123 650998 85151
rect 646922 85111 646928 85123
rect 650992 85111 650998 85123
rect 651050 85111 651056 85163
rect 146704 84963 146710 85015
rect 146762 85003 146768 85015
rect 204496 85003 204502 85015
rect 146762 84975 204502 85003
rect 146762 84963 146768 84975
rect 204496 84963 204502 84975
rect 204554 84963 204560 85015
rect 151408 83483 151414 83535
rect 151466 83523 151472 83535
rect 206224 83523 206230 83535
rect 151466 83495 206230 83523
rect 151466 83483 151472 83495
rect 206224 83483 206230 83495
rect 206282 83483 206288 83535
rect 165712 83409 165718 83461
rect 165770 83449 165776 83461
rect 206704 83449 206710 83461
rect 165770 83421 206710 83449
rect 165770 83409 165776 83421
rect 206704 83409 206710 83421
rect 206762 83409 206768 83461
rect 647920 83409 647926 83461
rect 647978 83449 647984 83461
rect 657040 83449 657046 83461
rect 647978 83421 657046 83449
rect 647978 83409 647984 83421
rect 657040 83409 657046 83421
rect 657098 83409 657104 83461
rect 168592 83335 168598 83387
rect 168650 83375 168656 83387
rect 205744 83375 205750 83387
rect 168650 83347 205750 83375
rect 168650 83335 168656 83347
rect 205744 83335 205750 83347
rect 205802 83335 205808 83387
rect 171472 83261 171478 83313
rect 171530 83301 171536 83313
rect 204496 83301 204502 83313
rect 171530 83273 204502 83301
rect 171530 83261 171536 83273
rect 204496 83261 204502 83273
rect 204554 83261 204560 83313
rect 146704 82077 146710 82129
rect 146762 82117 146768 82129
rect 204496 82117 204502 82129
rect 146762 82089 204502 82117
rect 146762 82077 146768 82089
rect 204496 82077 204502 82089
rect 204554 82077 204560 82129
rect 647920 81855 647926 81907
rect 647978 81895 647984 81907
rect 663280 81895 663286 81907
rect 647978 81867 663286 81895
rect 647978 81855 647984 81867
rect 663280 81855 663286 81867
rect 663338 81855 663344 81907
rect 645904 81781 645910 81833
rect 645962 81821 645968 81833
rect 663376 81821 663382 81833
rect 645962 81793 663382 81821
rect 645962 81781 645968 81793
rect 663376 81781 663382 81793
rect 663434 81781 663440 81833
rect 647632 81633 647638 81685
rect 647690 81673 647696 81685
rect 661072 81673 661078 81685
rect 647690 81645 661078 81673
rect 647690 81633 647696 81645
rect 661072 81633 661078 81645
rect 661130 81633 661136 81685
rect 647920 81263 647926 81315
rect 647978 81303 647984 81315
rect 657520 81303 657526 81315
rect 647978 81275 657526 81303
rect 647978 81263 647984 81275
rect 657520 81263 657526 81275
rect 657578 81263 657584 81315
rect 143920 80671 143926 80723
rect 143978 80711 143984 80723
rect 144688 80711 144694 80723
rect 143978 80683 144694 80711
rect 143978 80671 143984 80683
rect 144688 80671 144694 80683
rect 144746 80671 144752 80723
rect 659440 80671 659446 80723
rect 659498 80711 659504 80723
rect 659536 80711 659542 80723
rect 659498 80683 659542 80711
rect 659498 80671 659504 80683
rect 659536 80671 659542 80683
rect 659594 80671 659600 80723
rect 203152 80597 203158 80649
rect 203210 80637 203216 80649
rect 205264 80637 205270 80649
rect 203210 80609 205270 80637
rect 203210 80597 203216 80609
rect 205264 80597 205270 80609
rect 205322 80597 205328 80649
rect 200272 80523 200278 80575
rect 200330 80563 200336 80575
rect 204496 80563 204502 80575
rect 200330 80535 204502 80563
rect 200330 80523 200336 80535
rect 204496 80523 204502 80535
rect 204554 80523 204560 80575
rect 197392 80449 197398 80501
rect 197450 80489 197456 80501
rect 204592 80489 204598 80501
rect 197450 80461 204598 80489
rect 197450 80449 197456 80461
rect 204592 80449 204598 80461
rect 204650 80449 204656 80501
rect 194512 80375 194518 80427
rect 194570 80415 194576 80427
rect 204688 80415 204694 80427
rect 194570 80387 204694 80415
rect 194570 80375 194576 80387
rect 204688 80375 204694 80387
rect 204746 80375 204752 80427
rect 188752 80301 188758 80353
rect 188810 80341 188816 80353
rect 210160 80341 210166 80353
rect 188810 80313 210166 80341
rect 188810 80301 188816 80313
rect 210160 80301 210166 80313
rect 210218 80301 210224 80353
rect 647920 80153 647926 80205
rect 647978 80193 647984 80205
rect 656944 80193 656950 80205
rect 647978 80165 656950 80193
rect 647978 80153 647984 80165
rect 656944 80153 656950 80165
rect 657002 80153 657008 80205
rect 645424 79635 645430 79687
rect 645482 79675 645488 79687
rect 651184 79675 651190 79687
rect 645482 79647 651190 79675
rect 645482 79635 645488 79647
rect 651184 79635 651190 79647
rect 651242 79635 651248 79687
rect 647728 79265 647734 79317
rect 647786 79305 647792 79317
rect 658864 79305 658870 79317
rect 647786 79277 658870 79305
rect 647786 79265 647792 79277
rect 658864 79265 658870 79277
rect 658922 79265 658928 79317
rect 647824 78821 647830 78873
rect 647882 78861 647888 78873
rect 660688 78861 660694 78873
rect 647882 78833 660694 78861
rect 647882 78821 647888 78833
rect 660688 78821 660694 78833
rect 660746 78821 660752 78873
rect 647920 78303 647926 78355
rect 647978 78343 647984 78355
rect 662512 78343 662518 78355
rect 647978 78315 662518 78343
rect 647978 78303 647984 78315
rect 662512 78303 662518 78315
rect 662570 78303 662576 78355
rect 144304 77859 144310 77911
rect 144362 77899 144368 77911
rect 151120 77899 151126 77911
rect 144362 77871 151126 77899
rect 144362 77859 144368 77871
rect 151120 77859 151126 77871
rect 151178 77859 151184 77911
rect 146704 77785 146710 77837
rect 146762 77825 146768 77837
rect 146762 77797 190046 77825
rect 146762 77785 146768 77797
rect 146608 77711 146614 77763
rect 146666 77711 146672 77763
rect 157072 77711 157078 77763
rect 157130 77751 157136 77763
rect 189904 77751 189910 77763
rect 157130 77723 189910 77751
rect 157130 77711 157136 77723
rect 189904 77711 189910 77723
rect 189962 77711 189968 77763
rect 190018 77751 190046 77797
rect 204592 77751 204598 77763
rect 190018 77723 204598 77751
rect 204592 77711 204598 77723
rect 204650 77711 204656 77763
rect 647440 77711 647446 77763
rect 647498 77751 647504 77763
rect 659440 77751 659446 77763
rect 647498 77723 659446 77751
rect 647498 77711 647504 77723
rect 659440 77711 659446 77723
rect 659498 77711 659504 77763
rect 146626 77467 146654 77711
rect 159952 77637 159958 77689
rect 160010 77677 160016 77689
rect 206512 77677 206518 77689
rect 160010 77649 206518 77677
rect 160010 77637 160016 77649
rect 206512 77637 206518 77649
rect 206570 77637 206576 77689
rect 647920 77637 647926 77689
rect 647978 77677 647984 77689
rect 650992 77677 650998 77689
rect 647978 77649 650998 77677
rect 647978 77637 647984 77649
rect 650992 77637 650998 77649
rect 651050 77637 651056 77689
rect 162832 77563 162838 77615
rect 162890 77603 162896 77615
rect 204496 77603 204502 77615
rect 162890 77575 204502 77603
rect 162890 77563 162896 77575
rect 204496 77563 204502 77575
rect 204554 77563 204560 77615
rect 185872 77489 185878 77541
rect 185930 77529 185936 77541
rect 205936 77529 205942 77541
rect 185930 77501 205942 77529
rect 185930 77489 185936 77501
rect 205936 77489 205942 77501
rect 205994 77489 206000 77541
rect 146608 77415 146614 77467
rect 146666 77415 146672 77467
rect 189904 77415 189910 77467
rect 189962 77455 189968 77467
rect 204688 77455 204694 77467
rect 189962 77427 204694 77455
rect 189962 77415 189968 77427
rect 204688 77415 204694 77427
rect 204746 77415 204752 77467
rect 191632 77341 191638 77393
rect 191690 77381 191696 77393
rect 204784 77381 204790 77393
rect 191690 77353 204790 77381
rect 191690 77341 191696 77353
rect 204784 77341 204790 77353
rect 204842 77341 204848 77393
rect 647920 77267 647926 77319
rect 647978 77307 647984 77319
rect 662896 77307 662902 77319
rect 647978 77279 662902 77307
rect 647978 77267 647984 77279
rect 662896 77267 662902 77279
rect 662954 77267 662960 77319
rect 646480 76897 646486 76949
rect 646538 76937 646544 76949
rect 658288 76937 658294 76949
rect 646538 76909 658294 76937
rect 646538 76897 646544 76909
rect 658288 76897 658294 76909
rect 658346 76897 658352 76949
rect 646480 76749 646486 76801
rect 646538 76789 646544 76801
rect 650896 76789 650902 76801
rect 646538 76761 650902 76789
rect 646538 76749 646544 76761
rect 650896 76749 650902 76761
rect 650954 76749 650960 76801
rect 646096 75787 646102 75839
rect 646154 75827 646160 75839
rect 661744 75827 661750 75839
rect 646154 75799 661750 75827
rect 646154 75787 646160 75799
rect 661744 75787 661750 75799
rect 661802 75787 661808 75839
rect 646480 75417 646486 75469
rect 646538 75457 646544 75469
rect 656848 75457 656854 75469
rect 646538 75429 656854 75457
rect 646538 75417 646544 75429
rect 656848 75417 656854 75429
rect 656906 75417 656912 75469
rect 146512 75047 146518 75099
rect 146570 75087 146576 75099
rect 160144 75087 160150 75099
rect 146570 75059 160150 75087
rect 146570 75047 146576 75059
rect 160144 75047 160150 75059
rect 160202 75047 160208 75099
rect 144016 74973 144022 75025
rect 144074 75013 144080 75025
rect 156976 75013 156982 75025
rect 144074 74985 156982 75013
rect 144074 74973 144080 74985
rect 156976 74973 156982 74985
rect 157034 74973 157040 75025
rect 144304 74899 144310 74951
rect 144362 74939 144368 74951
rect 161488 74939 161494 74951
rect 144362 74911 161494 74939
rect 144362 74899 144368 74911
rect 161488 74899 161494 74911
rect 161546 74899 161552 74951
rect 154000 74825 154006 74877
rect 154058 74865 154064 74877
rect 204688 74865 204694 74877
rect 154058 74837 204694 74865
rect 154058 74825 154064 74837
rect 204688 74825 204694 74837
rect 204746 74825 204752 74877
rect 174448 74751 174454 74803
rect 174506 74791 174512 74803
rect 206800 74791 206806 74803
rect 174506 74763 206806 74791
rect 174506 74751 174512 74763
rect 206800 74751 206806 74763
rect 206858 74751 206864 74803
rect 177328 74677 177334 74729
rect 177386 74717 177392 74729
rect 204592 74717 204598 74729
rect 177386 74689 204598 74717
rect 177386 74677 177392 74689
rect 204592 74677 204598 74689
rect 204650 74677 204656 74729
rect 180112 74603 180118 74655
rect 180170 74643 180176 74655
rect 205744 74643 205750 74655
rect 180170 74615 205750 74643
rect 180170 74603 180176 74615
rect 205744 74603 205750 74615
rect 205802 74603 205808 74655
rect 182992 74529 182998 74581
rect 183050 74569 183056 74581
rect 204496 74569 204502 74581
rect 183050 74541 204502 74569
rect 183050 74529 183056 74541
rect 204496 74529 204502 74541
rect 204554 74529 204560 74581
rect 144304 74159 144310 74211
rect 144362 74199 144368 74211
rect 145456 74199 145462 74211
rect 144362 74171 145462 74199
rect 144362 74159 144368 74171
rect 145456 74159 145462 74171
rect 145514 74159 145520 74211
rect 144112 74085 144118 74137
rect 144170 74125 144176 74137
rect 148336 74125 148342 74137
rect 144170 74097 148342 74125
rect 144170 74085 144176 74097
rect 148336 74085 148342 74097
rect 148394 74085 148400 74137
rect 145456 74011 145462 74063
rect 145514 74051 145520 74063
rect 146032 74051 146038 74063
rect 145514 74023 146038 74051
rect 145514 74011 145520 74023
rect 146032 74011 146038 74023
rect 146090 74011 146096 74063
rect 647248 72531 647254 72583
rect 647306 72571 647312 72583
rect 663184 72571 663190 72583
rect 647306 72543 663190 72571
rect 647306 72531 647312 72543
rect 663184 72531 663190 72543
rect 663242 72531 663248 72583
rect 646864 72457 646870 72509
rect 646922 72497 646928 72509
rect 660112 72497 660118 72509
rect 646922 72469 660118 72497
rect 646922 72457 646928 72469
rect 660112 72457 660118 72469
rect 660170 72457 660176 72509
rect 646096 72235 646102 72287
rect 646154 72275 646160 72287
rect 663376 72275 663382 72287
rect 646154 72247 663382 72275
rect 646154 72235 646160 72247
rect 663376 72235 663382 72247
rect 663434 72235 663440 72287
rect 146032 72013 146038 72065
rect 146090 72053 146096 72065
rect 154672 72053 154678 72065
rect 146090 72025 154678 72053
rect 146090 72013 146096 72025
rect 154672 72013 154678 72025
rect 154730 72013 154736 72065
rect 151216 71939 151222 71991
rect 151274 71979 151280 71991
rect 206800 71979 206806 71991
rect 151274 71951 206806 71979
rect 151274 71939 151280 71951
rect 206800 71939 206806 71951
rect 206858 71939 206864 71991
rect 161488 71865 161494 71917
rect 161546 71905 161552 71917
rect 204976 71905 204982 71917
rect 161546 71877 204982 71905
rect 161546 71865 161552 71877
rect 204976 71865 204982 71877
rect 205034 71865 205040 71917
rect 165616 71791 165622 71843
rect 165674 71831 165680 71843
rect 205456 71831 205462 71843
rect 165674 71803 205462 71831
rect 165674 71791 165680 71803
rect 205456 71791 205462 71803
rect 205514 71791 205520 71843
rect 168496 71717 168502 71769
rect 168554 71757 168560 71769
rect 204592 71757 204598 71769
rect 168554 71729 204598 71757
rect 168554 71717 168560 71729
rect 204592 71717 204598 71729
rect 204650 71717 204656 71769
rect 171568 71643 171574 71695
rect 171626 71683 171632 71695
rect 204496 71683 204502 71695
rect 171626 71655 204502 71683
rect 171626 71643 171632 71655
rect 204496 71643 204502 71655
rect 204554 71643 204560 71695
rect 144016 70237 144022 70289
rect 144074 70277 144080 70289
rect 149776 70277 149782 70289
rect 144074 70249 149782 70277
rect 144074 70237 144080 70249
rect 149776 70237 149782 70249
rect 149834 70237 149840 70289
rect 146032 69201 146038 69253
rect 146090 69241 146096 69253
rect 146320 69241 146326 69253
rect 146090 69213 146326 69241
rect 146090 69201 146096 69213
rect 146320 69201 146326 69213
rect 146378 69201 146384 69253
rect 144016 69127 144022 69179
rect 144074 69167 144080 69179
rect 144074 69139 146942 69167
rect 144074 69127 144080 69139
rect 146914 69093 146942 69139
rect 206992 69127 206998 69179
rect 207050 69167 207056 69179
rect 207280 69167 207286 69179
rect 207050 69139 207286 69167
rect 207050 69127 207056 69139
rect 207280 69127 207286 69139
rect 207338 69127 207344 69179
rect 206512 69093 206518 69105
rect 146914 69065 206518 69093
rect 206512 69053 206518 69065
rect 206570 69053 206576 69105
rect 149776 68979 149782 69031
rect 149834 69019 149840 69031
rect 204112 69019 204118 69031
rect 149834 68991 204118 69019
rect 149834 68979 149840 68991
rect 204112 68979 204118 68991
rect 204170 68979 204176 69031
rect 205168 68979 205174 69031
rect 205226 69019 205232 69031
rect 207472 69019 207478 69031
rect 205226 68991 207478 69019
rect 205226 68979 205232 68991
rect 207472 68979 207478 68991
rect 207530 68979 207536 69031
rect 154672 68905 154678 68957
rect 154730 68945 154736 68957
rect 204592 68945 204598 68957
rect 154730 68917 204598 68945
rect 154730 68905 154736 68917
rect 204592 68905 204598 68917
rect 204650 68905 204656 68957
rect 156976 68831 156982 68883
rect 157034 68871 157040 68883
rect 206416 68871 206422 68883
rect 157034 68843 206422 68871
rect 157034 68831 157040 68843
rect 206416 68831 206422 68843
rect 206474 68831 206480 68883
rect 160144 68757 160150 68809
rect 160202 68797 160208 68809
rect 204496 68797 204502 68809
rect 160202 68769 204502 68797
rect 160202 68757 160208 68769
rect 204496 68757 204502 68769
rect 204554 68757 204560 68809
rect 144112 67203 144118 67255
rect 144170 67243 144176 67255
rect 152656 67243 152662 67255
rect 144170 67215 152662 67243
rect 144170 67203 144176 67215
rect 152656 67203 152662 67215
rect 152714 67203 152720 67255
rect 146320 66389 146326 66441
rect 146378 66429 146384 66441
rect 158320 66429 158326 66441
rect 146378 66401 158326 66429
rect 146378 66389 146384 66401
rect 158320 66389 158326 66401
rect 158378 66389 158384 66441
rect 146800 66241 146806 66293
rect 146858 66281 146864 66293
rect 146858 66253 149822 66281
rect 146858 66241 146864 66253
rect 144016 66167 144022 66219
rect 144074 66207 144080 66219
rect 144688 66207 144694 66219
rect 144074 66179 144694 66207
rect 144074 66167 144080 66179
rect 144688 66167 144694 66179
rect 144746 66167 144752 66219
rect 149794 66207 149822 66253
rect 205456 66207 205462 66219
rect 149794 66179 205462 66207
rect 205456 66167 205462 66179
rect 205514 66167 205520 66219
rect 152656 66093 152662 66145
rect 152714 66133 152720 66145
rect 206320 66133 206326 66145
rect 152714 66105 206326 66133
rect 152714 66093 152720 66105
rect 206320 66093 206326 66105
rect 206378 66093 206384 66145
rect 158320 66019 158326 66071
rect 158378 66059 158384 66071
rect 204496 66059 204502 66071
rect 158378 66031 204502 66059
rect 158378 66019 158384 66031
rect 204496 66019 204502 66031
rect 204554 66019 204560 66071
rect 145456 65871 145462 65923
rect 145514 65911 145520 65923
rect 146320 65911 146326 65923
rect 145514 65883 146326 65911
rect 145514 65871 145520 65883
rect 146320 65871 146326 65883
rect 146378 65871 146384 65923
rect 145072 65723 145078 65775
rect 145130 65763 145136 65775
rect 145456 65763 145462 65775
rect 145130 65735 145462 65763
rect 145130 65723 145136 65735
rect 145456 65723 145462 65735
rect 145514 65723 145520 65775
rect 144112 64983 144118 65035
rect 144170 65023 144176 65035
rect 144304 65023 144310 65035
rect 144170 64995 144310 65023
rect 144170 64983 144176 64995
rect 144304 64983 144310 64995
rect 144362 64983 144368 65035
rect 144304 64835 144310 64887
rect 144362 64875 144368 64887
rect 204592 64875 204598 64887
rect 144362 64847 204598 64875
rect 144362 64835 144368 64847
rect 204592 64835 204598 64847
rect 204650 64835 204656 64887
rect 144976 64761 144982 64813
rect 145034 64801 145040 64813
rect 204496 64801 204502 64813
rect 145034 64773 204502 64801
rect 145034 64761 145040 64773
rect 204496 64761 204502 64773
rect 204554 64761 204560 64813
rect 146896 63355 146902 63407
rect 146954 63395 146960 63407
rect 204496 63395 204502 63407
rect 146954 63367 204502 63395
rect 146954 63355 146960 63367
rect 204496 63355 204502 63367
rect 204554 63355 204560 63407
rect 144016 62911 144022 62963
rect 144074 62951 144080 62963
rect 144304 62951 144310 62963
rect 144074 62923 144310 62951
rect 144074 62911 144080 62923
rect 144304 62911 144310 62923
rect 144362 62911 144368 62963
rect 144016 62467 144022 62519
rect 144074 62507 144080 62519
rect 149776 62507 149782 62519
rect 144074 62479 149782 62507
rect 144074 62467 144080 62479
rect 149776 62467 149782 62479
rect 149834 62467 149840 62519
rect 160528 60765 160534 60817
rect 160586 60805 160592 60817
rect 204592 60805 204598 60817
rect 160586 60777 204598 60805
rect 160586 60765 160592 60777
rect 204592 60765 204598 60777
rect 204650 60765 204656 60817
rect 156304 60691 156310 60743
rect 156362 60731 156368 60743
rect 204688 60731 204694 60743
rect 156362 60703 204694 60731
rect 156362 60691 156368 60703
rect 204688 60691 204694 60703
rect 204746 60691 204752 60743
rect 152656 60617 152662 60669
rect 152714 60657 152720 60669
rect 204496 60657 204502 60669
rect 152714 60629 204502 60657
rect 152714 60617 152720 60629
rect 204496 60617 204502 60629
rect 204554 60617 204560 60669
rect 151216 60543 151222 60595
rect 151274 60583 151280 60595
rect 204880 60583 204886 60595
rect 151274 60555 204886 60583
rect 151274 60543 151280 60555
rect 204880 60543 204886 60555
rect 204938 60543 204944 60595
rect 148336 60469 148342 60521
rect 148394 60509 148400 60521
rect 204784 60509 204790 60521
rect 148394 60481 204790 60509
rect 148394 60469 148400 60481
rect 204784 60469 204790 60481
rect 204842 60469 204848 60521
rect 146896 60395 146902 60447
rect 146954 60435 146960 60447
rect 206800 60435 206806 60447
rect 146954 60407 206806 60435
rect 146954 60395 146960 60407
rect 206800 60395 206806 60407
rect 206858 60395 206864 60447
rect 149776 60321 149782 60373
rect 149834 60361 149840 60373
rect 204592 60361 204598 60373
rect 149834 60333 204598 60361
rect 149834 60321 149840 60333
rect 204592 60321 204598 60333
rect 204650 60321 204656 60373
rect 207760 60321 207766 60373
rect 207818 60361 207824 60373
rect 208720 60361 208726 60373
rect 207818 60333 208726 60361
rect 207818 60321 207824 60333
rect 208720 60321 208726 60333
rect 208778 60321 208784 60373
rect 207856 60247 207862 60299
rect 207914 60287 207920 60299
rect 208816 60287 208822 60299
rect 207914 60259 208822 60287
rect 207914 60247 207920 60259
rect 208816 60247 208822 60259
rect 208874 60247 208880 60299
rect 208816 59951 208822 60003
rect 208874 59991 208880 60003
rect 209104 59991 209110 60003
rect 208874 59963 209110 59991
rect 208874 59951 208880 59963
rect 209104 59951 209110 59963
rect 209162 59951 209168 60003
rect 209488 59951 209494 60003
rect 209546 59991 209552 60003
rect 209968 59991 209974 60003
rect 209546 59963 209974 59991
rect 209546 59951 209552 59963
rect 209968 59951 209974 59963
rect 210026 59951 210032 60003
rect 144016 59581 144022 59633
rect 144074 59621 144080 59633
rect 160528 59621 160534 59633
rect 144074 59593 160534 59621
rect 144074 59581 144080 59593
rect 160528 59581 160534 59593
rect 160586 59581 160592 59633
rect 144016 58989 144022 59041
rect 144074 59029 144080 59041
rect 204496 59029 204502 59041
rect 144074 59001 204502 59029
rect 144074 58989 144080 59001
rect 204496 58989 204502 59001
rect 204554 58989 204560 59041
rect 144016 57065 144022 57117
rect 144074 57105 144080 57117
rect 156304 57105 156310 57117
rect 144074 57077 156310 57105
rect 144074 57065 144080 57077
rect 156304 57065 156310 57077
rect 156362 57065 156368 57117
rect 144016 56473 144022 56525
rect 144074 56513 144080 56525
rect 152656 56513 152662 56525
rect 144074 56485 152662 56513
rect 144074 56473 144080 56485
rect 152656 56473 152662 56485
rect 152714 56473 152720 56525
rect 209968 54845 209974 54897
rect 210026 54845 210032 54897
rect 144016 54623 144022 54675
rect 144074 54663 144080 54675
rect 151216 54663 151222 54675
rect 144074 54635 151222 54663
rect 144074 54623 144080 54635
rect 151216 54623 151222 54635
rect 151274 54623 151280 54675
rect 209986 54589 210014 54845
rect 209986 54561 210110 54589
rect 210082 54441 210110 54561
rect 210082 54413 221054 54441
rect 221026 54305 221054 54413
rect 210160 54253 210166 54305
rect 210218 54293 210224 54305
rect 218992 54293 218998 54305
rect 210218 54265 218998 54293
rect 210218 54253 210224 54265
rect 218992 54253 218998 54265
rect 219050 54253 219056 54305
rect 221008 54253 221014 54305
rect 221066 54253 221072 54305
rect 207472 54179 207478 54231
rect 207530 54219 207536 54231
rect 216304 54219 216310 54231
rect 207530 54191 216310 54219
rect 207530 54179 207536 54191
rect 216304 54179 216310 54191
rect 216362 54179 216368 54231
rect 144016 54105 144022 54157
rect 144074 54145 144080 54157
rect 148336 54145 148342 54157
rect 144074 54117 148342 54145
rect 144074 54105 144080 54117
rect 148336 54105 148342 54117
rect 148394 54105 148400 54157
rect 210064 54105 210070 54157
rect 210122 54145 210128 54157
rect 219184 54145 219190 54157
rect 210122 54117 219190 54145
rect 210122 54105 210128 54117
rect 219184 54105 219190 54117
rect 219242 54105 219248 54157
rect 209200 54031 209206 54083
rect 209258 54071 209264 54083
rect 218992 54071 218998 54083
rect 209258 54043 218998 54071
rect 209258 54031 209264 54043
rect 218992 54031 218998 54043
rect 219050 54031 219056 54083
rect 209296 53957 209302 54009
rect 209354 53997 209360 54009
rect 218800 53997 218806 54009
rect 209354 53969 218806 53997
rect 209354 53957 209360 53969
rect 218800 53957 218806 53969
rect 218858 53957 218864 54009
rect 208432 53883 208438 53935
rect 208490 53923 208496 53935
rect 219184 53923 219190 53935
rect 208490 53895 219190 53923
rect 208490 53883 208496 53895
rect 219184 53883 219190 53895
rect 219242 53883 219248 53935
rect 208048 53809 208054 53861
rect 208106 53849 208112 53861
rect 216784 53849 216790 53861
rect 208106 53821 216790 53849
rect 208106 53809 208112 53821
rect 216784 53809 216790 53821
rect 216842 53809 216848 53861
rect 212368 53735 212374 53787
rect 212426 53775 212432 53787
rect 221200 53775 221206 53787
rect 212426 53747 221206 53775
rect 212426 53735 212432 53747
rect 221200 53735 221206 53747
rect 221258 53735 221264 53787
rect 210256 53661 210262 53713
rect 210314 53701 210320 53713
rect 293776 53701 293782 53713
rect 210314 53673 293782 53701
rect 210314 53661 210320 53673
rect 293776 53661 293782 53673
rect 293834 53661 293840 53713
rect 209968 53587 209974 53639
rect 210026 53627 210032 53639
rect 330928 53627 330934 53639
rect 210026 53599 330934 53627
rect 210026 53587 210032 53599
rect 330928 53587 330934 53599
rect 330986 53587 330992 53639
rect 211552 53513 211558 53565
rect 211610 53553 211616 53565
rect 216592 53553 216598 53565
rect 211610 53525 216598 53553
rect 211610 53513 211616 53525
rect 216592 53513 216598 53525
rect 216650 53513 216656 53565
rect 219184 53513 219190 53565
rect 219242 53553 219248 53565
rect 219808 53553 219814 53565
rect 219242 53525 219814 53553
rect 219242 53513 219248 53525
rect 219808 53513 219814 53525
rect 219866 53513 219872 53565
rect 221008 53513 221014 53565
rect 221066 53553 221072 53565
rect 403120 53553 403126 53565
rect 221066 53525 403126 53553
rect 221066 53513 221072 53525
rect 403120 53513 403126 53525
rect 403178 53513 403184 53565
rect 210352 53439 210358 53491
rect 210410 53479 210416 53491
rect 217792 53479 217798 53491
rect 210410 53451 217798 53479
rect 210410 53439 210416 53451
rect 217792 53439 217798 53451
rect 217850 53439 217856 53491
rect 218992 53439 218998 53491
rect 219050 53479 219056 53491
rect 452176 53479 452182 53491
rect 219050 53451 452182 53479
rect 219050 53439 219056 53451
rect 452176 53439 452182 53451
rect 452234 53439 452240 53491
rect 209584 53365 209590 53417
rect 209642 53405 209648 53417
rect 217456 53405 217462 53417
rect 209642 53377 217462 53405
rect 209642 53365 209648 53377
rect 217456 53365 217462 53377
rect 217514 53365 217520 53417
rect 218800 53365 218806 53417
rect 218858 53405 218864 53417
rect 466480 53405 466486 53417
rect 218858 53377 466486 53405
rect 218858 53365 218864 53377
rect 466480 53365 466486 53377
rect 466538 53365 466544 53417
rect 209392 53291 209398 53343
rect 209450 53331 209456 53343
rect 219664 53331 219670 53343
rect 209450 53303 219670 53331
rect 209450 53291 209456 53303
rect 219664 53291 219670 53303
rect 219722 53291 219728 53343
rect 219856 53291 219862 53343
rect 219914 53331 219920 53343
rect 517840 53331 517846 53343
rect 219914 53303 517846 53331
rect 219914 53291 219920 53303
rect 517840 53291 517846 53303
rect 517898 53291 517904 53343
rect 207184 53217 207190 53269
rect 207242 53257 207248 53269
rect 215536 53257 215542 53269
rect 207242 53229 215542 53257
rect 207242 53217 207248 53229
rect 215536 53217 215542 53229
rect 215594 53217 215600 53269
rect 308080 53257 308086 53269
rect 241954 53229 247742 53257
rect 209776 53143 209782 53195
rect 209834 53183 209840 53195
rect 213328 53183 213334 53195
rect 209834 53155 213334 53183
rect 209834 53143 209840 53155
rect 213328 53143 213334 53155
rect 213386 53143 213392 53195
rect 208144 53069 208150 53121
rect 208202 53109 208208 53121
rect 215728 53109 215734 53121
rect 208202 53081 215734 53109
rect 208202 53069 208208 53081
rect 215728 53069 215734 53081
rect 215786 53069 215792 53121
rect 216016 53069 216022 53121
rect 216074 53109 216080 53121
rect 241954 53109 241982 53229
rect 247714 53183 247742 53229
rect 267778 53229 287966 53257
rect 267778 53183 267806 53229
rect 247714 53155 267806 53183
rect 287938 53183 287966 53229
rect 291202 53229 308086 53257
rect 291202 53183 291230 53229
rect 308080 53217 308086 53229
rect 308138 53217 308144 53269
rect 348400 53257 348406 53269
rect 322498 53229 328286 53257
rect 287938 53155 291230 53183
rect 308176 53143 308182 53195
rect 308234 53183 308240 53195
rect 322498 53183 322526 53229
rect 308234 53155 322526 53183
rect 328258 53183 328286 53229
rect 331810 53229 348406 53257
rect 331810 53183 331838 53229
rect 348400 53217 348406 53229
rect 348458 53217 348464 53269
rect 420496 53257 420502 53269
rect 362818 53229 368606 53257
rect 328258 53155 331838 53183
rect 308234 53143 308240 53155
rect 348496 53143 348502 53195
rect 348554 53183 348560 53195
rect 362818 53183 362846 53229
rect 348554 53155 362846 53183
rect 348554 53143 348560 53155
rect 216074 53081 241982 53109
rect 216074 53069 216080 53081
rect 207952 52995 207958 53047
rect 208010 53035 208016 53047
rect 218128 53035 218134 53047
rect 208010 53007 218134 53035
rect 208010 52995 208016 53007
rect 218128 52995 218134 53007
rect 218186 52995 218192 53047
rect 368578 53035 368606 53229
rect 412370 53229 420502 53257
rect 412370 53109 412398 53229
rect 420496 53217 420502 53229
rect 420554 53217 420560 53269
rect 443536 53217 443542 53269
rect 443594 53257 443600 53269
rect 443594 53229 457982 53257
rect 443594 53217 443600 53229
rect 457954 53183 457982 53229
rect 463696 53217 463702 53269
rect 463754 53257 463760 53269
rect 483856 53257 483862 53269
rect 463754 53229 483862 53257
rect 463754 53217 463760 53229
rect 483856 53217 483862 53229
rect 483914 53217 483920 53269
rect 463600 53183 463606 53195
rect 457954 53155 463606 53183
rect 463600 53143 463606 53155
rect 463658 53143 463664 53195
rect 383074 53081 412398 53109
rect 383074 53035 383102 53081
rect 420592 53069 420598 53121
rect 420650 53109 420656 53121
rect 443440 53109 443446 53121
rect 420650 53081 443446 53109
rect 420650 53069 420656 53081
rect 443440 53069 443446 53081
rect 443498 53069 443504 53121
rect 368578 53007 383102 53035
rect 483856 52995 483862 53047
rect 483914 53035 483920 53047
rect 514000 53035 514006 53047
rect 483914 53007 514006 53035
rect 483914 52995 483920 53007
rect 514000 52995 514006 53007
rect 514058 52995 514064 53047
rect 207280 52847 207286 52899
rect 207338 52887 207344 52899
rect 219856 52887 219862 52899
rect 207338 52859 219862 52887
rect 207338 52847 207344 52859
rect 219856 52847 219862 52859
rect 219914 52847 219920 52899
rect 212176 52625 212182 52677
rect 212234 52665 212240 52677
rect 220912 52665 220918 52677
rect 212234 52637 220918 52665
rect 212234 52625 212240 52637
rect 220912 52625 220918 52637
rect 220970 52625 220976 52677
rect 151312 52551 151318 52603
rect 151370 52591 151376 52603
rect 217264 52591 217270 52603
rect 151370 52563 217270 52591
rect 151370 52551 151376 52563
rect 217264 52551 217270 52563
rect 217322 52551 217328 52603
rect 151120 52403 151126 52455
rect 151178 52443 151184 52455
rect 216112 52443 216118 52455
rect 151178 52415 216118 52443
rect 151178 52403 151184 52415
rect 216112 52403 216118 52415
rect 216170 52403 216176 52455
rect 211216 52329 211222 52381
rect 211274 52369 211280 52381
rect 227440 52369 227446 52381
rect 211274 52341 227446 52369
rect 211274 52329 211280 52341
rect 227440 52329 227446 52341
rect 227498 52329 227504 52381
rect 137488 52255 137494 52307
rect 137546 52295 137552 52307
rect 221776 52295 221782 52307
rect 137546 52267 221782 52295
rect 137546 52255 137552 52267
rect 221776 52255 221782 52267
rect 221834 52255 221840 52307
rect 227152 52221 227158 52233
rect 211618 52193 227158 52221
rect 146704 52107 146710 52159
rect 146762 52147 146768 52159
rect 161296 52147 161302 52159
rect 146762 52119 161302 52147
rect 146762 52107 146768 52119
rect 161296 52107 161302 52119
rect 161354 52107 161360 52159
rect 181360 52107 181366 52159
rect 181418 52147 181424 52159
rect 211618 52147 211646 52193
rect 227152 52181 227158 52193
rect 227210 52181 227216 52233
rect 225712 52147 225718 52159
rect 181418 52119 211646 52147
rect 212290 52119 225718 52147
rect 181418 52107 181424 52119
rect 144400 52033 144406 52085
rect 144458 52073 144464 52085
rect 212176 52073 212182 52085
rect 144458 52045 212182 52073
rect 144458 52033 144464 52045
rect 212176 52033 212182 52045
rect 212234 52033 212240 52085
rect 144592 51959 144598 52011
rect 144650 51999 144656 52011
rect 212290 51999 212318 52119
rect 225712 52107 225718 52119
rect 225770 52107 225776 52159
rect 212368 52033 212374 52085
rect 212426 52073 212432 52085
rect 213424 52073 213430 52085
rect 212426 52045 213430 52073
rect 212426 52033 212432 52045
rect 213424 52033 213430 52045
rect 213482 52033 213488 52085
rect 144650 51971 212318 51999
rect 213346 51971 213566 51999
rect 144650 51959 144656 51971
rect 146512 51885 146518 51937
rect 146570 51925 146576 51937
rect 213346 51925 213374 51971
rect 146570 51897 213374 51925
rect 213538 51925 213566 51971
rect 227536 51925 227542 51937
rect 213538 51897 227542 51925
rect 146570 51885 146576 51897
rect 227536 51885 227542 51897
rect 227594 51885 227600 51937
rect 423376 51885 423382 51937
rect 423434 51925 423440 51937
rect 432784 51925 432790 51937
rect 423434 51897 432790 51925
rect 423434 51885 423440 51897
rect 432784 51885 432790 51897
rect 432842 51885 432848 51937
rect 483856 51885 483862 51937
rect 483914 51925 483920 51937
rect 493840 51925 493846 51937
rect 483914 51897 493846 51925
rect 483914 51885 483920 51897
rect 493840 51885 493846 51897
rect 493898 51885 493904 51937
rect 544336 51885 544342 51937
rect 544394 51925 544400 51937
rect 552784 51925 552790 51937
rect 544394 51897 552790 51925
rect 544394 51885 544400 51897
rect 552784 51885 552790 51897
rect 552842 51885 552848 51937
rect 625744 51885 625750 51937
rect 625802 51925 625808 51937
rect 639664 51925 639670 51937
rect 625802 51897 639670 51925
rect 625802 51885 625808 51897
rect 639664 51885 639670 51897
rect 639722 51885 639728 51937
rect 213424 51811 213430 51863
rect 213482 51851 213488 51863
rect 645520 51851 645526 51863
rect 213482 51823 645526 51851
rect 213482 51811 213488 51823
rect 645520 51811 645526 51823
rect 645578 51811 645584 51863
rect 209680 51737 209686 51789
rect 209738 51777 209744 51789
rect 213712 51777 213718 51789
rect 209738 51749 213718 51777
rect 209738 51737 209744 51749
rect 213712 51737 213718 51749
rect 213770 51737 213776 51789
rect 216592 51737 216598 51789
rect 216650 51777 216656 51789
rect 645712 51777 645718 51789
rect 216650 51749 645718 51777
rect 216650 51737 216656 51749
rect 645712 51737 645718 51749
rect 645770 51737 645776 51789
rect 209872 51663 209878 51715
rect 209930 51703 209936 51715
rect 214096 51703 214102 51715
rect 209930 51675 214102 51703
rect 209930 51663 209936 51675
rect 214096 51663 214102 51675
rect 214154 51663 214160 51715
rect 287920 51703 287926 51715
rect 267778 51675 287926 51703
rect 221776 51589 221782 51641
rect 221834 51629 221840 51641
rect 243856 51629 243862 51641
rect 221834 51601 243862 51629
rect 221834 51589 221840 51601
rect 243856 51589 243862 51601
rect 243914 51589 243920 51641
rect 145360 51515 145366 51567
rect 145418 51555 145424 51567
rect 237616 51555 237622 51567
rect 145418 51527 237622 51555
rect 145418 51515 145424 51527
rect 237616 51515 237622 51527
rect 237674 51515 237680 51567
rect 145552 51441 145558 51493
rect 145610 51481 145616 51493
rect 236368 51481 236374 51493
rect 145610 51453 236374 51481
rect 145610 51441 145616 51453
rect 236368 51441 236374 51453
rect 236426 51441 236432 51493
rect 145936 51367 145942 51419
rect 145994 51407 146000 51419
rect 237136 51407 237142 51419
rect 145994 51379 237142 51407
rect 145994 51367 146000 51379
rect 237136 51367 237142 51379
rect 237194 51367 237200 51419
rect 267778 51407 267806 51675
rect 287920 51663 287926 51675
rect 287978 51663 287984 51715
rect 288016 51663 288022 51715
rect 288074 51703 288080 51715
rect 292048 51703 292054 51715
rect 288074 51675 292054 51703
rect 288074 51663 288080 51675
rect 292048 51663 292054 51675
rect 292106 51663 292112 51715
rect 348400 51703 348406 51715
rect 329890 51675 348406 51703
rect 302338 51601 302462 51629
rect 292048 51515 292054 51567
rect 292106 51555 292112 51567
rect 302338 51555 302366 51601
rect 302434 51567 302462 51601
rect 292106 51527 302366 51555
rect 292106 51515 292112 51527
rect 302416 51515 302422 51567
rect 302474 51515 302480 51567
rect 302512 51515 302518 51567
rect 302570 51555 302576 51567
rect 322576 51555 322582 51567
rect 302570 51527 322582 51555
rect 302570 51515 302576 51527
rect 322576 51515 322582 51527
rect 322634 51515 322640 51567
rect 252034 51379 267806 51407
rect 144304 51293 144310 51345
rect 144362 51333 144368 51345
rect 144362 51305 217502 51333
rect 144362 51293 144368 51305
rect 145648 51219 145654 51271
rect 145706 51259 145712 51271
rect 217474 51259 217502 51305
rect 227440 51293 227446 51345
rect 227498 51333 227504 51345
rect 227498 51305 247550 51333
rect 227498 51293 227504 51305
rect 233776 51259 233782 51271
rect 145706 51231 217406 51259
rect 217474 51231 233782 51259
rect 145706 51219 145712 51231
rect 145744 51145 145750 51197
rect 145802 51185 145808 51197
rect 217264 51185 217270 51197
rect 145802 51157 217270 51185
rect 145802 51145 145808 51157
rect 217264 51145 217270 51157
rect 217322 51145 217328 51197
rect 217378 51185 217406 51231
rect 233776 51219 233782 51231
rect 233834 51219 233840 51271
rect 247522 51259 247550 51305
rect 252034 51259 252062 51379
rect 322576 51367 322582 51419
rect 322634 51407 322640 51419
rect 329890 51407 329918 51675
rect 348400 51663 348406 51675
rect 348458 51663 348464 51715
rect 403312 51663 403318 51715
rect 403370 51703 403376 51715
rect 423376 51703 423382 51715
rect 403370 51675 423382 51703
rect 403370 51663 403376 51675
rect 423376 51663 423382 51675
rect 423434 51663 423440 51715
rect 469552 51663 469558 51715
rect 469610 51703 469616 51715
rect 483856 51703 483862 51715
rect 469610 51675 483862 51703
rect 469610 51663 469616 51675
rect 483856 51663 483862 51675
rect 483914 51663 483920 51715
rect 513250 51675 524222 51703
rect 330928 51589 330934 51641
rect 330986 51629 330992 51641
rect 348304 51629 348310 51641
rect 330986 51601 348310 51629
rect 330986 51589 330992 51601
rect 348304 51589 348310 51601
rect 348362 51589 348368 51641
rect 348496 51589 348502 51641
rect 348554 51629 348560 51641
rect 372016 51629 372022 51641
rect 348554 51601 372022 51629
rect 348554 51589 348560 51601
rect 372016 51589 372022 51601
rect 372074 51589 372080 51641
rect 382978 51601 383102 51629
rect 372112 51515 372118 51567
rect 372170 51555 372176 51567
rect 382978 51555 383006 51601
rect 372170 51527 383006 51555
rect 383074 51555 383102 51601
rect 432784 51589 432790 51641
rect 432842 51629 432848 51641
rect 452656 51629 452662 51641
rect 432842 51601 452662 51629
rect 432842 51589 432848 51601
rect 452656 51589 452662 51601
rect 452714 51589 452720 51641
rect 469360 51629 469366 51641
rect 463618 51601 469366 51629
rect 403120 51555 403126 51567
rect 383074 51527 403126 51555
rect 372170 51515 372176 51527
rect 403120 51515 403126 51527
rect 403178 51515 403184 51567
rect 452752 51515 452758 51567
rect 452810 51555 452816 51567
rect 463618 51555 463646 51601
rect 469360 51589 469366 51601
rect 469418 51589 469424 51641
rect 503938 51601 504062 51629
rect 452810 51527 463646 51555
rect 452810 51515 452816 51527
rect 493840 51515 493846 51567
rect 493898 51555 493904 51567
rect 503938 51555 503966 51601
rect 493898 51527 503966 51555
rect 504034 51555 504062 51601
rect 513250 51555 513278 51675
rect 504034 51527 513278 51555
rect 524194 51555 524222 51675
rect 552784 51663 552790 51715
rect 552842 51703 552848 51715
rect 610480 51703 610486 51715
rect 552842 51675 564542 51703
rect 552842 51663 552848 51675
rect 544336 51589 544342 51641
rect 544394 51589 544400 51641
rect 544354 51555 544382 51589
rect 524194 51527 544382 51555
rect 564514 51555 564542 51675
rect 593986 51675 610486 51703
rect 593986 51555 594014 51675
rect 610480 51663 610486 51675
rect 610538 51663 610544 51715
rect 610672 51589 610678 51641
rect 610730 51629 610736 51641
rect 625744 51629 625750 51641
rect 610730 51601 625750 51629
rect 610730 51589 610736 51601
rect 625744 51589 625750 51601
rect 625802 51589 625808 51641
rect 564514 51527 594014 51555
rect 493898 51515 493904 51527
rect 322634 51379 329918 51407
rect 322634 51367 322640 51379
rect 247522 51231 252062 51259
rect 235408 51185 235414 51197
rect 217378 51157 235414 51185
rect 235408 51145 235414 51157
rect 235466 51145 235472 51197
rect 146128 51071 146134 51123
rect 146186 51111 146192 51123
rect 232336 51111 232342 51123
rect 146186 51083 232342 51111
rect 146186 51071 146192 51083
rect 232336 51071 232342 51083
rect 232394 51071 232400 51123
rect 146224 50997 146230 51049
rect 146282 51037 146288 51049
rect 232720 51037 232726 51049
rect 146282 51009 232726 51037
rect 146282 50997 146288 51009
rect 232720 50997 232726 51009
rect 232778 50997 232784 51049
rect 146416 50923 146422 50975
rect 146474 50963 146480 50975
rect 231952 50963 231958 50975
rect 146474 50935 231958 50963
rect 146474 50923 146480 50935
rect 231952 50923 231958 50935
rect 232010 50923 232016 50975
rect 146608 50849 146614 50901
rect 146666 50889 146672 50901
rect 230992 50889 230998 50901
rect 146666 50861 230998 50889
rect 146666 50849 146672 50861
rect 230992 50849 230998 50861
rect 231050 50849 231056 50901
rect 146800 50775 146806 50827
rect 146858 50815 146864 50827
rect 230608 50815 230614 50827
rect 146858 50787 230614 50815
rect 146858 50775 146864 50787
rect 230608 50775 230614 50787
rect 230666 50775 230672 50827
rect 144880 50701 144886 50753
rect 144938 50741 144944 50753
rect 228784 50741 228790 50753
rect 144938 50713 228790 50741
rect 144938 50701 144944 50713
rect 228784 50701 228790 50713
rect 228842 50701 228848 50753
rect 145072 50627 145078 50679
rect 145130 50667 145136 50679
rect 228304 50667 228310 50679
rect 145130 50639 228310 50667
rect 145130 50627 145136 50639
rect 228304 50627 228310 50639
rect 228362 50627 228368 50679
rect 145264 50553 145270 50605
rect 145322 50593 145328 50605
rect 229744 50593 229750 50605
rect 145322 50565 229750 50593
rect 145322 50553 145328 50565
rect 229744 50553 229750 50565
rect 229802 50553 229808 50605
rect 145168 50479 145174 50531
rect 145226 50519 145232 50531
rect 229360 50519 229366 50531
rect 145226 50491 229366 50519
rect 145226 50479 145232 50491
rect 229360 50479 229366 50491
rect 229418 50479 229424 50531
rect 145456 50405 145462 50457
rect 145514 50445 145520 50457
rect 228400 50445 228406 50457
rect 145514 50417 228406 50445
rect 145514 50405 145520 50417
rect 228400 50405 228406 50417
rect 228458 50405 228464 50457
rect 144496 50331 144502 50383
rect 144554 50371 144560 50383
rect 208144 50371 208150 50383
rect 144554 50343 208150 50371
rect 144554 50331 144560 50343
rect 208144 50331 208150 50343
rect 208202 50331 208208 50383
rect 208240 50331 208246 50383
rect 208298 50371 208304 50383
rect 216880 50371 216886 50383
rect 208298 50343 216886 50371
rect 208298 50331 208304 50343
rect 216880 50331 216886 50343
rect 216938 50331 216944 50383
rect 146032 50257 146038 50309
rect 146090 50297 146096 50309
rect 207952 50297 207958 50309
rect 146090 50269 207958 50297
rect 146090 50257 146096 50269
rect 207952 50257 207958 50269
rect 208010 50257 208016 50309
rect 224272 50297 224278 50309
rect 217186 50269 224278 50297
rect 144208 50183 144214 50235
rect 144266 50223 144272 50235
rect 217186 50223 217214 50269
rect 224272 50257 224278 50269
rect 224330 50257 224336 50309
rect 144266 50195 217214 50223
rect 144266 50183 144272 50195
rect 217264 50183 217270 50235
rect 217322 50223 217328 50235
rect 235984 50223 235990 50235
rect 217322 50195 235990 50223
rect 217322 50183 217328 50195
rect 235984 50183 235990 50195
rect 236042 50183 236048 50235
rect 144976 50109 144982 50161
rect 145034 50149 145040 50161
rect 234544 50149 234550 50161
rect 145034 50121 234550 50149
rect 145034 50109 145040 50121
rect 234544 50109 234550 50121
rect 234602 50109 234608 50161
rect 145840 50035 145846 50087
rect 145898 50075 145904 50087
rect 234928 50075 234934 50087
rect 145898 50047 234934 50075
rect 145898 50035 145904 50047
rect 234928 50035 234934 50047
rect 234986 50035 234992 50087
rect 144112 49961 144118 50013
rect 144170 50001 144176 50013
rect 237232 50001 237238 50013
rect 144170 49973 237238 50001
rect 144170 49961 144176 49973
rect 237232 49961 237238 49973
rect 237290 49961 237296 50013
rect 146320 49887 146326 49939
rect 146378 49927 146384 49939
rect 232816 49927 232822 49939
rect 146378 49899 232822 49927
rect 146378 49887 146384 49899
rect 232816 49887 232822 49899
rect 232874 49887 232880 49939
rect 209104 49813 209110 49865
rect 209162 49853 209168 49865
rect 221488 49853 221494 49865
rect 209162 49825 221494 49853
rect 209162 49813 209168 49825
rect 221488 49813 221494 49825
rect 221546 49813 221552 49865
rect 208144 49739 208150 49791
rect 208202 49779 208208 49791
rect 225328 49779 225334 49791
rect 208202 49751 225334 49779
rect 208202 49739 208208 49751
rect 225328 49739 225334 49751
rect 225386 49739 225392 49791
rect 207952 49665 207958 49717
rect 208010 49705 208016 49717
rect 226576 49705 226582 49717
rect 208010 49677 226582 49705
rect 208010 49665 208016 49677
rect 226576 49665 226582 49677
rect 226634 49665 226640 49717
rect 208336 49591 208342 49643
rect 208394 49631 208400 49643
rect 219472 49631 219478 49643
rect 208394 49603 219478 49631
rect 208394 49591 208400 49603
rect 219472 49591 219478 49603
rect 219530 49591 219536 49643
rect 223696 48925 223702 48977
rect 223754 48965 223760 48977
rect 229648 48965 229654 48977
rect 223754 48937 229654 48965
rect 223754 48925 223760 48937
rect 229648 48925 229654 48937
rect 229706 48925 229712 48977
rect 208528 48851 208534 48903
rect 208586 48891 208592 48903
rect 220528 48891 220534 48903
rect 208586 48863 220534 48891
rect 208586 48851 208592 48863
rect 220528 48851 220534 48863
rect 220586 48851 220592 48903
rect 222928 48851 222934 48903
rect 222986 48891 222992 48903
rect 645328 48891 645334 48903
rect 222986 48863 645334 48891
rect 222986 48851 222992 48863
rect 645328 48851 645334 48863
rect 645386 48851 645392 48903
rect 209008 48777 209014 48829
rect 209066 48817 209072 48829
rect 222064 48817 222070 48829
rect 209066 48789 222070 48817
rect 209066 48777 209072 48789
rect 222064 48777 222070 48789
rect 222122 48777 222128 48829
rect 222256 48777 222262 48829
rect 222314 48817 222320 48829
rect 645232 48817 645238 48829
rect 222314 48789 645238 48817
rect 222314 48777 222320 48789
rect 645232 48777 645238 48789
rect 645290 48777 645296 48829
rect 208624 48703 208630 48755
rect 208682 48743 208688 48755
rect 221680 48743 221686 48755
rect 208682 48715 221686 48743
rect 208682 48703 208688 48715
rect 221680 48703 221686 48715
rect 221738 48703 221744 48755
rect 224080 48703 224086 48755
rect 224138 48743 224144 48755
rect 645136 48743 645142 48755
rect 224138 48715 645142 48743
rect 224138 48703 224144 48715
rect 645136 48703 645142 48715
rect 645194 48703 645200 48755
rect 208912 48629 208918 48681
rect 208970 48669 208976 48681
rect 222352 48669 222358 48681
rect 208970 48641 222358 48669
rect 208970 48629 208976 48641
rect 222352 48629 222358 48641
rect 222410 48629 222416 48681
rect 148432 48555 148438 48607
rect 148490 48595 148496 48607
rect 235024 48595 235030 48607
rect 148490 48567 235030 48595
rect 148490 48555 148496 48567
rect 235024 48555 235030 48567
rect 235082 48555 235088 48607
rect 208816 48481 208822 48533
rect 208874 48521 208880 48533
rect 222736 48521 222742 48533
rect 208874 48493 222742 48521
rect 208874 48481 208880 48493
rect 222736 48481 222742 48493
rect 222794 48481 222800 48533
rect 188560 48407 188566 48459
rect 188618 48447 188624 48459
rect 241168 48447 241174 48459
rect 188618 48419 241174 48447
rect 188618 48407 188624 48419
rect 241168 48407 241174 48419
rect 241226 48407 241232 48459
rect 208720 48333 208726 48385
rect 208778 48373 208784 48385
rect 223888 48373 223894 48385
rect 208778 48345 223894 48373
rect 208778 48333 208784 48345
rect 223888 48333 223894 48345
rect 223946 48333 223952 48385
rect 197200 48259 197206 48311
rect 197258 48299 197264 48311
rect 241552 48299 241558 48311
rect 197258 48271 241558 48299
rect 197258 48259 197264 48271
rect 241552 48259 241558 48271
rect 241610 48259 241616 48311
rect 149104 48185 149110 48237
rect 149162 48225 149168 48237
rect 226096 48225 226102 48237
rect 149162 48197 226102 48225
rect 149162 48185 149168 48197
rect 226096 48185 226102 48197
rect 226154 48185 226160 48237
rect 149200 48111 149206 48163
rect 149258 48151 149264 48163
rect 224560 48151 224566 48163
rect 149258 48123 224566 48151
rect 149258 48111 149264 48123
rect 224560 48111 224566 48123
rect 224618 48111 224624 48163
rect 149392 48037 149398 48089
rect 149450 48077 149456 48089
rect 223120 48077 223126 48089
rect 149450 48049 223126 48077
rect 149450 48037 149456 48049
rect 223120 48037 223126 48049
rect 223178 48037 223184 48089
rect 149296 47963 149302 48015
rect 149354 48003 149360 48015
rect 223504 48003 223510 48015
rect 149354 47975 223510 48003
rect 149354 47963 149360 47975
rect 223504 47963 223510 47975
rect 223562 47963 223568 48015
rect 149584 47889 149590 47941
rect 149642 47929 149648 47941
rect 220144 47929 220150 47941
rect 149642 47901 220150 47929
rect 149642 47889 149648 47901
rect 220144 47889 220150 47901
rect 220202 47889 220208 47941
rect 149488 47815 149494 47867
rect 149546 47855 149552 47867
rect 221296 47855 221302 47867
rect 149546 47827 221302 47855
rect 149546 47815 149552 47827
rect 221296 47815 221302 47827
rect 221354 47815 221360 47867
rect 149680 47741 149686 47793
rect 149738 47781 149744 47793
rect 219088 47781 219094 47793
rect 149738 47753 219094 47781
rect 149738 47741 149744 47753
rect 219088 47741 219094 47753
rect 219146 47741 219152 47793
rect 147760 47667 147766 47719
rect 147818 47707 147824 47719
rect 216496 47707 216502 47719
rect 147818 47679 216502 47707
rect 147818 47667 147824 47679
rect 216496 47667 216502 47679
rect 216554 47667 216560 47719
rect 147856 47593 147862 47645
rect 147914 47633 147920 47645
rect 217648 47633 217654 47645
rect 147914 47605 217654 47633
rect 147914 47593 147920 47605
rect 217648 47593 217654 47605
rect 217706 47593 217712 47645
rect 147952 47519 147958 47571
rect 148010 47559 148016 47571
rect 217936 47559 217942 47571
rect 148010 47531 217942 47559
rect 148010 47519 148016 47531
rect 217936 47519 217942 47531
rect 217994 47519 218000 47571
rect 514000 47519 514006 47571
rect 514058 47559 514064 47571
rect 525904 47559 525910 47571
rect 514058 47531 525910 47559
rect 514058 47519 514064 47531
rect 525904 47519 525910 47531
rect 525962 47519 525968 47571
rect 148048 47445 148054 47497
rect 148106 47485 148112 47497
rect 218320 47485 218326 47497
rect 148106 47457 218326 47485
rect 148106 47445 148112 47457
rect 218320 47445 218326 47457
rect 218378 47445 218384 47497
rect 148144 47371 148150 47423
rect 148202 47411 148208 47423
rect 218704 47411 218710 47423
rect 148202 47383 218710 47411
rect 148202 47371 148208 47383
rect 218704 47371 218710 47383
rect 218762 47371 218768 47423
rect 179920 47297 179926 47349
rect 179978 47337 179984 47349
rect 238576 47337 238582 47349
rect 179978 47309 238582 47337
rect 179978 47297 179984 47309
rect 238576 47297 238582 47309
rect 238634 47297 238640 47349
rect 185680 47223 185686 47275
rect 185738 47263 185744 47275
rect 240400 47263 240406 47275
rect 185738 47235 240406 47263
rect 185738 47223 185744 47235
rect 240400 47223 240406 47235
rect 240458 47223 240464 47275
rect 202960 47149 202966 47201
rect 203018 47189 203024 47201
rect 239344 47189 239350 47201
rect 203018 47161 239350 47189
rect 203018 47149 203024 47161
rect 239344 47149 239350 47161
rect 239402 47149 239408 47201
rect 148816 47075 148822 47127
rect 148874 47115 148880 47127
rect 233296 47115 233302 47127
rect 148874 47087 233302 47115
rect 148874 47075 148880 47087
rect 233296 47075 233302 47087
rect 233354 47075 233360 47127
rect 200080 47001 200086 47053
rect 200138 47041 200144 47053
rect 238960 47041 238966 47053
rect 200138 47013 238966 47041
rect 200138 47001 200144 47013
rect 238960 47001 238966 47013
rect 239018 47001 239024 47053
rect 194320 46927 194326 46979
rect 194378 46967 194384 46979
rect 240784 46967 240790 46979
rect 194378 46939 240790 46967
rect 194378 46927 194384 46939
rect 240784 46927 240790 46939
rect 240842 46927 240848 46979
rect 148912 46853 148918 46905
rect 148970 46893 148976 46905
rect 230128 46893 230134 46905
rect 148970 46865 230134 46893
rect 148970 46853 148976 46865
rect 230128 46853 230134 46865
rect 230186 46853 230192 46905
rect 148528 46779 148534 46831
rect 148586 46819 148592 46831
rect 231568 46819 231574 46831
rect 148586 46791 231574 46819
rect 148586 46779 148592 46791
rect 231568 46779 231574 46791
rect 231626 46779 231632 46831
rect 207856 46705 207862 46757
rect 207914 46745 207920 46757
rect 224944 46745 224950 46757
rect 207914 46717 224950 46745
rect 207914 46705 207920 46717
rect 224944 46705 224950 46717
rect 225002 46705 225008 46757
rect 225040 46705 225046 46757
rect 225098 46745 225104 46757
rect 227920 46745 227926 46757
rect 225098 46717 227926 46745
rect 225098 46705 225104 46717
rect 227920 46705 227926 46717
rect 227978 46705 227984 46757
rect 149008 46631 149014 46683
rect 149066 46671 149072 46683
rect 226480 46671 226486 46683
rect 149066 46643 226486 46671
rect 149066 46631 149072 46643
rect 226480 46631 226486 46643
rect 226538 46631 226544 46683
rect 148720 46557 148726 46609
rect 148778 46597 148784 46609
rect 234160 46597 234166 46609
rect 148778 46569 234166 46597
rect 148778 46557 148784 46569
rect 234160 46557 234166 46569
rect 234218 46557 234224 46609
rect 148624 46483 148630 46535
rect 148682 46523 148688 46535
rect 230512 46523 230518 46535
rect 148682 46495 230518 46523
rect 148682 46483 148688 46495
rect 230512 46483 230518 46495
rect 230570 46483 230576 46535
rect 218512 46409 218518 46461
rect 218570 46449 218576 46461
rect 645616 46449 645622 46461
rect 218570 46421 645622 46449
rect 218570 46409 218576 46421
rect 645616 46409 645622 46421
rect 645674 46409 645680 46461
rect 159760 46335 159766 46387
rect 159818 46375 159824 46387
rect 239440 46375 239446 46387
rect 159818 46347 239446 46375
rect 159818 46335 159824 46347
rect 239440 46335 239446 46347
rect 239498 46335 239504 46387
rect 207760 46261 207766 46313
rect 207818 46301 207824 46313
rect 225040 46301 225046 46313
rect 207818 46273 225046 46301
rect 207818 46261 207824 46273
rect 225040 46261 225046 46273
rect 225098 46261 225104 46313
rect 148240 46187 148246 46239
rect 148298 46227 148304 46239
rect 236752 46227 236758 46239
rect 148298 46199 236758 46227
rect 148298 46187 148304 46199
rect 236752 46187 236758 46199
rect 236810 46187 236816 46239
rect 162640 46113 162646 46165
rect 162698 46153 162704 46165
rect 239824 46153 239830 46165
rect 162698 46125 239830 46153
rect 162698 46113 162704 46125
rect 239824 46113 239830 46125
rect 239882 46113 239888 46165
rect 293776 45817 293782 45869
rect 293834 45857 293840 45869
rect 302320 45857 302326 45869
rect 293834 45829 302326 45857
rect 293834 45817 293840 45829
rect 302320 45817 302326 45829
rect 302378 45817 302384 45869
rect 211696 45299 211702 45351
rect 211754 45339 211760 45351
rect 327280 45339 327286 45351
rect 211754 45311 327286 45339
rect 211754 45299 211760 45311
rect 327280 45299 327286 45311
rect 327338 45299 327344 45351
rect 211408 45225 211414 45277
rect 211466 45265 211472 45277
rect 328048 45265 328054 45277
rect 211466 45237 328054 45265
rect 211466 45225 211472 45237
rect 328048 45225 328054 45237
rect 328106 45225 328112 45277
rect 213904 45151 213910 45203
rect 213962 45191 213968 45203
rect 446896 45191 446902 45203
rect 213962 45163 446902 45191
rect 213962 45151 213968 45163
rect 446896 45151 446902 45163
rect 446954 45151 446960 45203
rect 214672 45077 214678 45129
rect 214730 45117 214736 45129
rect 506800 45117 506806 45129
rect 214730 45089 506806 45117
rect 214730 45077 214736 45089
rect 506800 45077 506806 45089
rect 506858 45077 506864 45129
rect 215056 45003 215062 45055
rect 215114 45043 215120 45055
rect 506704 45043 506710 45055
rect 215114 45015 506710 45043
rect 215114 45003 215120 45015
rect 506704 45003 506710 45015
rect 506762 45003 506768 45055
rect 215440 44929 215446 44981
rect 215498 44969 215504 44981
rect 526960 44969 526966 44981
rect 215498 44941 526966 44969
rect 215498 44929 215504 44941
rect 526960 44929 526966 44941
rect 527018 44929 527024 44981
rect 452176 43523 452182 43575
rect 452234 43563 452240 43575
rect 461104 43563 461110 43575
rect 452234 43535 461110 43563
rect 452234 43523 452240 43535
rect 461104 43523 461110 43535
rect 461162 43523 461168 43575
rect 213232 43227 213238 43279
rect 213290 43267 213296 43279
rect 410992 43267 410998 43279
rect 213290 43239 410998 43267
rect 213290 43227 213296 43239
rect 410992 43227 410998 43239
rect 411050 43227 411056 43279
rect 446896 43153 446902 43205
rect 446954 43193 446960 43205
rect 454960 43193 454966 43205
rect 446954 43165 454966 43193
rect 446954 43153 446960 43165
rect 454960 43153 454966 43165
rect 455018 43153 455024 43205
rect 348304 42857 348310 42909
rect 348362 42897 348368 42909
rect 357424 42897 357430 42909
rect 348362 42869 357430 42897
rect 348362 42857 348368 42869
rect 357424 42857 357430 42869
rect 357482 42857 357488 42909
rect 133648 42783 133654 42835
rect 133706 42823 133712 42835
rect 136528 42823 136534 42835
rect 133706 42795 136534 42823
rect 133706 42783 133712 42795
rect 136528 42783 136534 42795
rect 136586 42783 136592 42835
rect 212464 42339 212470 42391
rect 212522 42379 212528 42391
rect 310096 42379 310102 42391
rect 212522 42351 310102 42379
rect 212522 42339 212528 42351
rect 310096 42339 310102 42351
rect 310154 42339 310160 42391
rect 206896 42117 206902 42169
rect 206954 42157 206960 42169
rect 405232 42157 405238 42169
rect 206954 42129 405238 42157
rect 206954 42117 206960 42129
rect 405232 42117 405238 42129
rect 405290 42117 405296 42169
rect 213616 42043 213622 42095
rect 213674 42083 213680 42095
rect 460048 42083 460054 42095
rect 213674 42055 460054 42083
rect 213674 42043 213680 42055
rect 460048 42043 460054 42055
rect 460106 42043 460112 42095
rect 214288 41969 214294 42021
rect 214346 42009 214352 42021
rect 514864 42009 514870 42021
rect 214346 41981 514870 42009
rect 214346 41969 214352 41981
rect 514864 41969 514870 41981
rect 514922 41969 514928 42021
rect 521584 42009 521590 42021
rect 514978 41981 521590 42009
rect 506800 41895 506806 41947
rect 506858 41935 506864 41947
rect 514978 41935 515006 41981
rect 521584 41969 521590 41981
rect 521642 41969 521648 42021
rect 506858 41907 515006 41935
rect 506858 41895 506864 41907
rect 403408 41821 403414 41873
rect 403466 41861 403472 41873
rect 403466 41833 409406 41861
rect 403466 41821 403472 41833
rect 506704 41747 506710 41799
rect 506762 41787 506768 41799
rect 518512 41787 518518 41799
rect 506762 41759 518518 41787
rect 506762 41747 506768 41759
rect 518512 41747 518518 41759
rect 518570 41747 518576 41799
<< via1 >>
rect 93910 1010925 93962 1010977
rect 97078 1010925 97130 1010977
rect 440662 1005671 440714 1005723
rect 446614 1005671 446666 1005723
rect 93718 1005523 93770 1005575
rect 115702 1005597 115754 1005649
rect 439222 1005523 439274 1005575
rect 446422 1005523 446474 1005575
rect 97078 1005449 97130 1005501
rect 118198 1005449 118250 1005501
rect 298486 1005449 298538 1005501
rect 312790 1005449 312842 1005501
rect 365110 1005449 365162 1005501
rect 383638 1005449 383690 1005501
rect 433174 1005449 433226 1005501
rect 460822 1005449 460874 1005501
rect 558742 1005449 558794 1005501
rect 572854 1005449 572906 1005501
rect 92566 1005375 92618 1005427
rect 102166 1005375 102218 1005427
rect 298390 1005375 298442 1005427
rect 313846 1005375 313898 1005427
rect 430870 1005375 430922 1005427
rect 446038 1005375 446090 1005427
rect 446614 1005375 446666 1005427
rect 469846 1005375 469898 1005427
rect 554518 1005375 554570 1005427
rect 570454 1005375 570506 1005427
rect 92662 1005301 92714 1005353
rect 101494 1005301 101546 1005353
rect 298678 1005301 298730 1005353
rect 309622 1005301 309674 1005353
rect 358678 1005301 358730 1005353
rect 366262 1005301 366314 1005353
rect 431542 1005301 431594 1005353
rect 446326 1005301 446378 1005353
rect 446422 1005301 446474 1005353
rect 470038 1005301 470090 1005353
rect 556918 1005301 556970 1005353
rect 574486 1005301 574538 1005353
rect 92950 1005227 93002 1005279
rect 114166 1005227 114218 1005279
rect 298774 1005227 298826 1005279
rect 308758 1005227 308810 1005279
rect 318646 1005227 318698 1005279
rect 328726 1005227 328778 1005279
rect 359926 1005227 359978 1005279
rect 92470 1005153 92522 1005205
rect 105430 1005153 105482 1005205
rect 195478 1005153 195530 1005205
rect 209014 1005153 209066 1005205
rect 299542 1005153 299594 1005205
rect 310294 1005153 310346 1005205
rect 325462 1005153 325514 1005205
rect 331222 1005153 331274 1005205
rect 357046 1005153 357098 1005205
rect 368566 1005153 368618 1005205
rect 381718 1005227 381770 1005279
rect 425302 1005227 425354 1005279
rect 463606 1005227 463658 1005279
rect 500662 1005227 500714 1005279
rect 512566 1005227 512618 1005279
rect 364246 1005079 364298 1005131
rect 427606 1005153 427658 1005205
rect 466582 1005153 466634 1005205
rect 501142 1005153 501194 1005205
rect 512470 1005153 512522 1005205
rect 553750 1005153 553802 1005205
rect 558742 1005153 558794 1005205
rect 562486 1005153 562538 1005205
rect 570550 1005153 570602 1005205
rect 382966 1005079 383018 1005131
rect 435574 1005079 435626 1005131
rect 440662 1005079 440714 1005131
rect 428086 1003895 428138 1003947
rect 457846 1003895 457898 1003947
rect 357622 1003821 357674 1003873
rect 380086 1003821 380138 1003873
rect 426454 1003821 426506 1003873
rect 456310 1003821 456362 1003873
rect 554902 1003821 554954 1003873
rect 567190 1003821 567242 1003873
rect 359062 1003747 359114 1003799
rect 378262 1003747 378314 1003799
rect 423382 1003747 423434 1003799
rect 466486 1003747 466538 1003799
rect 498166 1003747 498218 1003799
rect 515734 1003747 515786 1003799
rect 92374 1003673 92426 1003725
rect 108886 1003673 108938 1003725
rect 355990 1003673 356042 1003725
rect 379318 1003673 379370 1003725
rect 425782 1003673 425834 1003725
rect 471766 1003673 471818 1003725
rect 555670 1003673 555722 1003725
rect 567286 1003673 567338 1003725
rect 501046 1002563 501098 1002615
rect 519286 1002563 519338 1002615
rect 143734 1002489 143786 1002541
rect 157942 1002489 157994 1002541
rect 503446 1002489 503498 1002541
rect 97846 1002415 97898 1002467
rect 102838 1002415 102890 1002467
rect 144022 1002415 144074 1002467
rect 151222 1002415 151274 1002467
rect 99766 1002341 99818 1002393
rect 103798 1002341 103850 1002393
rect 143926 1002341 143978 1002393
rect 150358 1002341 150410 1002393
rect 559126 1002489 559178 1002541
rect 566134 1002489 566186 1002541
rect 560566 1002415 560618 1002467
rect 566422 1002415 566474 1002467
rect 517174 1002341 517226 1002393
rect 560086 1002341 560138 1002393
rect 564694 1002341 564746 1002393
rect 564790 1002341 564842 1002393
rect 567670 1002341 567722 1002393
rect 97750 1002267 97802 1002319
rect 100534 1002267 100586 1002319
rect 100726 1002267 100778 1002319
rect 104470 1002267 104522 1002319
rect 144118 1002267 144170 1002319
rect 178486 1002267 178538 1002319
rect 446038 1002267 446090 1002319
rect 446518 1002267 446570 1002319
rect 505078 1002267 505130 1002319
rect 523606 1002267 523658 1002319
rect 561526 1002267 561578 1002319
rect 565174 1002267 565226 1002319
rect 378262 1001897 378314 1001949
rect 380470 1001897 380522 1001949
rect 446518 1001157 446570 1001209
rect 467062 1001157 467114 1001209
rect 434038 1001083 434090 1001135
rect 472630 1001083 472682 1001135
rect 195286 1001009 195338 1001061
rect 208342 1001009 208394 1001061
rect 446422 1001009 446474 1001061
rect 472342 1001009 472394 1001061
rect 564694 1001009 564746 1001061
rect 570166 1001009 570218 1001061
rect 432502 1000935 432554 1000987
rect 472630 1000935 472682 1000987
rect 361558 1000861 361610 1000913
rect 383638 1000861 383690 1000913
rect 428950 1000861 429002 1000913
rect 472534 1000861 472586 1000913
rect 565174 1000861 565226 1000913
rect 568342 1000861 568394 1000913
rect 143830 1000787 143882 1000839
rect 160246 1000787 160298 1000839
rect 195382 1000787 195434 1000839
rect 211702 1000787 211754 1000839
rect 360694 1000787 360746 1000839
rect 383542 1000787 383594 1000839
rect 424150 1000787 424202 1000839
rect 471958 1000787 472010 1000839
rect 463702 1000713 463754 1000765
rect 472150 1000713 472202 1000765
rect 509398 1000639 509450 1000691
rect 516694 1000639 516746 1000691
rect 456310 1000269 456362 1000321
rect 458806 1000269 458858 1000321
rect 298102 999973 298154 1000025
rect 308086 999973 308138 1000025
rect 503062 999899 503114 999951
rect 516694 999899 516746 999951
rect 509878 999751 509930 999803
rect 521686 999751 521738 999803
rect 298294 999677 298346 999729
rect 298582 999529 298634 999581
rect 315478 999529 315530 999581
rect 92758 999455 92810 999507
rect 97750 999455 97802 999507
rect 246934 999455 246986 999507
rect 256438 999455 256490 999507
rect 298198 999455 298250 999507
rect 314710 999455 314762 999507
rect 92854 999381 92906 999433
rect 126646 999381 126698 999433
rect 143734 999381 143786 999433
rect 156886 999381 156938 999433
rect 195766 999381 195818 999433
rect 224662 999381 224714 999433
rect 246550 999381 246602 999433
rect 259510 999381 259562 999433
rect 298102 999381 298154 999433
rect 311446 999381 311498 999433
rect 506230 999677 506282 999729
rect 516790 999677 516842 999729
rect 616054 999677 616106 999729
rect 625750 999677 625802 999729
rect 507766 999603 507818 999655
rect 521590 999603 521642 999655
rect 540310 999603 540362 999655
rect 502390 999529 502442 999581
rect 516790 999529 516842 999581
rect 466582 999455 466634 999507
rect 472438 999455 472490 999507
rect 508630 999455 508682 999507
rect 523990 999455 524042 999507
rect 331798 999381 331850 999433
rect 399958 999381 400010 999433
rect 471670 999381 471722 999433
rect 488950 999381 489002 999433
rect 368566 999307 368618 999359
rect 383062 999307 383114 999359
rect 422518 999307 422570 999359
rect 429142 999307 429194 999359
rect 497590 999307 497642 999359
rect 516886 999307 516938 999359
rect 552982 999381 553034 999433
rect 555862 999381 555914 999433
rect 616150 999603 616202 999655
rect 625846 999603 625898 999655
rect 600406 999529 600458 999581
rect 598774 999455 598826 999507
rect 616054 999455 616106 999507
rect 625654 999455 625706 999507
rect 572470 999381 572522 999433
rect 596086 999381 596138 999433
rect 616150 999381 616202 999433
rect 616246 999381 616298 999433
rect 625846 999381 625898 999433
rect 521302 999307 521354 999359
rect 366262 999233 366314 999285
rect 383254 999233 383306 999285
rect 512470 999233 512522 999285
rect 521782 999233 521834 999285
rect 566134 999233 566186 999285
rect 573046 999233 573098 999285
rect 567190 999159 567242 999211
rect 575350 999159 575402 999211
rect 460822 999085 460874 999137
rect 471862 999085 471914 999137
rect 567382 998567 567434 998619
rect 575446 998567 575498 998619
rect 568342 998271 568394 998323
rect 572950 998271 573002 998323
rect 320950 997901 321002 997953
rect 367894 997901 367946 997953
rect 380182 997901 380234 997953
rect 572470 997901 572522 997953
rect 617782 997901 617834 997953
rect 331798 997827 331850 997879
rect 383158 997827 383210 997879
rect 557302 997827 557354 997879
rect 596086 997827 596138 997879
rect 302422 997753 302474 997805
rect 348694 997753 348746 997805
rect 566422 997753 566474 997805
rect 598774 997753 598826 997805
rect 328726 997679 328778 997731
rect 369046 997679 369098 997731
rect 457942 997679 457994 997731
rect 472246 997679 472298 997731
rect 574486 997679 574538 997731
rect 619126 997679 619178 997731
rect 570550 997605 570602 997657
rect 600406 997605 600458 997657
rect 570454 997531 570506 997583
rect 616246 997531 616298 997583
rect 458806 996791 458858 996843
rect 472054 996791 472106 996843
rect 195190 996495 195242 996547
rect 204214 996495 204266 996547
rect 251254 996495 251306 996547
rect 263062 996495 263114 996547
rect 512662 996495 512714 996547
rect 521494 996495 521546 996547
rect 555862 996495 555914 996547
rect 561430 996495 561482 996547
rect 319798 996421 319850 996473
rect 367126 996421 367178 996473
rect 604822 996347 604874 996399
rect 624886 996347 624938 996399
rect 511894 996199 511946 996251
rect 115318 996051 115370 996103
rect 127510 996051 127562 996103
rect 163126 996125 163178 996177
rect 214102 996125 214154 996177
rect 265942 996125 265994 996177
rect 127414 995977 127466 996029
rect 93910 995829 93962 995881
rect 97846 995829 97898 995881
rect 115222 995829 115274 995881
rect 127414 995829 127466 995881
rect 127510 995829 127562 995881
rect 162262 996051 162314 996103
rect 213334 996051 213386 996103
rect 215638 996051 215690 996103
rect 266998 996051 267050 996103
rect 270742 996125 270794 996177
rect 318646 996125 318698 996177
rect 368662 996125 368714 996177
rect 436342 996125 436394 996177
rect 436438 996125 436490 996177
rect 513430 996125 513482 996177
rect 563734 996125 563786 996177
rect 317110 996051 317162 996103
rect 320950 996051 321002 996103
rect 380182 996051 380234 996103
rect 440662 996051 440714 996103
rect 470038 996051 470090 996103
rect 511126 996051 511178 996103
rect 562870 996051 562922 996103
rect 164086 995977 164138 996029
rect 164182 995977 164234 996029
rect 215446 995977 215498 996029
rect 81622 995755 81674 995807
rect 89014 995755 89066 995807
rect 91510 995755 91562 995807
rect 92470 995755 92522 995807
rect 106102 995755 106154 995807
rect 113302 995755 113354 995807
rect 113398 995755 113450 995807
rect 118102 995755 118154 995807
rect 137590 995755 137642 995807
rect 89782 995681 89834 995733
rect 92374 995681 92426 995733
rect 133654 995681 133706 995733
rect 151990 995903 152042 995955
rect 198646 995903 198698 995955
rect 203446 995903 203498 995955
rect 213046 995903 213098 995955
rect 217078 995903 217130 995955
rect 264694 995977 264746 996029
rect 267766 995977 267818 996029
rect 267862 995977 267914 996029
rect 316342 995977 316394 996029
rect 319702 995977 319754 996029
rect 367126 995977 367178 996029
rect 434134 995977 434186 996029
rect 439222 995977 439274 996029
rect 469846 995977 469898 996029
rect 511894 995977 511946 996029
rect 513334 995977 513386 996029
rect 564790 995977 564842 996029
rect 144022 995829 144074 995881
rect 155350 995829 155402 995881
rect 195478 995829 195530 995881
rect 213334 995829 213386 995881
rect 250486 995903 250538 995955
rect 258838 995903 258890 995955
rect 250102 995829 250154 995881
rect 255574 995829 255626 995881
rect 299446 995903 299498 995955
rect 472054 995903 472106 995955
rect 298774 995829 298826 995881
rect 382966 995829 383018 995881
rect 472438 995829 472490 995881
rect 524086 995903 524138 995955
rect 523702 995829 523754 995881
rect 142966 995755 143018 995807
rect 143734 995755 143786 995807
rect 146806 995755 146858 995807
rect 154294 995755 154346 995807
rect 164086 995755 164138 995807
rect 165622 995755 165674 995807
rect 187702 995755 187754 995807
rect 190582 995755 190634 995807
rect 204982 995755 205034 995807
rect 224662 995755 224714 995807
rect 141046 995681 141098 995733
rect 143830 995681 143882 995733
rect 151702 995681 151754 995733
rect 156310 995681 156362 995733
rect 163990 995681 164042 995733
rect 166198 995681 166250 995733
rect 188086 995681 188138 995733
rect 202870 995681 202922 995733
rect 194422 995607 194474 995659
rect 195286 995607 195338 995659
rect 201622 995607 201674 995659
rect 206998 995607 207050 995659
rect 236470 995755 236522 995807
rect 254806 995755 254858 995807
rect 268246 995755 268298 995807
rect 273718 995755 273770 995807
rect 283798 995755 283850 995807
rect 289462 995755 289514 995807
rect 291190 995755 291242 995807
rect 305590 995755 305642 995807
rect 366646 995755 366698 995807
rect 371830 995755 371882 995807
rect 383638 995755 383690 995807
rect 384982 995755 385034 995807
rect 387478 995755 387530 995807
rect 396598 995755 396650 995807
rect 399958 995755 400010 995807
rect 438742 995755 438794 995807
rect 444502 995755 444554 995807
rect 472630 995755 472682 995807
rect 473302 995755 473354 995807
rect 477718 995755 477770 995807
rect 483862 995755 483914 995807
rect 485686 995755 485738 995807
rect 488950 995755 489002 995807
rect 504694 995755 504746 995807
rect 518710 995755 518762 995807
rect 523894 995755 523946 995807
rect 525334 995755 525386 995807
rect 529846 995755 529898 995807
rect 567094 995903 567146 995955
rect 570262 995903 570314 995955
rect 625846 995903 625898 995955
rect 562870 995829 562922 995881
rect 567382 995829 567434 995881
rect 619126 995829 619178 995881
rect 533398 995755 533450 995807
rect 537142 995755 537194 995807
rect 540310 995755 540362 995807
rect 566326 995755 566378 995807
rect 570358 995755 570410 995807
rect 625750 995755 625802 995807
rect 626518 995755 626570 995807
rect 630166 995755 630218 995807
rect 635254 995755 635306 995807
rect 245686 995681 245738 995733
rect 246550 995681 246602 995733
rect 247606 995681 247658 995733
rect 257494 995681 257546 995733
rect 291766 995681 291818 995733
rect 307414 995681 307466 995733
rect 365878 995681 365930 995733
rect 377398 995681 377450 995733
rect 383542 995681 383594 995733
rect 388054 995681 388106 995733
rect 472534 995681 472586 995733
rect 474070 995681 474122 995733
rect 523798 995681 523850 995733
rect 524758 995681 524810 995733
rect 563734 995681 563786 995733
rect 567478 995681 567530 995733
rect 625942 995681 625994 995733
rect 627094 995681 627146 995733
rect 237238 995607 237290 995659
rect 253078 995607 253130 995659
rect 258262 995607 258314 995659
rect 297334 995607 297386 995659
rect 298102 995607 298154 995659
rect 383734 995607 383786 995659
rect 384406 995607 384458 995659
rect 472726 995607 472778 995659
rect 474646 995607 474698 995659
rect 523606 995607 523658 995659
rect 528406 995607 528458 995659
rect 625654 995607 625706 995659
rect 627862 995607 627914 995659
rect 132406 995533 132458 995585
rect 144022 995533 144074 995585
rect 192502 995533 192554 995585
rect 195382 995533 195434 995585
rect 295414 995533 295466 995585
rect 298198 995533 298250 995585
rect 383062 995533 383114 995585
rect 392374 995533 392426 995585
rect 472342 995533 472394 995585
rect 476374 995533 476426 995585
rect 617782 995533 617834 995585
rect 629206 995533 629258 995585
rect 82294 995459 82346 995511
rect 92758 995459 92810 995511
rect 284374 995459 284426 995511
rect 133078 995385 133130 995437
rect 136246 995385 136298 995437
rect 143638 995385 143690 995437
rect 286774 995385 286826 995437
rect 293686 995459 293738 995511
rect 298006 995459 298058 995511
rect 380470 995459 380522 995511
rect 394870 995459 394922 995511
rect 466582 995459 466634 995511
rect 482710 995459 482762 995511
rect 521782 995459 521834 995511
rect 532822 995459 532874 995511
rect 146806 995311 146858 995363
rect 133990 995237 134042 995289
rect 143926 995237 143978 995289
rect 201718 995237 201770 995289
rect 206518 995237 206570 995289
rect 82582 995163 82634 995215
rect 141238 995163 141290 995215
rect 161206 995163 161258 995215
rect 181462 995163 181514 995215
rect 201526 995163 201578 995215
rect 287158 995163 287210 995215
rect 289462 995163 289514 995215
rect 298582 995385 298634 995437
rect 471958 995385 472010 995437
rect 481366 995385 481418 995437
rect 523510 995385 523562 995437
rect 531094 995385 531146 995437
rect 561718 995385 561770 995437
rect 581686 995385 581738 995437
rect 521302 995311 521354 995363
rect 640726 995311 640778 995363
rect 443542 995237 443594 995289
rect 463606 995237 463658 995289
rect 515734 995237 515786 995289
rect 642646 995237 642698 995289
rect 298678 995163 298730 995215
rect 471670 995163 471722 995215
rect 643414 995163 643466 995215
rect 69142 995089 69194 995141
rect 302422 995089 302474 995141
rect 383158 995089 383210 995141
rect 636502 995089 636554 995141
rect 118198 995015 118250 995067
rect 561526 995015 561578 995067
rect 584758 995015 584810 995067
rect 604726 995015 604778 995067
rect 247414 994941 247466 994993
rect 259126 994941 259178 994993
rect 287830 994941 287882 994993
rect 306454 994941 306506 994993
rect 290326 994793 290378 994845
rect 311926 994793 311978 994845
rect 289270 994497 289322 994549
rect 296662 994497 296714 994549
rect 131830 994127 131882 994179
rect 158806 994127 158858 994179
rect 244822 994053 244874 994105
rect 279286 994053 279338 994105
rect 234934 993905 234986 993957
rect 253078 993905 253130 993957
rect 61846 993831 61898 993883
rect 82582 993831 82634 993883
rect 238678 993831 238730 993883
rect 260758 993831 260810 993883
rect 558166 993831 558218 993883
rect 641014 993831 641066 993883
rect 77686 993757 77738 993809
rect 100726 993757 100778 993809
rect 129334 993757 129386 993809
rect 151702 993757 151754 993809
rect 180502 993757 180554 993809
rect 201622 993757 201674 993809
rect 231478 993757 231530 993809
rect 262390 993757 262442 993809
rect 78358 993683 78410 993735
rect 109846 993683 109898 993735
rect 181366 993683 181418 993735
rect 212662 993683 212714 993735
rect 232534 993683 232586 993735
rect 264022 993683 264074 993735
rect 506614 993683 506666 993735
rect 538966 993683 539018 993735
rect 77302 993609 77354 993661
rect 108214 993609 108266 993661
rect 128470 993609 128522 993661
rect 159574 993609 159626 993661
rect 179830 993609 179882 993661
rect 211030 993609 211082 993661
rect 237430 993609 237482 993661
rect 289270 993609 289322 993661
rect 362326 993609 362378 993661
rect 398806 993609 398858 993661
rect 429718 993609 429770 993661
rect 487798 993609 487850 993661
rect 531190 993609 531242 993661
rect 633046 993609 633098 993661
rect 126646 993535 126698 993587
rect 134614 993535 134666 993587
rect 186166 993535 186218 993587
rect 195766 993535 195818 993587
rect 279286 993535 279338 993587
rect 288118 993535 288170 993587
rect 390166 993535 390218 993587
rect 479158 993535 479210 993587
rect 501046 993535 501098 993587
rect 636502 993535 636554 993587
rect 643606 993535 643658 993587
rect 642646 993461 642698 993513
rect 649462 993461 649514 993513
rect 331222 992573 331274 992625
rect 332566 992573 332618 992625
rect 640726 990723 640778 990775
rect 645142 990649 645194 990701
rect 89590 990501 89642 990553
rect 93718 990501 93770 990553
rect 219478 990501 219530 990553
rect 221782 990501 221834 990553
rect 444502 990501 444554 990553
rect 462742 990501 462794 990553
rect 521398 989465 521450 989517
rect 374422 989391 374474 989443
rect 397846 989391 397898 989443
rect 154486 989317 154538 989369
rect 163990 989317 164042 989369
rect 222934 989317 222986 989369
rect 235606 989317 235658 989369
rect 273622 989317 273674 989369
rect 284278 989317 284330 989369
rect 328246 989317 328298 989369
rect 349174 989317 349226 989369
rect 377302 989317 377354 989369
rect 414070 989317 414122 989369
rect 446230 989317 446282 989369
rect 478966 989317 479018 989369
rect 518518 989317 518570 989369
rect 527638 989317 527690 989369
rect 570262 989465 570314 989517
rect 592438 989465 592490 989517
rect 573142 989391 573194 989443
rect 608758 989391 608810 989443
rect 543766 989317 543818 989369
rect 570358 989317 570410 989369
rect 624982 989317 625034 989369
rect 73462 989243 73514 989295
rect 92950 989243 93002 989295
rect 138262 989243 138314 989295
rect 164086 989243 164138 989295
rect 273718 989243 273770 989295
rect 300502 989243 300554 989295
rect 325270 989243 325322 989295
rect 365398 989243 365450 989295
rect 374518 989243 374570 989295
rect 430294 989243 430346 989295
rect 440758 989243 440810 989295
rect 495190 989243 495242 989295
rect 518710 989243 518762 989295
rect 560086 989243 560138 989295
rect 567670 989243 567722 989295
rect 658006 989243 658058 989295
rect 203158 988799 203210 988851
rect 213046 988799 213098 988851
rect 288022 988651 288074 988703
rect 299158 988651 299210 988703
rect 47638 988281 47690 988333
rect 122038 988281 122090 988333
rect 44758 988207 44810 988259
rect 186934 988207 186986 988259
rect 561526 988207 561578 988259
rect 576310 988207 576362 988259
rect 44854 988133 44906 988185
rect 251830 988133 251882 988185
rect 44950 988059 45002 988111
rect 316726 988059 316778 988111
rect 45046 987985 45098 988037
rect 381622 987985 381674 988037
rect 45142 987911 45194 987963
rect 446518 987911 446570 987963
rect 43126 987837 43178 987889
rect 511414 987837 511466 987889
rect 244726 987763 244778 987815
rect 247510 987763 247562 987815
rect 640534 987763 640586 987815
rect 649558 987763 649610 987815
rect 643606 987689 643658 987741
rect 650134 987689 650186 987741
rect 643414 987615 643466 987667
rect 649654 987615 649706 987667
rect 640918 987541 640970 987593
rect 650038 987541 650090 987593
rect 47926 986653 47978 986705
rect 115318 986653 115370 986705
rect 47734 986579 47786 986631
rect 115222 986579 115274 986631
rect 629206 986579 629258 986631
rect 649750 986579 649802 986631
rect 47446 986505 47498 986557
rect 118102 986505 118154 986557
rect 567382 986505 567434 986557
rect 660886 986505 660938 986557
rect 63286 986431 63338 986483
rect 145270 986431 145322 986483
rect 567478 986431 567530 986483
rect 660982 986431 661034 986483
rect 65206 986357 65258 986409
rect 195094 986357 195146 986409
rect 544246 986357 544298 986409
rect 650998 986357 651050 986409
rect 277942 985099 277994 985151
rect 288022 985099 288074 985151
rect 65110 984951 65162 985003
rect 94966 984951 95018 985003
rect 645142 984877 645194 984929
rect 649942 984877 649994 984929
rect 64822 984137 64874 984189
rect 69046 984137 69098 984189
rect 632374 983619 632426 983671
rect 674518 983619 674570 983671
rect 64918 983545 64970 983597
rect 244726 983545 244778 983597
rect 633046 983545 633098 983597
rect 674326 983545 674378 983597
rect 65014 983471 65066 983523
rect 277942 983471 277994 983523
rect 429142 983471 429194 983523
rect 649366 983471 649418 983523
rect 50518 973481 50570 973533
rect 59446 973481 59498 973533
rect 42166 967265 42218 967317
rect 43126 967265 43178 967317
rect 42166 960975 42218 961027
rect 42454 960975 42506 961027
rect 46102 959051 46154 959103
rect 59542 959051 59594 959103
rect 675094 958163 675146 958215
rect 675382 958163 675434 958215
rect 675190 956979 675242 957031
rect 675478 956979 675530 957031
rect 42070 955203 42122 955255
rect 42838 955203 42890 955255
rect 669526 954685 669578 954737
rect 675382 954685 675434 954737
rect 41782 954611 41834 954663
rect 41782 954389 41834 954441
rect 673942 953945 673994 953997
rect 675478 953945 675530 953997
rect 37366 952169 37418 952221
rect 41782 952169 41834 952221
rect 674038 952021 674090 952073
rect 675478 952021 675530 952073
rect 42358 948395 42410 948447
rect 53206 948395 53258 948447
rect 42646 947877 42698 947929
rect 46102 947877 46154 947929
rect 42454 947433 42506 947485
rect 57814 947433 57866 947485
rect 655222 944843 655274 944895
rect 674518 944843 674570 944895
rect 655126 944621 655178 944673
rect 674518 944621 674570 944673
rect 658006 942031 658058 942083
rect 674518 942031 674570 942083
rect 660982 941957 661034 942009
rect 674422 941957 674474 942009
rect 654454 941883 654506 941935
rect 674902 941883 674954 941935
rect 660886 941143 660938 941195
rect 674422 941143 674474 941195
rect 674038 938997 674090 939049
rect 676822 938997 676874 939049
rect 53206 933077 53258 933129
rect 59542 933077 59594 933129
rect 42358 930931 42410 930983
rect 44662 930931 44714 930983
rect 654454 927453 654506 927505
rect 666742 927453 666794 927505
rect 40054 927379 40106 927431
rect 40246 927379 40298 927431
rect 649558 927379 649610 927431
rect 679798 927379 679850 927431
rect 53398 915835 53450 915887
rect 59542 915835 59594 915887
rect 653974 915835 654026 915887
rect 660982 915835 661034 915887
rect 654454 904365 654506 904417
rect 663958 904365 664010 904417
rect 50326 901479 50378 901531
rect 59542 901479 59594 901531
rect 39958 892821 40010 892873
rect 40150 892821 40202 892873
rect 53206 887123 53258 887175
rect 59542 887123 59594 887175
rect 653974 881277 654026 881329
rect 660886 881277 660938 881329
rect 673174 872841 673226 872893
rect 675382 872841 675434 872893
rect 47542 872619 47594 872671
rect 59542 872619 59594 872671
rect 673366 872101 673418 872153
rect 675478 872101 675530 872153
rect 674038 871657 674090 871709
rect 675094 871657 675146 871709
rect 675382 871657 675434 871709
rect 674230 871435 674282 871487
rect 675190 871435 675242 871487
rect 675382 871435 675434 871487
rect 654454 869807 654506 869859
rect 663766 869807 663818 869859
rect 673078 869141 673130 869193
rect 675478 869141 675530 869193
rect 674518 868327 674570 868379
rect 675382 868327 675434 868379
rect 673270 867809 673322 867861
rect 675382 867809 675434 867861
rect 674134 866477 674186 866529
rect 675382 866477 675434 866529
rect 666646 865293 666698 865345
rect 675382 865293 675434 865345
rect 40054 863961 40106 864013
rect 40246 863961 40298 864013
rect 47446 858263 47498 858315
rect 58582 858263 58634 858315
rect 654166 858263 654218 858315
rect 661078 858263 661130 858315
rect 53302 843833 53354 843885
rect 59542 843833 59594 843885
rect 653974 835175 654026 835227
rect 669718 835175 669770 835227
rect 40246 832363 40298 832415
rect 40054 832289 40106 832341
rect 47734 829477 47786 829529
rect 59542 829477 59594 829529
rect 40054 826591 40106 826643
rect 40246 826591 40298 826643
rect 42166 823853 42218 823905
rect 53206 823853 53258 823905
rect 653974 823705 654026 823757
rect 672502 823705 672554 823757
rect 42166 823113 42218 823165
rect 47542 823113 47594 823165
rect 42166 822225 42218 822277
rect 50326 822225 50378 822277
rect 50422 815047 50474 815099
rect 59542 815047 59594 815099
rect 654454 812161 654506 812213
rect 664054 812161 664106 812213
rect 42166 810459 42218 810511
rect 43030 810459 43082 810511
rect 42454 807055 42506 807107
rect 42838 807055 42890 807107
rect 42838 805427 42890 805479
rect 53206 805427 53258 805479
rect 40150 803429 40202 803481
rect 42838 803429 42890 803481
rect 41974 802023 42026 802075
rect 42454 802023 42506 802075
rect 43414 800617 43466 800669
rect 45142 800617 45194 800669
rect 50326 800617 50378 800669
rect 59542 800617 59594 800669
rect 41494 800543 41546 800595
rect 43606 800543 43658 800595
rect 41590 800469 41642 800521
rect 43510 800469 43562 800521
rect 41878 800173 41930 800225
rect 42166 800173 42218 800225
rect 43318 800173 43370 800225
rect 41878 799951 41930 800003
rect 43030 798471 43082 798523
rect 42838 798323 42890 798375
rect 42166 798101 42218 798153
rect 42742 798027 42794 798079
rect 42070 797287 42122 797339
rect 43414 797287 43466 797339
rect 42166 796251 42218 796303
rect 42742 796251 42794 796303
rect 42742 796103 42794 796155
rect 43318 796103 43370 796155
rect 42166 794993 42218 795045
rect 43126 794993 43178 795045
rect 43126 794845 43178 794897
rect 43510 794845 43562 794897
rect 42166 792995 42218 793047
rect 42742 792995 42794 793047
rect 42742 792847 42794 792899
rect 43126 792847 43178 792899
rect 42166 790627 42218 790679
rect 42742 790627 42794 790679
rect 42166 789887 42218 789939
rect 43606 789887 43658 789939
rect 42166 789443 42218 789495
rect 42454 789443 42506 789495
rect 674038 789147 674090 789199
rect 675094 789147 675146 789199
rect 42166 787001 42218 787053
rect 42934 787001 42986 787053
rect 42166 786409 42218 786461
rect 42838 786409 42890 786461
rect 47542 786261 47594 786313
rect 59542 786261 59594 786313
rect 654070 786261 654122 786313
rect 666838 786261 666890 786313
rect 42070 785743 42122 785795
rect 42742 785743 42794 785795
rect 672310 784263 672362 784315
rect 675478 784263 675530 784315
rect 671926 783449 671978 783501
rect 675382 783449 675434 783501
rect 672790 783079 672842 783131
rect 675094 783079 675146 783131
rect 675478 783079 675530 783131
rect 672598 782931 672650 782983
rect 675382 782931 675434 782983
rect 672406 782487 672458 782539
rect 674230 782487 674282 782539
rect 675478 782487 675530 782539
rect 663862 780489 663914 780541
rect 675094 780489 675146 780541
rect 42742 780415 42794 780467
rect 47734 780415 47786 780467
rect 672886 779897 672938 779949
rect 675382 779897 675434 779949
rect 42742 779675 42794 779727
rect 50422 779675 50474 779727
rect 42742 778861 42794 778913
rect 53302 778861 53354 778913
rect 672982 778565 673034 778617
rect 675382 778565 675434 778617
rect 675094 777011 675146 777063
rect 675382 777011 675434 777063
rect 654070 774717 654122 774769
rect 666934 774717 666986 774769
rect 53494 771831 53546 771883
rect 59542 771831 59594 771883
rect 660982 767465 661034 767517
rect 674422 767465 674474 767517
rect 666742 766873 666794 766925
rect 674614 766873 674666 766925
rect 42934 765985 42986 766037
rect 43798 765985 43850 766037
rect 663958 765837 664010 765889
rect 674422 765837 674474 765889
rect 672118 763469 672170 763521
rect 674422 763469 674474 763521
rect 653974 763247 654026 763299
rect 661174 763247 661226 763299
rect 672694 763247 672746 763299
rect 673846 763247 673898 763299
rect 42166 761915 42218 761967
rect 53302 761915 53354 761967
rect 672214 760361 672266 760413
rect 673846 760361 673898 760413
rect 38998 760287 39050 760339
rect 43030 760287 43082 760339
rect 43222 757475 43274 757527
rect 45046 757475 45098 757527
rect 53686 757475 53738 757527
rect 59542 757475 59594 757527
rect 41494 757401 41546 757453
rect 43702 757401 43754 757453
rect 41398 757327 41450 757379
rect 43606 757327 43658 757379
rect 41686 757253 41738 757305
rect 43510 757253 43562 757305
rect 41878 756957 41930 757009
rect 41878 756735 41930 756787
rect 42070 754885 42122 754937
rect 43030 754885 43082 754937
rect 42166 754071 42218 754123
rect 43222 754071 43274 754123
rect 43702 751851 43754 751903
rect 43126 751777 43178 751829
rect 43414 751777 43466 751829
rect 43030 751703 43082 751755
rect 42934 751629 42986 751681
rect 43222 751629 43274 751681
rect 42166 750371 42218 750423
rect 43126 750371 43178 750423
rect 43126 750223 43178 750275
rect 43798 750223 43850 750275
rect 42070 749779 42122 749831
rect 43030 749779 43082 749831
rect 42454 749261 42506 749313
rect 43606 749261 43658 749313
rect 649654 748817 649706 748869
rect 679798 748817 679850 748869
rect 672790 748743 672842 748795
rect 673846 748743 673898 748795
rect 42166 746893 42218 746945
rect 42934 746893 42986 746945
rect 42070 746079 42122 746131
rect 42454 746079 42506 746131
rect 42166 745487 42218 745539
rect 42454 745487 42506 745539
rect 42166 743785 42218 743837
rect 43126 743785 43178 743837
rect 42070 743045 42122 743097
rect 43030 743045 43082 743097
rect 53590 743045 53642 743097
rect 59542 743045 59594 743097
rect 672406 742971 672458 743023
rect 675094 742971 675146 743023
rect 42166 742601 42218 742653
rect 42934 742601 42986 742653
rect 653974 740159 654026 740211
rect 672406 740159 672458 740211
rect 674710 738013 674762 738065
rect 675382 738013 675434 738065
rect 673846 737421 673898 737473
rect 675478 737421 675530 737473
rect 660982 737273 661034 737325
rect 674518 737273 674570 737325
rect 42838 737199 42890 737251
rect 53494 737199 53546 737251
rect 42166 736681 42218 736733
rect 53686 736681 53738 736733
rect 674614 736607 674666 736659
rect 675094 736607 675146 736659
rect 675382 736607 675434 736659
rect 42838 735645 42890 735697
rect 47542 735645 47594 735697
rect 675094 735423 675146 735475
rect 675478 735423 675530 735475
rect 673366 734757 673418 734809
rect 675382 734757 675434 734809
rect 672022 734387 672074 734439
rect 675382 734387 675434 734439
rect 673174 733573 673226 733625
rect 675478 733573 675530 733625
rect 672790 732315 672842 732367
rect 675478 732315 675530 732367
rect 674518 732019 674570 732071
rect 675382 732019 675434 732071
rect 674518 730465 674570 730517
rect 675478 730465 675530 730517
rect 47542 728615 47594 728667
rect 59542 728615 59594 728667
rect 674230 728615 674282 728667
rect 675478 728615 675530 728667
rect 675094 727875 675146 727927
rect 675574 727875 675626 727927
rect 663766 722473 663818 722525
rect 674422 722473 674474 722525
rect 660886 721881 660938 721933
rect 674710 721881 674762 721933
rect 661078 720845 661130 720897
rect 674422 720845 674474 720897
rect 672694 720253 672746 720305
rect 674710 720253 674762 720305
rect 672694 718995 672746 719047
rect 674710 718995 674762 719047
rect 42454 718699 42506 718751
rect 53494 718699 53546 718751
rect 654262 717145 654314 717197
rect 663958 717145 664010 717197
rect 40246 717071 40298 717123
rect 42454 717071 42506 717123
rect 672214 716997 672266 717049
rect 673942 716997 673994 717049
rect 43510 714259 43562 714311
rect 44950 714259 45002 714311
rect 50422 714259 50474 714311
rect 59542 714259 59594 714311
rect 41590 714037 41642 714089
rect 43702 714037 43754 714089
rect 41974 713889 42026 713941
rect 43414 713889 43466 713941
rect 41878 713815 41930 713867
rect 42070 713815 42122 713867
rect 43318 713815 43370 713867
rect 41878 713519 41930 713571
rect 42454 713223 42506 713275
rect 41878 711669 41930 711721
rect 672310 711521 672362 711573
rect 674710 711521 674762 711573
rect 43126 711447 43178 711499
rect 43606 711447 43658 711499
rect 43414 711373 43466 711425
rect 43702 711373 43754 711425
rect 42166 710855 42218 710907
rect 43510 710855 43562 710907
rect 671926 710485 671978 710537
rect 674422 710485 674474 710537
rect 42166 709893 42218 709945
rect 43126 709893 43178 709945
rect 672598 708413 672650 708465
rect 674710 708413 674762 708465
rect 42166 707377 42218 707429
rect 43318 707377 43370 707429
rect 672886 707377 672938 707429
rect 674422 707377 674474 707429
rect 672982 706785 673034 706837
rect 674710 706785 674762 706837
rect 42166 704269 42218 704321
rect 43030 704269 43082 704321
rect 43030 704121 43082 704173
rect 43414 704121 43466 704173
rect 42070 703529 42122 703581
rect 43126 703529 43178 703581
rect 43126 703381 43178 703433
rect 43606 703381 43658 703433
rect 42166 702863 42218 702915
rect 43030 702863 43082 702915
rect 649750 702715 649802 702767
rect 679798 702715 679850 702767
rect 673846 702641 673898 702693
rect 674710 702641 674762 702693
rect 42166 702419 42218 702471
rect 42742 702419 42794 702471
rect 42070 700421 42122 700473
rect 43126 700421 43178 700473
rect 42166 700051 42218 700103
rect 42454 700051 42506 700103
rect 42454 699829 42506 699881
rect 59542 699829 59594 699881
rect 42166 699163 42218 699215
rect 43030 699163 43082 699215
rect 674326 698941 674378 698993
rect 675574 698941 675626 698993
rect 654454 694057 654506 694109
rect 669814 694057 669866 694109
rect 42838 693983 42890 694035
rect 50422 693983 50474 694035
rect 672310 692873 672362 692925
rect 675382 692873 675434 692925
rect 42454 692725 42506 692777
rect 47542 692725 47594 692777
rect 672982 692429 673034 692481
rect 674710 692429 674762 692481
rect 675478 692429 675530 692481
rect 674614 692281 674666 692333
rect 675382 692281 675434 692333
rect 674806 690653 674858 690705
rect 675478 690653 675530 690705
rect 674902 689765 674954 689817
rect 675382 689765 675434 689817
rect 673078 688581 673130 688633
rect 675478 688581 675530 688633
rect 674902 687323 674954 687375
rect 675478 687323 675530 687375
rect 669622 686213 669674 686265
rect 675382 686213 675434 686265
rect 47542 685473 47594 685525
rect 59542 685473 59594 685525
rect 674422 685473 674474 685525
rect 675478 685473 675530 685525
rect 674038 683623 674090 683675
rect 675478 683623 675530 683675
rect 674902 681921 674954 681973
rect 675478 681921 675530 681973
rect 672118 681329 672170 681381
rect 673750 681329 673802 681381
rect 672502 677481 672554 677533
rect 674710 677481 674762 677533
rect 672694 676741 672746 676793
rect 673846 676741 673898 676793
rect 669718 676667 669770 676719
rect 674710 676667 674762 676719
rect 674710 676001 674762 676053
rect 674998 676001 675050 676053
rect 664054 675853 664106 675905
rect 674710 675853 674762 675905
rect 42454 675779 42506 675831
rect 53686 675779 53738 675831
rect 42166 674965 42218 675017
rect 42454 674965 42506 675017
rect 41782 674521 41834 674573
rect 41974 674521 42026 674573
rect 43606 673707 43658 673759
rect 44854 673707 44906 673759
rect 40150 672227 40202 672279
rect 41782 672227 41834 672279
rect 50422 671043 50474 671095
rect 59542 671043 59594 671095
rect 654454 671043 654506 671095
rect 661078 671043 661130 671095
rect 40918 670895 40970 670947
rect 43318 670895 43370 670947
rect 41686 670821 41738 670873
rect 42166 670821 42218 670873
rect 41878 670673 41930 670725
rect 43030 670673 43082 670725
rect 41782 670599 41834 670651
rect 43126 670599 43178 670651
rect 42454 670081 42506 670133
rect 43414 670081 43466 670133
rect 43030 668897 43082 668949
rect 42742 668675 42794 668727
rect 42838 668675 42890 668727
rect 43318 668675 43370 668727
rect 42166 668527 42218 668579
rect 43126 668527 43178 668579
rect 42166 667861 42218 667913
rect 43702 667861 43754 667913
rect 42166 666677 42218 666729
rect 43126 666677 43178 666729
rect 43606 665271 43658 665323
rect 43894 665271 43946 665323
rect 672790 665197 672842 665249
rect 673846 665197 673898 665249
rect 674038 665197 674090 665249
rect 674326 665197 674378 665249
rect 42166 664827 42218 664879
rect 43606 664827 43658 664879
rect 672022 664309 672074 664361
rect 673846 664309 673898 664361
rect 42070 664161 42122 664213
rect 43126 664161 43178 664213
rect 42166 663495 42218 663547
rect 42838 663495 42890 663547
rect 674614 660905 674666 660957
rect 674998 660905 675050 660957
rect 42070 660831 42122 660883
rect 42742 660831 42794 660883
rect 42166 659647 42218 659699
rect 42838 659647 42890 659699
rect 42070 657353 42122 657405
rect 42454 657353 42506 657405
rect 674902 656761 674954 656813
rect 675478 656761 675530 656813
rect 42454 656687 42506 656739
rect 59542 656687 59594 656739
rect 649846 656687 649898 656739
rect 679702 656687 679754 656739
rect 42166 656169 42218 656221
rect 43126 656169 43178 656221
rect 672982 653727 673034 653779
rect 674230 653727 674282 653779
rect 42454 649731 42506 649783
rect 51862 649731 51914 649783
rect 42454 649509 42506 649561
rect 50422 649509 50474 649561
rect 673366 648251 673418 648303
rect 675382 648251 675434 648303
rect 654262 648029 654314 648081
rect 672598 648029 672650 648081
rect 672214 647955 672266 648007
rect 675382 647955 675434 648007
rect 674230 647067 674282 647119
rect 675382 647067 675434 647119
rect 674806 646401 674858 646453
rect 675382 646401 675434 646453
rect 672790 644551 672842 644603
rect 675478 644551 675530 644603
rect 51862 644477 51914 644529
rect 59254 644477 59306 644529
rect 672694 644033 672746 644085
rect 675478 644033 675530 644085
rect 672886 643367 672938 643419
rect 675382 643367 675434 643419
rect 672502 642257 672554 642309
rect 675478 642257 675530 642309
rect 666742 641073 666794 641125
rect 675478 641073 675530 641125
rect 674806 638187 674858 638239
rect 675574 638187 675626 638239
rect 674710 638113 674762 638165
rect 675382 638113 675434 638165
rect 666934 632489 666986 632541
rect 674518 632489 674570 632541
rect 666838 631749 666890 631801
rect 674518 631749 674570 631801
rect 43126 630787 43178 630839
rect 43702 630787 43754 630839
rect 42454 630713 42506 630765
rect 56086 630713 56138 630765
rect 661174 630639 661226 630691
rect 674134 630639 674186 630691
rect 43414 627901 43466 627953
rect 44758 627901 44810 627953
rect 671926 627901 671978 627953
rect 673750 627901 673802 627953
rect 39862 627827 39914 627879
rect 43030 627827 43082 627879
rect 43126 627827 43178 627879
rect 43318 627827 43370 627879
rect 50422 627827 50474 627879
rect 59542 627827 59594 627879
rect 672022 627827 672074 627879
rect 673846 627827 673898 627879
rect 41494 627753 41546 627805
rect 43510 627753 43562 627805
rect 673270 627753 673322 627805
rect 675382 627753 675434 627805
rect 41686 627679 41738 627731
rect 43126 627679 43178 627731
rect 41878 627383 41930 627435
rect 41974 627383 42026 627435
rect 42934 627383 42986 627435
rect 41878 627161 41930 627213
rect 42166 625311 42218 625363
rect 43030 625311 43082 625363
rect 43030 625163 43082 625215
rect 43318 625163 43370 625215
rect 42166 624645 42218 624697
rect 43414 624645 43466 624697
rect 674902 623757 674954 623809
rect 675382 623757 675434 623809
rect 42166 623461 42218 623513
rect 42934 623461 42986 623513
rect 42934 623313 42986 623365
rect 43510 623313 43562 623365
rect 42166 622203 42218 622255
rect 43030 622203 43082 622255
rect 654358 622055 654410 622107
rect 669718 622055 669770 622107
rect 42166 620353 42218 620405
rect 43126 620353 43178 620405
rect 672310 617985 672362 618037
rect 674422 617985 674474 618037
rect 42166 617319 42218 617371
rect 43318 617319 43370 617371
rect 42166 615839 42218 615891
rect 43126 615839 43178 615891
rect 42166 614137 42218 614189
rect 43702 614137 43754 614189
rect 42742 613471 42794 613523
rect 59542 613471 59594 613523
rect 649942 613471 649994 613523
rect 679702 613471 679754 613523
rect 654358 613397 654410 613449
rect 669526 613397 669578 613449
rect 674998 613397 675050 613449
rect 675574 613397 675626 613449
rect 674230 613323 674282 613375
rect 675094 613323 675146 613375
rect 42166 607847 42218 607899
rect 42742 607847 42794 607899
rect 42742 607699 42794 607751
rect 51862 607699 51914 607751
rect 42742 606811 42794 606863
rect 53878 606811 53930 606863
rect 672982 604073 673034 604125
rect 675478 604073 675530 604125
rect 673078 603259 673130 603311
rect 675382 603259 675434 603311
rect 673750 603037 673802 603089
rect 675094 603037 675146 603089
rect 675382 603037 675434 603089
rect 671638 602889 671690 602941
rect 675478 602889 675530 602941
rect 672310 602445 672362 602497
rect 674998 602445 675050 602497
rect 675382 602445 675434 602497
rect 663766 601927 663818 601979
rect 674422 601927 674474 601979
rect 51862 601853 51914 601905
rect 59542 601853 59594 601905
rect 673558 599559 673610 599611
rect 675382 599559 675434 599611
rect 671830 599263 671882 599315
rect 675382 599263 675434 599315
rect 654454 599041 654506 599093
rect 666838 599041 666890 599093
rect 673174 598375 673226 598427
rect 675478 598375 675530 598427
rect 672118 597117 672170 597169
rect 675478 597117 675530 597169
rect 674422 596821 674474 596873
rect 675382 596821 675434 596873
rect 674902 595267 674954 595319
rect 675478 595267 675530 595319
rect 53878 587423 53930 587475
rect 58198 587423 58250 587475
rect 672406 587423 672458 587475
rect 673846 587423 673898 587475
rect 672022 586165 672074 586217
rect 673846 586165 673898 586217
rect 41878 586091 41930 586143
rect 42742 586091 42794 586143
rect 40054 585943 40106 585995
rect 41878 585943 41930 585995
rect 663958 585425 664010 585477
rect 674422 585425 674474 585477
rect 655222 584759 655274 584811
rect 674614 584759 674666 584811
rect 43126 584685 43178 584737
rect 47638 584685 47690 584737
rect 41782 584241 41834 584293
rect 43222 584241 43274 584293
rect 41974 584167 42026 584219
rect 42166 584167 42218 584219
rect 43318 584167 43370 584219
rect 41974 583945 42026 583997
rect 671734 583353 671786 583405
rect 671926 583353 671978 583405
rect 674614 583353 674666 583405
rect 672022 581873 672074 581925
rect 673270 581873 673322 581925
rect 671926 581799 671978 581851
rect 673846 581799 673898 581851
rect 43030 581503 43082 581555
rect 43318 581503 43370 581555
rect 42070 581429 42122 581481
rect 43126 581429 43178 581481
rect 42934 578395 42986 578447
rect 42070 578247 42122 578299
rect 42166 577655 42218 577707
rect 43030 577655 43082 577707
rect 654454 576027 654506 576079
rect 672406 576027 672458 576079
rect 672694 575953 672746 576005
rect 673846 575953 673898 576005
rect 672502 574325 672554 574377
rect 674422 574325 674474 574377
rect 42166 574103 42218 574155
rect 43126 574103 43178 574155
rect 42070 573215 42122 573267
rect 42454 573215 42506 573267
rect 672886 573067 672938 573119
rect 673846 573067 673898 573119
rect 672214 572845 672266 572897
rect 674422 572845 674474 572897
rect 42166 572771 42218 572823
rect 42934 572771 42986 572823
rect 42454 572623 42506 572675
rect 42934 572623 42986 572675
rect 672790 571957 672842 572009
rect 674422 571957 674474 572009
rect 42166 570995 42218 571047
rect 43030 570995 43082 571047
rect 42166 570329 42218 570381
rect 43126 570329 43178 570381
rect 42838 570255 42890 570307
rect 59542 570255 59594 570307
rect 42070 569737 42122 569789
rect 42934 569737 42986 569789
rect 650038 567369 650090 567421
rect 679798 567369 679850 567421
rect 654358 567295 654410 567347
rect 666646 567295 666698 567347
rect 34486 564483 34538 564535
rect 51862 564483 51914 564535
rect 673750 564113 673802 564165
rect 675094 564113 675146 564165
rect 42166 563447 42218 563499
rect 48886 563447 48938 563499
rect 672310 563447 672362 563499
rect 674998 563447 675050 563499
rect 51862 561523 51914 561575
rect 59446 561523 59498 561575
rect 674710 559525 674762 559577
rect 675382 559525 675434 559577
rect 675094 557823 675146 557875
rect 675382 557823 675434 557875
rect 675094 557083 675146 557135
rect 675478 557083 675530 557135
rect 660886 555825 660938 555877
rect 674998 555825 675050 555877
rect 674230 555233 674282 555285
rect 675478 555233 675530 555285
rect 674422 553753 674474 553805
rect 675478 553753 675530 553805
rect 673750 553161 673802 553213
rect 675382 553161 675434 553213
rect 654454 552939 654506 552991
rect 663958 552939 664010 552991
rect 674326 551903 674378 551955
rect 675478 551903 675530 551955
rect 674998 551607 675050 551659
rect 675382 551607 675434 551659
rect 674998 550053 675050 550105
rect 675478 550053 675530 550105
rect 674518 548203 674570 548255
rect 675478 548203 675530 548255
rect 674038 546353 674090 546405
rect 674326 546353 674378 546405
rect 43318 544799 43370 544851
rect 44566 544799 44618 544851
rect 48886 544651 48938 544703
rect 59542 544651 59594 544703
rect 41878 544503 41930 544555
rect 42166 544503 42218 544555
rect 42166 544355 42218 544407
rect 42454 544355 42506 544407
rect 40246 544207 40298 544259
rect 41014 544207 41066 544259
rect 42934 541617 42986 541669
rect 43318 541617 43370 541669
rect 654166 541543 654218 541595
rect 661174 541543 661226 541595
rect 42934 541469 42986 541521
rect 50518 541469 50570 541521
rect 655414 541469 655466 541521
rect 674326 541469 674378 541521
rect 669814 541395 669866 541447
rect 674614 541395 674666 541447
rect 41398 541321 41450 541373
rect 43510 541321 43562 541373
rect 41974 540951 42026 541003
rect 42070 540951 42122 541003
rect 42454 540951 42506 541003
rect 41974 540729 42026 540781
rect 661078 540729 661130 540781
rect 674614 540729 674666 540781
rect 671926 539841 671978 539893
rect 674614 539841 674666 539893
rect 673942 539767 673994 539819
rect 674230 539767 674282 539819
rect 674518 539249 674570 539301
rect 675094 539249 675146 539301
rect 42166 538287 42218 538339
rect 42934 538287 42986 538339
rect 42934 538139 42986 538191
rect 43318 538139 43370 538191
rect 42070 535771 42122 535823
rect 43030 535771 43082 535823
rect 43030 535623 43082 535675
rect 43510 535623 43562 535675
rect 672022 535623 672074 535675
rect 676630 535623 676682 535675
rect 671734 535549 671786 535601
rect 676534 535549 676586 535601
rect 42166 534587 42218 534639
rect 42934 534587 42986 534639
rect 42166 531479 42218 531531
rect 42454 531479 42506 531531
rect 672982 531109 673034 531161
rect 674806 531109 674858 531161
rect 42166 530887 42218 530939
rect 43030 530887 43082 530939
rect 42070 530147 42122 530199
rect 42934 530147 42986 530199
rect 43030 529925 43082 529977
rect 59542 529925 59594 529977
rect 654070 529925 654122 529977
rect 672502 529925 672554 529977
rect 674038 529925 674090 529977
rect 674422 529925 674474 529977
rect 672118 529481 672170 529533
rect 674806 529481 674858 529533
rect 42166 529407 42218 529459
rect 42454 529407 42506 529459
rect 671830 528889 671882 528941
rect 674806 528889 674858 528941
rect 671638 528001 671690 528053
rect 674806 528001 674858 528053
rect 42166 527631 42218 527683
rect 43126 527631 43178 527683
rect 42070 527187 42122 527239
rect 42934 527187 42986 527239
rect 650134 521267 650186 521319
rect 679798 521267 679850 521319
rect 41878 519787 41930 519839
rect 43030 519787 43082 519839
rect 654070 519343 654122 519395
rect 663862 519343 663914 519395
rect 53878 515495 53930 515547
rect 59542 515495 59594 515547
rect 656374 506911 656426 506963
rect 669526 506911 669578 506963
rect 47638 501139 47690 501191
rect 59542 501139 59594 501191
rect 674422 497439 674474 497491
rect 674902 497439 674954 497491
rect 672598 497291 672650 497343
rect 674422 497291 674474 497343
rect 669718 496477 669770 496529
rect 674422 496477 674474 496529
rect 655318 495515 655370 495567
rect 674710 495515 674762 495567
rect 44758 486709 44810 486761
rect 58582 486709 58634 486761
rect 654262 483823 654314 483875
rect 666934 483823 666986 483875
rect 650230 478125 650282 478177
rect 679798 478125 679850 478177
rect 44854 472353 44906 472405
rect 59542 472353 59594 472405
rect 654454 472205 654506 472257
rect 660982 472205 661034 472257
rect 50518 457923 50570 457975
rect 59542 457923 59594 457975
rect 654454 457923 654506 457975
rect 661078 457923 661130 457975
rect 654358 446379 654410 446431
rect 663862 446379 663914 446431
rect 53974 443567 54026 443619
rect 59542 443567 59594 443619
rect 42262 437129 42314 437181
rect 53878 437129 53930 437181
rect 42262 436241 42314 436293
rect 47638 436241 47690 436293
rect 654454 434909 654506 434961
rect 664054 434909 664106 434961
rect 47638 429137 47690 429189
rect 59542 429137 59594 429189
rect 654454 426177 654506 426229
rect 669622 426177 669674 426229
rect 42358 418407 42410 418459
rect 53878 418407 53930 418459
rect 37366 416483 37418 416535
rect 42454 416483 42506 416535
rect 40246 415373 40298 415425
rect 42934 415373 42986 415425
rect 40150 415151 40202 415203
rect 43030 415151 43082 415203
rect 43222 414855 43274 414907
rect 43702 414855 43754 414907
rect 37270 414707 37322 414759
rect 43222 414707 43274 414759
rect 45046 414707 45098 414759
rect 58390 414707 58442 414759
rect 41782 413375 41834 413427
rect 41782 413153 41834 413205
rect 653878 411821 653930 411873
rect 669622 411821 669674 411873
rect 42358 411451 42410 411503
rect 42166 411303 42218 411355
rect 42550 409823 42602 409875
rect 42166 409675 42218 409727
rect 42550 409675 42602 409727
rect 42166 409453 42218 409505
rect 42358 409453 42410 409505
rect 42358 409305 42410 409357
rect 42934 409305 42986 409357
rect 42934 409157 42986 409209
rect 666838 409157 666890 409209
rect 674422 409157 674474 409209
rect 655126 409083 655178 409135
rect 674710 409083 674762 409135
rect 672406 408343 672458 408395
rect 674710 408343 674762 408395
rect 42166 408195 42218 408247
rect 43126 408195 43178 408247
rect 42070 407455 42122 407507
rect 43030 407455 43082 407507
rect 42166 407011 42218 407063
rect 42358 407011 42410 407063
rect 42550 406049 42602 406101
rect 53398 406049 53450 406101
rect 42166 403829 42218 403881
rect 43222 403829 43274 403881
rect 42166 403311 42218 403363
rect 42934 403311 42986 403363
rect 56278 400351 56330 400403
rect 57622 400351 57674 400403
rect 654454 400351 654506 400403
rect 666646 400351 666698 400403
rect 42358 393913 42410 393965
rect 44854 393913 44906 393965
rect 42646 392877 42698 392929
rect 50518 392877 50570 392929
rect 42358 392285 42410 392337
rect 44758 392285 44810 392337
rect 650326 391693 650378 391745
rect 679702 391693 679754 391745
rect 654454 388807 654506 388859
rect 669718 388807 669770 388859
rect 675382 386365 675434 386417
rect 675382 386143 675434 386195
rect 44950 385921 45002 385973
rect 59254 385921 59306 385973
rect 675190 385403 675242 385455
rect 675478 385403 675530 385455
rect 674326 385107 674378 385159
rect 675190 385107 675242 385159
rect 674038 384811 674090 384863
rect 675382 384811 675434 384863
rect 673942 383109 673994 383161
rect 675286 383109 675338 383161
rect 674614 382443 674666 382495
rect 675478 382443 675530 382495
rect 654454 380075 654506 380127
rect 666742 380075 666794 380127
rect 675094 378965 675146 379017
rect 675286 378965 675338 379017
rect 674998 378151 675050 378203
rect 675382 378151 675434 378203
rect 674902 377559 674954 377611
rect 675382 377559 675434 377611
rect 674710 376819 674762 376871
rect 675478 376819 675530 376871
rect 674134 375709 674186 375761
rect 675478 375709 675530 375761
rect 42262 375191 42314 375243
rect 44758 375191 44810 375243
rect 37366 373193 37418 373245
rect 43318 373193 43370 373245
rect 40054 373045 40106 373097
rect 43030 373045 43082 373097
rect 40150 372527 40202 372579
rect 42838 372527 42890 372579
rect 40246 372231 40298 372283
rect 42934 372231 42986 372283
rect 37270 371565 37322 371617
rect 38326 371565 38378 371617
rect 47734 371565 47786 371617
rect 59542 371565 59594 371617
rect 41974 370159 42026 370211
rect 42166 369937 42218 369989
rect 42358 369937 42410 369989
rect 42358 369789 42410 369841
rect 42070 368087 42122 368139
rect 42358 368087 42410 368139
rect 42070 367347 42122 367399
rect 47446 367347 47498 367399
rect 42070 366237 42122 366289
rect 42838 366237 42890 366289
rect 654454 365793 654506 365845
rect 660982 365793 661034 365845
rect 42166 364979 42218 365031
rect 43126 364979 43178 365031
rect 661174 364905 661226 364957
rect 674710 364905 674762 364957
rect 42070 364239 42122 364291
rect 43030 364239 43082 364291
rect 663958 363869 664010 363921
rect 674422 363869 674474 363921
rect 42166 363647 42218 363699
rect 42934 363647 42986 363699
rect 672502 363277 672554 363329
rect 674710 363277 674762 363329
rect 42166 360613 42218 360665
rect 43318 360613 43370 360665
rect 56182 357357 56234 357409
rect 60214 357357 60266 357409
rect 42358 350697 42410 350749
rect 47638 350697 47690 350749
rect 42358 349957 42410 350009
rect 45046 349957 45098 350009
rect 42358 349069 42410 349121
rect 53974 349069 54026 349121
rect 650422 345591 650474 345643
rect 679798 345591 679850 345643
rect 674710 344407 674762 344459
rect 676822 344407 676874 344459
rect 50518 342779 50570 342831
rect 58390 342779 58442 342831
rect 654454 342705 654506 342757
rect 666742 342705 666794 342757
rect 674614 340929 674666 340981
rect 675478 340929 675530 340981
rect 673942 339523 673994 339575
rect 675382 339523 675434 339575
rect 674326 336563 674378 336615
rect 675382 336563 675434 336615
rect 674038 332715 674090 332767
rect 675382 332715 675434 332767
rect 674230 332345 674282 332397
rect 675478 332345 675530 332397
rect 654454 332271 654506 332323
rect 663766 332271 663818 332323
rect 42262 331975 42314 332027
rect 45046 331975 45098 332027
rect 674134 331531 674186 331583
rect 675382 331531 675434 331583
rect 41878 330643 41930 330695
rect 42550 330643 42602 330695
rect 674710 330495 674762 330547
rect 675478 330495 675530 330547
rect 37174 329755 37226 329807
rect 43126 329755 43178 329807
rect 40054 328793 40106 328845
rect 42934 328793 42986 328845
rect 39958 328497 40010 328549
rect 43318 328497 43370 328549
rect 37366 328423 37418 328475
rect 43030 328423 43082 328475
rect 40246 328349 40298 328401
rect 42838 328349 42890 328401
rect 53398 328349 53450 328401
rect 57814 328349 57866 328401
rect 41782 327017 41834 327069
rect 41782 326721 41834 326773
rect 42070 324871 42122 324923
rect 42550 324871 42602 324923
rect 42166 324131 42218 324183
rect 50326 324131 50378 324183
rect 42166 323095 42218 323147
rect 43126 323095 43178 323147
rect 42070 321763 42122 321815
rect 42550 321763 42602 321815
rect 42166 321023 42218 321075
rect 42934 321023 42986 321075
rect 42934 320875 42986 320927
rect 43318 320875 43370 320927
rect 42166 320579 42218 320631
rect 42838 320579 42890 320631
rect 655222 319691 655274 319743
rect 674422 319691 674474 319743
rect 669526 318877 669578 318929
rect 674422 318877 674474 318929
rect 42262 318729 42314 318781
rect 43030 318729 43082 318781
rect 666934 318285 666986 318337
rect 674710 318285 674762 318337
rect 42070 316583 42122 316635
rect 42934 316583 42986 316635
rect 44854 313919 44906 313971
rect 58006 313919 58058 313971
rect 42358 307481 42410 307533
rect 44950 307481 45002 307533
rect 42358 306741 42410 306793
rect 47734 306741 47786 306793
rect 42358 305483 42410 305535
rect 56278 305483 56330 305535
rect 44950 299563 45002 299615
rect 59446 299563 59498 299615
rect 650518 299563 650570 299615
rect 679798 299563 679850 299615
rect 674710 299489 674762 299541
rect 676822 299489 676874 299541
rect 674806 299415 674858 299467
rect 676918 299415 676970 299467
rect 674038 294753 674090 294805
rect 675190 294753 675242 294805
rect 674230 294235 674282 294287
rect 675094 294235 675146 294287
rect 673942 292903 673994 292955
rect 675382 292903 675434 292955
rect 674614 291719 674666 291771
rect 675094 291719 675146 291771
rect 674326 291053 674378 291105
rect 675094 291053 675146 291105
rect 41782 289795 41834 289847
rect 42262 289795 42314 289847
rect 674806 288537 674858 288589
rect 675478 288537 675530 288589
rect 42262 288019 42314 288071
rect 56278 288019 56330 288071
rect 674422 287723 674474 287775
rect 675382 287723 675434 287775
rect 674710 287353 674762 287405
rect 675478 287353 675530 287405
rect 37270 286761 37322 286813
rect 40534 286761 40586 286813
rect 674134 286539 674186 286591
rect 675382 286539 675434 286591
rect 40054 285281 40106 285333
rect 42262 285281 42314 285333
rect 40150 285207 40202 285259
rect 43126 285207 43178 285259
rect 40246 285133 40298 285185
rect 43030 285133 43082 285185
rect 45142 285133 45194 285185
rect 58102 285133 58154 285185
rect 654454 284911 654506 284963
rect 660886 284911 660938 284963
rect 41782 283801 41834 283853
rect 41782 283505 41834 283557
rect 42166 281729 42218 281781
rect 42358 281729 42410 281781
rect 42070 280101 42122 280153
rect 42358 280101 42410 280153
rect 42166 278547 42218 278599
rect 42934 278547 42986 278599
rect 64918 278547 64970 278599
rect 67606 278547 67658 278599
rect 299254 278547 299306 278599
rect 299494 278547 299546 278599
rect 226678 278473 226730 278525
rect 329782 278473 329834 278525
rect 350326 278473 350378 278525
rect 219574 278399 219626 278451
rect 326518 278399 326570 278451
rect 339862 278399 339914 278451
rect 384406 278547 384458 278599
rect 393814 278547 393866 278599
rect 407542 278547 407594 278599
rect 432406 278547 432458 278599
rect 351766 278473 351818 278525
rect 372502 278473 372554 278525
rect 372886 278473 372938 278525
rect 374614 278473 374666 278525
rect 374710 278473 374762 278525
rect 366358 278399 366410 278451
rect 378358 278399 378410 278451
rect 292054 278325 292106 278377
rect 374806 278325 374858 278377
rect 375286 278325 375338 278377
rect 380182 278399 380234 278451
rect 380278 278399 380330 278451
rect 400918 278399 400970 278451
rect 408118 278399 408170 278451
rect 378550 278325 378602 278377
rect 384694 278325 384746 278377
rect 302806 278251 302858 278303
rect 460438 278251 460490 278303
rect 293206 278177 293258 278229
rect 382006 278177 382058 278229
rect 382390 278177 382442 278229
rect 384022 278177 384074 278229
rect 384406 278177 384458 278229
rect 407542 278177 407594 278229
rect 300790 278103 300842 278155
rect 446326 278103 446378 278155
rect 301846 278029 301898 278081
rect 453238 278029 453290 278081
rect 291670 277955 291722 278007
rect 371350 277955 371402 278007
rect 371926 277955 371978 278007
rect 397366 277955 397418 278007
rect 64822 277881 64874 277933
rect 191446 277881 191498 277933
rect 287734 277881 287786 277933
rect 339094 277881 339146 277933
rect 352918 277881 352970 277933
rect 415318 277881 415370 277933
rect 569878 277881 569930 277933
rect 649462 277881 649514 277933
rect 42166 277807 42218 277859
rect 43126 277807 43178 277859
rect 283798 277807 283850 277859
rect 336310 277807 336362 277859
rect 354454 277807 354506 277859
rect 429526 277807 429578 277859
rect 288406 277733 288458 277785
rect 342742 277733 342794 277785
rect 355798 277733 355850 277785
rect 443830 277733 443882 277785
rect 289270 277659 289322 277711
rect 350038 277659 350090 277711
rect 358774 277659 358826 277711
rect 384406 277659 384458 277711
rect 384502 277659 384554 277711
rect 454774 277659 454826 277711
rect 294742 277585 294794 277637
rect 396502 277585 396554 277637
rect 289942 277511 289994 277563
rect 357238 277511 357290 277563
rect 368278 277511 368330 277563
rect 375190 277511 375242 277563
rect 375286 277511 375338 277563
rect 383830 277511 383882 277563
rect 383926 277511 383978 277563
rect 384310 277511 384362 277563
rect 384406 277511 384458 277563
rect 465526 277511 465578 277563
rect 295798 277437 295850 277489
rect 403606 277437 403658 277489
rect 42070 277363 42122 277415
rect 43030 277363 43082 277415
rect 296470 277363 296522 277415
rect 410806 277363 410858 277415
rect 240694 277289 240746 277341
rect 331318 277289 331370 277341
rect 351094 277289 351146 277341
rect 380278 277289 380330 277341
rect 380374 277289 380426 277341
rect 384118 277289 384170 277341
rect 384214 277289 384266 277341
rect 479734 277289 479786 277341
rect 297526 277215 297578 277267
rect 417910 277215 417962 277267
rect 317974 277141 318026 277193
rect 439318 277141 439370 277193
rect 298198 277067 298250 277119
rect 425014 277067 425066 277119
rect 254902 276993 254954 277045
rect 332758 276993 332810 277045
rect 360502 276993 360554 277045
rect 384214 276993 384266 277045
rect 384406 276993 384458 277045
rect 391606 276993 391658 277045
rect 297814 276919 297866 276971
rect 338134 276919 338186 276971
rect 365878 276919 365930 276971
rect 269206 276845 269258 276897
rect 334486 276845 334538 276897
rect 357718 276845 357770 276897
rect 384310 276845 384362 276897
rect 384502 276919 384554 276971
rect 508342 276919 508394 276971
rect 398998 276845 399050 276897
rect 262102 276771 262154 276823
rect 333910 276771 333962 276823
rect 362134 276771 362186 276823
rect 403222 276771 403274 276823
rect 247894 276697 247946 276749
rect 332182 276697 332234 276749
rect 349174 276697 349226 276749
rect 239446 276623 239498 276675
rect 252310 276623 252362 276675
rect 290806 276623 290858 276675
rect 364438 276623 364490 276675
rect 212182 276549 212234 276601
rect 327382 276549 327434 276601
rect 375190 276697 375242 276749
rect 379990 276697 380042 276749
rect 380086 276697 380138 276749
rect 381142 276697 381194 276749
rect 381238 276697 381290 276749
rect 372982 276623 373034 276675
rect 384502 276623 384554 276675
rect 386230 276697 386282 276749
rect 400054 276697 400106 276749
rect 386998 276549 387050 276601
rect 387190 276623 387242 276675
rect 615382 276623 615434 276675
rect 640342 276549 640394 276601
rect 194326 276475 194378 276527
rect 325750 276475 325802 276527
rect 374326 276475 374378 276527
rect 639094 276475 639146 276527
rect 42358 276401 42410 276453
rect 53590 276401 53642 276453
rect 231766 276401 231818 276453
rect 334582 276401 334634 276453
rect 365014 276401 365066 276453
rect 369142 276401 369194 276453
rect 371350 276401 371402 276453
rect 374134 276401 374186 276453
rect 374230 276401 374282 276453
rect 375478 276401 375530 276453
rect 375670 276401 375722 276453
rect 384118 276401 384170 276453
rect 384214 276401 384266 276453
rect 384886 276401 384938 276453
rect 385078 276401 385130 276453
rect 561814 276401 561866 276453
rect 232342 276327 232394 276379
rect 341782 276327 341834 276379
rect 372502 276327 372554 276379
rect 374710 276327 374762 276379
rect 375574 276327 375626 276379
rect 391702 276327 391754 276379
rect 395062 276327 395114 276379
rect 568918 276327 568970 276379
rect 244726 276253 244778 276305
rect 441718 276253 441770 276305
rect 245398 276179 245450 276231
rect 448822 276179 448874 276231
rect 233398 276105 233450 276157
rect 348982 276105 349034 276157
rect 367510 276105 367562 276157
rect 375382 276105 375434 276157
rect 376342 276105 376394 276157
rect 383926 276105 383978 276157
rect 384694 276105 384746 276157
rect 576118 276105 576170 276157
rect 246358 276031 246410 276083
rect 455926 276031 455978 276083
rect 234070 275957 234122 276009
rect 356086 275957 356138 276009
rect 368086 275957 368138 276009
rect 375670 275957 375722 276009
rect 375766 275957 375818 276009
rect 379894 275957 379946 276009
rect 379990 275957 380042 276009
rect 383542 275957 383594 276009
rect 384310 275957 384362 276009
rect 583222 275957 583274 276009
rect 247414 275883 247466 275935
rect 463126 275883 463178 275935
rect 204982 275809 205034 275861
rect 317590 275809 317642 275861
rect 317686 275809 317738 275861
rect 324022 275809 324074 275861
rect 324502 275809 324554 275861
rect 374326 275809 374378 275861
rect 374614 275809 374666 275861
rect 377974 275809 378026 275861
rect 378070 275809 378122 275861
rect 384310 275809 384362 275861
rect 384406 275809 384458 275861
rect 590326 275809 590378 275861
rect 248086 275735 248138 275787
rect 470230 275735 470282 275787
rect 235030 275661 235082 275713
rect 363190 275661 363242 275713
rect 364246 275661 364298 275713
rect 372982 275661 373034 275713
rect 374038 275661 374090 275713
rect 384406 275661 384458 275713
rect 384790 275661 384842 275713
rect 385078 275661 385130 275713
rect 385174 275661 385226 275713
rect 604630 275661 604682 275713
rect 235990 275587 236042 275639
rect 370294 275587 370346 275639
rect 377782 275587 377834 275639
rect 390550 275587 390602 275639
rect 398902 275587 398954 275639
rect 618838 275587 618890 275639
rect 226294 275513 226346 275565
rect 291862 275513 291914 275565
rect 317590 275513 317642 275565
rect 326998 275513 327050 275565
rect 327094 275513 327146 275565
rect 557014 275513 557066 275565
rect 227446 275439 227498 275491
rect 298966 275439 299018 275491
rect 315382 275439 315434 275491
rect 564214 275439 564266 275491
rect 200182 275365 200234 275417
rect 267670 275365 267722 275417
rect 267766 275365 267818 275417
rect 270262 275365 270314 275417
rect 315958 275365 316010 275417
rect 571318 275365 571370 275417
rect 236758 275291 236810 275343
rect 377494 275291 377546 275343
rect 377590 275291 377642 275343
rect 385174 275291 385226 275343
rect 385270 275291 385322 275343
rect 394486 275291 394538 275343
rect 398806 275291 398858 275343
rect 636694 275291 636746 275343
rect 196726 275217 196778 275269
rect 257590 275217 257642 275269
rect 317590 275217 317642 275269
rect 578518 275217 578570 275269
rect 228022 275143 228074 275195
rect 257494 275143 257546 275195
rect 257878 275143 257930 275195
rect 306070 275143 306122 275195
rect 314326 275143 314378 275195
rect 317686 275143 317738 275195
rect 318646 275143 318698 275195
rect 193078 275069 193130 275121
rect 257590 275069 257642 275121
rect 257782 275069 257834 275121
rect 267670 275069 267722 275121
rect 267766 275069 267818 275121
rect 272470 275069 272522 275121
rect 284950 275069 285002 275121
rect 314422 275069 314474 275121
rect 319798 275069 319850 275121
rect 338422 275143 338474 275195
rect 585622 275143 585674 275195
rect 229078 274995 229130 275047
rect 313270 274995 313322 275047
rect 318166 274995 318218 275047
rect 330166 274995 330218 275047
rect 592726 275069 592778 275121
rect 599830 274995 599882 275047
rect 243766 274921 243818 274973
rect 434518 274921 434570 274973
rect 663862 274921 663914 274973
rect 674710 274921 674762 274973
rect 242998 274847 243050 274899
rect 427414 274847 427466 274899
rect 233494 274773 233546 274825
rect 318166 274773 318218 274825
rect 318262 274773 318314 274825
rect 335638 274773 335690 274825
rect 362710 274773 362762 274825
rect 375766 274773 375818 274825
rect 377878 274773 377930 274825
rect 554710 274773 554762 274825
rect 242230 274699 242282 274751
rect 420214 274699 420266 274751
rect 241078 274625 241130 274677
rect 413206 274625 413258 274677
rect 429238 274625 429290 274677
rect 449110 274625 449162 274677
rect 153814 274551 153866 274603
rect 161206 274551 161258 274603
rect 240502 274551 240554 274603
rect 406006 274551 406058 274603
rect 619126 274551 619178 274603
rect 627286 274551 627338 274603
rect 239350 274477 239402 274529
rect 398614 274477 398666 274529
rect 238486 274403 238538 274455
rect 375574 274403 375626 274455
rect 375766 274403 375818 274455
rect 377590 274403 377642 274455
rect 237814 274329 237866 274381
rect 376342 274329 376394 274381
rect 377302 274329 377354 274381
rect 379126 274403 379178 274455
rect 379222 274403 379274 274455
rect 385078 274403 385130 274455
rect 593302 274403 593354 274455
rect 613366 274403 613418 274455
rect 378550 274329 378602 274381
rect 383734 274329 383786 274381
rect 383830 274329 383882 274381
rect 384406 274329 384458 274381
rect 384502 274329 384554 274381
rect 394390 274329 394442 274381
rect 394486 274329 394538 274381
rect 398806 274329 398858 274381
rect 230230 274255 230282 274307
rect 323638 274255 323690 274307
rect 324022 274255 324074 274307
rect 327094 274255 327146 274307
rect 230614 274181 230666 274233
rect 327478 274181 327530 274233
rect 207382 274107 207434 274159
rect 271318 274107 271370 274159
rect 276406 274107 276458 274159
rect 318262 274107 318314 274159
rect 318454 274107 318506 274159
rect 338422 274255 338474 274307
rect 368470 274255 368522 274307
rect 368854 274255 368906 274307
rect 369622 274255 369674 274307
rect 377878 274255 377930 274307
rect 377974 274255 378026 274307
rect 383926 274255 383978 274307
rect 359734 274181 359786 274233
rect 472630 274255 472682 274307
rect 384502 274181 384554 274233
rect 458326 274181 458378 274233
rect 469558 274181 469610 274233
rect 477622 274181 477674 274233
rect 552982 274181 553034 274233
rect 573046 274181 573098 274233
rect 355702 274107 355754 274159
rect 440470 274107 440522 274159
rect 214582 274033 214634 274085
rect 252214 274033 252266 274085
rect 252310 274033 252362 274085
rect 275254 274033 275306 274085
rect 287062 274033 287114 274085
rect 336694 274033 336746 274085
rect 353494 274033 353546 274085
rect 422614 274033 422666 274085
rect 661078 274033 661130 274085
rect 674710 274033 674762 274085
rect 225430 273959 225482 274011
rect 284662 273959 284714 274011
rect 317014 273959 317066 274011
rect 335446 273959 335498 274011
rect 358102 273959 358154 274011
rect 384502 273959 384554 274011
rect 384598 273959 384650 274011
rect 392854 273959 392906 274011
rect 225238 273885 225290 273937
rect 281110 273885 281162 273937
rect 301270 273885 301322 273937
rect 338710 273885 338762 273937
rect 370966 273885 371018 273937
rect 396118 273885 396170 273937
rect 224086 273811 224138 273863
rect 274006 273811 274058 273863
rect 274102 273811 274154 273863
rect 223030 273737 223082 273789
rect 158806 273663 158858 273715
rect 178294 273663 178346 273715
rect 252214 273737 252266 273789
rect 267766 273737 267818 273789
rect 269398 273737 269450 273789
rect 286006 273737 286058 273789
rect 286678 273811 286730 273863
rect 328726 273811 328778 273863
rect 343126 273811 343178 273863
rect 359638 273811 359690 273863
rect 361942 273811 361994 273863
rect 400342 273811 400394 273863
rect 370390 273737 370442 273789
rect 373366 273737 373418 273789
rect 378070 273737 378122 273789
rect 378166 273737 378218 273789
rect 383638 273737 383690 273789
rect 383734 273737 383786 273789
rect 398902 273737 398954 273789
rect 263350 273663 263402 273715
rect 267190 273663 267242 273715
rect 372406 273663 372458 273715
rect 372502 273663 372554 273715
rect 377686 273663 377738 273715
rect 143158 273589 143210 273641
rect 160726 273589 160778 273641
rect 267862 273589 267914 273641
rect 270742 273589 270794 273641
rect 270838 273589 270890 273641
rect 274102 273589 274154 273641
rect 102646 273515 102698 273567
rect 211606 273515 211658 273567
rect 228790 273515 228842 273567
rect 274198 273515 274250 273567
rect 275158 273515 275210 273567
rect 279670 273515 279722 273567
rect 67030 273441 67082 273493
rect 209686 273441 209738 273493
rect 209782 273441 209834 273493
rect 216118 273441 216170 273493
rect 218230 273441 218282 273493
rect 223990 273441 224042 273493
rect 224566 273441 224618 273493
rect 277558 273441 277610 273493
rect 278806 273441 278858 273493
rect 280054 273441 280106 273493
rect 280726 273441 280778 273493
rect 282358 273441 282410 273493
rect 284470 273441 284522 273493
rect 286006 273589 286058 273641
rect 378838 273663 378890 273715
rect 378934 273663 378986 273715
rect 379702 273663 379754 273715
rect 380086 273663 380138 273715
rect 394486 273663 394538 273715
rect 378646 273589 378698 273641
rect 379030 273589 379082 273641
rect 379126 273589 379178 273641
rect 387190 273589 387242 273641
rect 388630 273589 388682 273641
rect 391222 273589 391274 273641
rect 310870 273515 310922 273567
rect 319126 273515 319178 273567
rect 323734 273515 323786 273567
rect 323830 273515 323882 273567
rect 553462 273515 553514 273567
rect 285526 273441 285578 273493
rect 321526 273441 321578 273493
rect 321622 273441 321674 273493
rect 334102 273441 334154 273493
rect 336982 273441 337034 273493
rect 343030 273441 343082 273493
rect 347446 273441 347498 273493
rect 349846 273441 349898 273493
rect 351190 273441 351242 273493
rect 362038 273441 362090 273493
rect 368662 273441 368714 273493
rect 369142 273441 369194 273493
rect 370006 273441 370058 273493
rect 378646 273441 378698 273493
rect 379126 273441 379178 273493
rect 161014 273367 161066 273419
rect 377974 273367 378026 273419
rect 378358 273367 378410 273419
rect 389014 273367 389066 273419
rect 391222 273441 391274 273493
rect 622486 273441 622538 273493
rect 393622 273367 393674 273419
rect 393718 273367 393770 273419
rect 402550 273367 402602 273419
rect 403222 273367 403274 273419
rect 494038 273367 494090 273419
rect 144406 273293 144458 273345
rect 146806 273293 146858 273345
rect 157462 273293 157514 273345
rect 404086 273293 404138 273345
rect 664054 273293 664106 273345
rect 674710 273293 674762 273345
rect 65878 273219 65930 273271
rect 212374 273219 212426 273271
rect 213334 273219 213386 273271
rect 216694 273219 216746 273271
rect 217558 273219 217610 273271
rect 220438 273219 220490 273271
rect 229750 273219 229802 273271
rect 320374 273219 320426 273271
rect 320470 273219 320522 273271
rect 323638 273219 323690 273271
rect 323734 273219 323786 273271
rect 340534 273219 340586 273271
rect 340630 273219 340682 273271
rect 343510 273219 343562 273271
rect 344662 273219 344714 273271
rect 347734 273219 347786 273271
rect 347926 273219 347978 273271
rect 349750 273219 349802 273271
rect 349846 273219 349898 273271
rect 372694 273219 372746 273271
rect 374422 273219 374474 273271
rect 376246 273219 376298 273271
rect 376342 273219 376394 273271
rect 379318 273219 379370 273271
rect 379414 273219 379466 273271
rect 388630 273219 388682 273271
rect 388726 273219 388778 273271
rect 395350 273219 395402 273271
rect 396022 273219 396074 273271
rect 161302 273145 161354 273197
rect 147958 273071 148010 273123
rect 149686 273071 149738 273123
rect 152662 273071 152714 273123
rect 155350 273071 155402 273123
rect 156214 273071 156266 273123
rect 158326 273071 158378 273123
rect 162166 273071 162218 273123
rect 164086 273071 164138 273123
rect 164278 273145 164330 273197
rect 378358 273145 378410 273197
rect 378742 273145 378794 273197
rect 397078 273145 397130 273197
rect 397366 273145 397418 273197
rect 398710 273145 398762 273197
rect 398902 273219 398954 273271
rect 629686 273219 629738 273271
rect 399862 273145 399914 273197
rect 400342 273145 400394 273197
rect 490486 273145 490538 273197
rect 362998 273071 363050 273123
rect 363382 273071 363434 273123
rect 403318 273071 403370 273123
rect 501238 273071 501290 273123
rect 617686 273071 617738 273123
rect 139606 272997 139658 273049
rect 68182 272849 68234 272901
rect 69046 272849 69098 272901
rect 75382 272849 75434 272901
rect 77686 272849 77738 272901
rect 98038 272849 98090 272901
rect 100726 272849 100778 272901
rect 101494 272849 101546 272901
rect 103606 272849 103658 272901
rect 115798 272849 115850 272901
rect 118006 272849 118058 272901
rect 119350 272849 119402 272901
rect 120886 272849 120938 272901
rect 122902 272849 122954 272901
rect 123766 272849 123818 272901
rect 130102 272849 130154 272901
rect 132406 272849 132458 272901
rect 133558 272849 133610 272901
rect 135286 272849 135338 272901
rect 137206 272849 137258 272901
rect 138166 272849 138218 272901
rect 138358 272849 138410 272901
rect 140950 272849 141002 272901
rect 142006 272849 142058 272901
rect 143926 272849 143978 272901
rect 178486 272997 178538 273049
rect 302422 272997 302474 273049
rect 322486 272997 322538 273049
rect 339574 272997 339626 273049
rect 339766 272997 339818 273049
rect 362902 272997 362954 273049
rect 146710 272923 146762 272975
rect 158806 272923 158858 272975
rect 279382 272923 279434 272975
rect 279574 272923 279626 272975
rect 379510 272997 379562 273049
rect 379606 272997 379658 273049
rect 398614 272997 398666 273049
rect 363190 272923 363242 272975
rect 161206 272849 161258 272901
rect 378166 272849 378218 272901
rect 378742 272923 378794 272975
rect 394198 272923 394250 272975
rect 394390 272923 394442 272975
rect 540406 272997 540458 273049
rect 398998 272923 399050 272975
rect 407638 272923 407690 272975
rect 407734 272923 407786 272975
rect 533206 272923 533258 272975
rect 378934 272849 378986 272901
rect 135958 272775 136010 272827
rect 370390 272775 370442 272827
rect 373078 272775 373130 272827
rect 128950 272701 129002 272753
rect 160534 272701 160586 272753
rect 161206 272701 161258 272753
rect 378550 272701 378602 272753
rect 379318 272849 379370 272901
rect 388726 272849 388778 272901
rect 388822 272849 388874 272901
rect 392470 272775 392522 272827
rect 394486 272849 394538 272901
rect 518998 272849 519050 272901
rect 407542 272775 407594 272827
rect 407638 272775 407690 272827
rect 522550 272775 522602 272827
rect 105046 272627 105098 272679
rect 106486 272627 106538 272679
rect 114646 272627 114698 272679
rect 111094 272479 111146 272531
rect 125302 272627 125354 272679
rect 377974 272627 378026 272679
rect 378358 272627 378410 272679
rect 118102 272553 118154 272605
rect 378646 272553 378698 272605
rect 378838 272627 378890 272679
rect 391702 272701 391754 272753
rect 391798 272701 391850 272753
rect 396022 272701 396074 272753
rect 396118 272701 396170 272753
rect 504694 272701 504746 272753
rect 402358 272627 402410 272679
rect 418966 272627 419018 272679
rect 501142 272627 501194 272679
rect 505270 272627 505322 272679
rect 621238 272627 621290 272679
rect 103894 272405 103946 272457
rect 379030 272479 379082 272531
rect 373078 272405 373130 272457
rect 373174 272405 373226 272457
rect 378358 272405 378410 272457
rect 390934 272553 390986 272605
rect 379318 272479 379370 272531
rect 389878 272479 389930 272531
rect 389974 272479 390026 272531
rect 404950 272553 405002 272605
rect 405046 272553 405098 272605
rect 497590 272553 497642 272605
rect 497686 272553 497738 272605
rect 614230 272553 614282 272605
rect 393142 272479 393194 272531
rect 526102 272479 526154 272531
rect 379798 272405 379850 272457
rect 398806 272405 398858 272457
rect 107446 272257 107498 272309
rect 99190 272183 99242 272235
rect 370198 272183 370250 272235
rect 370390 272257 370442 272309
rect 378550 272183 378602 272235
rect 378646 272183 378698 272235
rect 378934 272183 378986 272235
rect 379510 272257 379562 272309
rect 391990 272331 392042 272383
rect 529750 272405 529802 272457
rect 398998 272331 399050 272383
rect 399190 272257 399242 272309
rect 399862 272257 399914 272309
rect 84886 272109 84938 272161
rect 86326 272109 86378 272161
rect 100342 272109 100394 272161
rect 379126 272109 379178 272161
rect 399670 272183 399722 272235
rect 89590 272035 89642 272087
rect 92086 272035 92138 272087
rect 145558 272035 145610 272087
rect 146710 272035 146762 272087
rect 150262 272035 150314 272087
rect 164278 272035 164330 272087
rect 165814 272035 165866 272087
rect 166966 272035 167018 272087
rect 170518 272035 170570 272087
rect 172726 272035 172778 272087
rect 174070 272035 174122 272087
rect 175510 272035 175562 272087
rect 177622 272035 177674 272087
rect 178390 272035 178442 272087
rect 180022 272035 180074 272087
rect 181366 272035 181418 272087
rect 181462 272035 181514 272087
rect 390550 272035 390602 272087
rect 400630 272109 400682 272161
rect 401302 272035 401354 272087
rect 401590 272331 401642 272383
rect 547606 272331 547658 272383
rect 560086 272331 560138 272383
rect 643894 272331 643946 272383
rect 406006 272257 406058 272309
rect 418966 272257 419018 272309
rect 486742 272257 486794 272309
rect 641494 272257 641546 272309
rect 407734 272183 407786 272235
rect 480982 272183 481034 272235
rect 634294 272183 634346 272235
rect 406102 272109 406154 272161
rect 609430 272109 609482 272161
rect 406774 272035 406826 272087
rect 409078 272035 409130 272087
rect 486838 272035 486890 272087
rect 164566 271961 164618 272013
rect 405526 271961 405578 272013
rect 411286 271961 411338 272013
rect 468982 271961 469034 272013
rect 172918 271887 172970 271939
rect 175606 271887 175658 271939
rect 176470 271887 176522 271939
rect 178486 271887 178538 271939
rect 179446 271887 179498 271939
rect 388822 271887 388874 271939
rect 388918 271887 388970 271939
rect 408214 271887 408266 271939
rect 106294 271813 106346 271865
rect 109846 271739 109898 271791
rect 190582 271739 190634 271791
rect 190774 271813 190826 271865
rect 192886 271813 192938 271865
rect 209686 271813 209738 271865
rect 213238 271813 213290 271865
rect 232438 271813 232490 271865
rect 271222 271813 271274 271865
rect 271606 271813 271658 271865
rect 279478 271813 279530 271865
rect 283798 271813 283850 271865
rect 307318 271813 307370 271865
rect 312118 271813 312170 271865
rect 321622 271813 321674 271865
rect 205846 271739 205898 271791
rect 220822 271739 220874 271791
rect 245494 271739 245546 271791
rect 250198 271739 250250 271791
rect 267958 271739 268010 271791
rect 268054 271739 268106 271791
rect 278998 271739 279050 271791
rect 283414 271739 283466 271791
rect 303670 271739 303722 271791
rect 313654 271739 313706 271791
rect 549910 271813 549962 271865
rect 321814 271739 321866 271791
rect 329878 271739 329930 271791
rect 329974 271739 330026 271791
rect 341782 271739 341834 271791
rect 347254 271739 347306 271791
rect 358486 271739 358538 271791
rect 358582 271739 358634 271791
rect 374422 271739 374474 271791
rect 375574 271739 375626 271791
rect 378070 271739 378122 271791
rect 378166 271739 378218 271791
rect 388630 271739 388682 271791
rect 388726 271739 388778 271791
rect 608182 271739 608234 271791
rect 171670 271665 171722 271717
rect 179446 271665 179498 271717
rect 175318 271591 175370 271643
rect 388822 271665 388874 271717
rect 388918 271665 388970 271717
rect 396214 271665 396266 271717
rect 397366 271665 397418 271717
rect 405046 271665 405098 271717
rect 141142 271517 141194 271569
rect 147190 271517 147242 271569
rect 178870 271517 178922 271569
rect 409270 271591 409322 271643
rect 182422 271517 182474 271569
rect 409942 271517 409994 271569
rect 124150 271443 124202 271495
rect 212182 271443 212234 271495
rect 246646 271443 246698 271495
rect 276118 271443 276170 271495
rect 282742 271443 282794 271495
rect 296662 271443 296714 271495
rect 308470 271443 308522 271495
rect 321814 271443 321866 271495
rect 323062 271443 323114 271495
rect 325558 271443 325610 271495
rect 325654 271443 325706 271495
rect 328054 271443 328106 271495
rect 328150 271443 328202 271495
rect 329014 271443 329066 271495
rect 329878 271443 329930 271495
rect 339382 271443 339434 271495
rect 346774 271443 346826 271495
rect 349654 271443 349706 271495
rect 349750 271443 349802 271495
rect 358582 271443 358634 271495
rect 362998 271443 363050 271495
rect 365398 271443 365450 271495
rect 370006 271443 370058 271495
rect 383254 271443 383306 271495
rect 383350 271443 383402 271495
rect 601078 271443 601130 271495
rect 127702 271369 127754 271421
rect 141142 271369 141194 271421
rect 151414 271369 151466 271421
rect 152566 271369 152618 271421
rect 190582 271369 190634 271421
rect 206998 271369 207050 271421
rect 207094 271369 207146 271421
rect 411958 271369 412010 271421
rect 131254 271295 131306 271347
rect 134806 270999 134858 271051
rect 168118 271295 168170 271347
rect 181462 271295 181514 271347
rect 185974 271295 186026 271347
rect 410998 271295 411050 271347
rect 147190 271221 147242 271273
rect 177046 271221 177098 271273
rect 184726 271221 184778 271273
rect 187030 271221 187082 271273
rect 195190 271221 195242 271273
rect 211894 271221 211946 271273
rect 220342 271221 220394 271273
rect 241846 271221 241898 271273
rect 271222 271221 271274 271273
rect 274678 271221 274730 271273
rect 282934 271221 282986 271273
rect 300118 271221 300170 271273
rect 316342 271221 316394 271273
rect 332278 271221 332330 271273
rect 334102 271221 334154 271273
rect 339862 271221 339914 271273
rect 349558 271221 349610 271273
rect 351190 271221 351242 271273
rect 351286 271221 351338 271273
rect 151126 271073 151178 271125
rect 211702 271147 211754 271199
rect 219766 271147 219818 271199
rect 238294 271147 238346 271199
rect 267958 271147 268010 271199
rect 276790 271147 276842 271199
rect 281206 271147 281258 271199
rect 285814 271147 285866 271199
rect 316822 271147 316874 271199
rect 327190 271147 327242 271199
rect 328342 271147 328394 271199
rect 331222 271147 331274 271199
rect 345718 271147 345770 271199
rect 151126 270777 151178 270829
rect 189622 271073 189674 271125
rect 212086 271073 212138 271125
rect 213046 271073 213098 271125
rect 189526 270999 189578 271051
rect 207094 270999 207146 271051
rect 207190 270999 207242 271051
rect 213814 270999 213866 271051
rect 195478 270925 195530 270977
rect 214486 270925 214538 270977
rect 177046 270851 177098 270903
rect 195190 270851 195242 270903
rect 199126 270851 199178 270903
rect 214966 270851 215018 270903
rect 189622 270777 189674 270829
rect 202582 270777 202634 270829
rect 215446 270777 215498 270829
rect 67606 270703 67658 270755
rect 191926 270703 191978 270755
rect 81814 270629 81866 270681
rect 206230 270703 206282 270755
rect 215542 270703 215594 270755
rect 219286 271073 219338 271125
rect 234646 271073 234698 271125
rect 264502 271073 264554 271125
rect 278518 271073 278570 271125
rect 315670 271073 315722 271125
rect 324598 271073 324650 271125
rect 324694 271073 324746 271125
rect 325654 271073 325706 271125
rect 326326 271073 326378 271125
rect 341494 271073 341546 271125
rect 345238 271073 345290 271125
rect 354838 271073 354890 271125
rect 355222 271147 355274 271199
rect 370006 271147 370058 271199
rect 370198 271221 370250 271273
rect 389398 271221 389450 271273
rect 390454 271221 390506 271273
rect 394390 271221 394442 271273
rect 394486 271221 394538 271273
rect 511894 271221 511946 271273
rect 383158 271147 383210 271199
rect 385462 271147 385514 271199
rect 389302 271147 389354 271199
rect 358390 271073 358442 271125
rect 358486 271073 358538 271125
rect 365014 271073 365066 271125
rect 367030 271073 367082 271125
rect 371926 271073 371978 271125
rect 372886 271073 372938 271125
rect 398038 271147 398090 271199
rect 398230 271147 398282 271199
rect 483286 271147 483338 271199
rect 218902 270999 218954 271051
rect 231190 270999 231242 271051
rect 253750 270999 253802 271051
rect 277270 270999 277322 271051
rect 282166 270999 282218 271051
rect 293014 270999 293066 271051
rect 300214 270999 300266 271051
rect 317974 270999 318026 271051
rect 320374 270999 320426 271051
rect 325366 270999 325418 271051
rect 325558 270999 325610 271051
rect 341302 270999 341354 271051
rect 344758 270999 344810 271051
rect 350998 270999 351050 271051
rect 218710 270925 218762 270977
rect 227638 270925 227690 270977
rect 268726 270925 268778 270977
rect 270550 270925 270602 270977
rect 281686 270925 281738 270977
rect 289462 270925 289514 270977
rect 313846 270925 313898 270977
rect 320470 270925 320522 270977
rect 320566 270925 320618 270977
rect 327958 270925 328010 270977
rect 328054 270925 328106 270977
rect 340438 270925 340490 270977
rect 346390 270925 346442 270977
rect 349558 270925 349610 270977
rect 349654 270925 349706 270977
rect 362998 270999 363050 271051
rect 363094 270999 363146 271051
rect 377974 270999 378026 271051
rect 378070 270999 378122 271051
rect 358486 270925 358538 270977
rect 378934 270999 378986 271051
rect 379414 270999 379466 271051
rect 379510 270999 379562 271051
rect 379798 270999 379850 271051
rect 379894 270999 379946 271051
rect 380086 270999 380138 271051
rect 380278 270999 380330 271051
rect 380950 270999 381002 271051
rect 381430 270999 381482 271051
rect 388918 270999 388970 271051
rect 221014 270851 221066 270903
rect 249046 270851 249098 270903
rect 253462 270851 253514 270903
rect 259702 270851 259754 270903
rect 260950 270851 261002 270903
rect 277942 270851 277994 270903
rect 279958 270851 280010 270903
rect 284854 270851 284906 270903
rect 296758 270851 296810 270903
rect 381142 270925 381194 270977
rect 381238 270925 381290 270977
rect 390646 271073 390698 271125
rect 409558 271073 409610 271125
rect 410422 271073 410474 271125
rect 416662 271073 416714 271125
rect 398806 270999 398858 271051
rect 516598 270999 516650 271051
rect 527350 270925 527402 270977
rect 257302 270777 257354 270829
rect 277462 270777 277514 270829
rect 317206 270777 317258 270829
rect 327094 270777 327146 270829
rect 327190 270777 327242 270829
rect 372886 270777 372938 270829
rect 372982 270777 373034 270829
rect 377782 270777 377834 270829
rect 382006 270851 382058 270903
rect 383158 270851 383210 270903
rect 383638 270851 383690 270903
rect 385942 270851 385994 270903
rect 390454 270851 390506 270903
rect 390550 270851 390602 270903
rect 406678 270851 406730 270903
rect 406774 270851 406826 270903
rect 543958 270851 544010 270903
rect 392086 270777 392138 270829
rect 394390 270777 394442 270829
rect 402454 270777 402506 270829
rect 402550 270777 402602 270829
rect 536854 270777 536906 270829
rect 358486 270703 358538 270755
rect 364150 270703 364202 270755
rect 369046 270703 369098 270755
rect 207190 270629 207242 270681
rect 231286 270629 231338 270681
rect 328150 270629 328202 270681
rect 328246 270629 328298 270681
rect 338902 270629 338954 270681
rect 341974 270629 342026 270681
rect 373462 270703 373514 270755
rect 374998 270703 375050 270755
rect 369238 270629 369290 270681
rect 380374 270629 380426 270681
rect 381238 270703 381290 270755
rect 383350 270703 383402 270755
rect 383638 270703 383690 270755
rect 387766 270703 387818 270755
rect 389014 270703 389066 270755
rect 411478 270703 411530 270755
rect 414838 270703 414890 270755
rect 434806 270703 434858 270755
rect 385942 270629 385994 270681
rect 386038 270629 386090 270681
rect 565462 270629 565514 270681
rect 245302 270555 245354 270607
rect 445270 270555 445322 270607
rect 231958 270481 232010 270533
rect 328342 270481 328394 270533
rect 331222 270481 331274 270533
rect 338230 270481 338282 270533
rect 338326 270481 338378 270533
rect 348214 270481 348266 270533
rect 348406 270481 348458 270533
rect 362710 270481 362762 270533
rect 365206 270481 365258 270533
rect 368470 270481 368522 270533
rect 245878 270407 245930 270459
rect 368566 270407 368618 270459
rect 232822 270333 232874 270385
rect 328342 270333 328394 270385
rect 328438 270333 328490 270385
rect 334102 270333 334154 270385
rect 233974 270259 234026 270311
rect 352438 270333 352490 270385
rect 353302 270333 353354 270385
rect 378550 270481 378602 270533
rect 378646 270481 378698 270533
rect 394486 270481 394538 270533
rect 394582 270481 394634 270533
rect 403126 270481 403178 270533
rect 427606 270481 427658 270533
rect 437686 270481 437738 270533
rect 368854 270407 368906 270459
rect 452374 270407 452426 270459
rect 552982 270407 553034 270459
rect 573046 270407 573098 270459
rect 590422 270407 590474 270459
rect 600502 270407 600554 270459
rect 336598 270259 336650 270311
rect 343126 270259 343178 270311
rect 359446 270259 359498 270311
rect 388438 270333 388490 270385
rect 388534 270333 388586 270385
rect 579670 270333 579722 270385
rect 369046 270259 369098 270311
rect 383638 270259 383690 270311
rect 383926 270259 383978 270311
rect 586774 270259 586826 270311
rect 247030 270185 247082 270237
rect 348310 270185 348362 270237
rect 234550 270111 234602 270163
rect 323158 270111 323210 270163
rect 323350 270111 323402 270163
rect 336886 270111 336938 270163
rect 235702 270037 235754 270089
rect 342166 270111 342218 270163
rect 341878 270037 341930 270089
rect 348118 270037 348170 270089
rect 348310 270037 348362 270089
rect 459574 270185 459626 270237
rect 355414 270111 355466 270163
rect 364150 270111 364202 270163
rect 364342 270111 364394 270163
rect 378166 270111 378218 270163
rect 355606 270037 355658 270089
rect 370006 270037 370058 270089
rect 370198 270037 370250 270089
rect 374998 270037 375050 270089
rect 375094 270037 375146 270089
rect 380278 270111 380330 270163
rect 380374 270111 380426 270163
rect 381046 270111 381098 270163
rect 381142 270111 381194 270163
rect 593974 270111 594026 270163
rect 378550 270037 378602 270089
rect 380086 270037 380138 270089
rect 380470 270037 380522 270089
rect 380854 270037 380906 270089
rect 380950 270037 381002 270089
rect 427606 270037 427658 270089
rect 159862 269963 159914 270015
rect 161110 269963 161162 270015
rect 247606 269963 247658 270015
rect 437686 270037 437738 270089
rect 597526 270037 597578 270089
rect 466582 269963 466634 270015
rect 573142 269963 573194 270015
rect 589174 269963 589226 270015
rect 216022 269889 216074 269941
rect 243286 269889 243338 269941
rect 248566 269889 248618 269941
rect 226966 269815 227018 269867
rect 295414 269815 295466 269867
rect 295510 269815 295562 269867
rect 302518 269815 302570 269867
rect 308182 269815 308234 269867
rect 311926 269815 311978 269867
rect 312022 269815 312074 269867
rect 316342 269815 316394 269867
rect 316438 269815 316490 269867
rect 327862 269815 327914 269867
rect 327958 269815 328010 269867
rect 338326 269815 338378 269867
rect 342166 269815 342218 269867
rect 427606 269889 427658 269941
rect 437590 269889 437642 269941
rect 473782 269889 473834 269941
rect 348214 269815 348266 269867
rect 437110 269815 437162 269867
rect 437494 269815 437546 269867
rect 539254 269815 539306 269867
rect 249622 269741 249674 269793
rect 250294 269667 250346 269719
rect 341878 269667 341930 269719
rect 342550 269741 342602 269793
rect 481078 269741 481130 269793
rect 483958 269741 484010 269793
rect 518326 269741 518378 269793
rect 348118 269667 348170 269719
rect 365206 269667 365258 269719
rect 365302 269667 365354 269719
rect 379702 269667 379754 269719
rect 379798 269667 379850 269719
rect 437974 269667 438026 269719
rect 438166 269667 438218 269719
rect 488086 269667 488138 269719
rect 251350 269593 251402 269645
rect 336214 269593 336266 269645
rect 342838 269593 342890 269645
rect 437398 269593 437450 269645
rect 437590 269593 437642 269645
rect 437782 269593 437834 269645
rect 437878 269593 437930 269645
rect 495190 269593 495242 269645
rect 85270 269519 85322 269571
rect 86518 269519 86570 269571
rect 227542 269519 227594 269571
rect 295510 269519 295562 269571
rect 297910 269519 297962 269571
rect 308182 269519 308234 269571
rect 308278 269519 308330 269571
rect 316822 269519 316874 269571
rect 318166 269519 318218 269571
rect 326806 269519 326858 269571
rect 328054 269519 328106 269571
rect 236278 269445 236330 269497
rect 341974 269445 342026 269497
rect 417718 269519 417770 269571
rect 437686 269519 437738 269571
rect 458230 269519 458282 269571
rect 478006 269519 478058 269571
rect 501046 269519 501098 269571
rect 501142 269519 501194 269571
rect 509878 269593 509930 269645
rect 529846 269519 529898 269571
rect 560662 269519 560714 269571
rect 573142 269519 573194 269571
rect 593206 269519 593258 269571
rect 360982 269445 361034 269497
rect 378550 269445 378602 269497
rect 378646 269445 378698 269497
rect 393142 269445 393194 269497
rect 398806 269445 398858 269497
rect 437494 269445 437546 269497
rect 437590 269445 437642 269497
rect 457942 269445 457994 269497
rect 458614 269445 458666 269497
rect 532822 269445 532874 269497
rect 533110 269445 533162 269497
rect 626038 269445 626090 269497
rect 228502 269371 228554 269423
rect 229558 269297 229610 269349
rect 297910 269297 297962 269349
rect 304918 269371 304970 269423
rect 327958 269371 328010 269423
rect 328438 269371 328490 269423
rect 437302 269371 437354 269423
rect 437398 269371 437450 269423
rect 437782 269371 437834 269423
rect 309718 269297 309770 269349
rect 311926 269297 311978 269349
rect 316054 269297 316106 269349
rect 316150 269297 316202 269349
rect 327574 269297 327626 269349
rect 327862 269297 327914 269349
rect 438262 269371 438314 269423
rect 567766 269371 567818 269423
rect 53878 269223 53930 269275
rect 205942 269223 205994 269275
rect 221494 269223 221546 269275
rect 252502 269223 252554 269275
rect 254134 269223 254186 269275
rect 342070 269223 342122 269275
rect 342454 269223 342506 269275
rect 380182 269223 380234 269275
rect 244150 269149 244202 269201
rect 341974 269149 342026 269201
rect 342550 269149 342602 269201
rect 381622 269223 381674 269275
rect 574870 269297 574922 269349
rect 467926 269223 467978 269275
rect 520150 269223 520202 269275
rect 632086 269223 632138 269275
rect 649366 269223 649418 269275
rect 203830 269075 203882 269127
rect 270934 269075 270986 269127
rect 272758 269075 272810 269127
rect 316150 269075 316202 269127
rect 316246 269075 316298 269127
rect 336118 269075 336170 269127
rect 336214 269075 336266 269127
rect 342646 269075 342698 269127
rect 342742 269075 342794 269127
rect 366742 269075 366794 269127
rect 367318 269075 367370 269127
rect 378646 269075 378698 269127
rect 378742 269075 378794 269127
rect 438358 269149 438410 269201
rect 457942 269149 457994 269201
rect 509878 269149 509930 269201
rect 529846 269149 529898 269201
rect 243286 269001 243338 269053
rect 558262 269075 558314 269127
rect 242614 268927 242666 268979
rect 431062 269001 431114 269053
rect 458038 269001 458090 269053
rect 467926 269001 467978 269053
rect 237142 268853 237194 268905
rect 355414 268853 355466 268905
rect 355510 268853 355562 268905
rect 360886 268853 360938 268905
rect 362710 268853 362762 268905
rect 377590 268853 377642 268905
rect 378358 268853 378410 268905
rect 423862 268927 423914 268979
rect 458518 268927 458570 268979
rect 478006 268927 478058 268979
rect 398806 268853 398858 268905
rect 417718 268853 417770 268905
rect 437686 268853 437738 268905
rect 241558 268779 241610 268831
rect 380182 268779 380234 268831
rect 240886 268705 240938 268757
rect 380854 268779 380906 268831
rect 238294 268631 238346 268683
rect 379894 268631 379946 268683
rect 380182 268631 380234 268683
rect 380854 268631 380906 268683
rect 390646 268705 390698 268757
rect 410422 268779 410474 268831
rect 381238 268631 381290 268683
rect 483958 268853 484010 268905
rect 483862 268779 483914 268831
rect 560086 268779 560138 268831
rect 238870 268557 238922 268609
rect 368662 268557 368714 268609
rect 240022 268483 240074 268535
rect 370198 268557 370250 268609
rect 370294 268557 370346 268609
rect 378742 268557 378794 268609
rect 378838 268557 378890 268609
rect 380278 268557 380330 268609
rect 380566 268557 380618 268609
rect 388534 268557 388586 268609
rect 388822 268557 388874 268609
rect 389398 268557 389450 268609
rect 389494 268557 389546 268609
rect 400726 268557 400778 268609
rect 368854 268483 368906 268535
rect 387670 268483 387722 268535
rect 387766 268483 387818 268535
rect 397366 268483 397418 268535
rect 225814 268409 225866 268461
rect 288214 268409 288266 268461
rect 294262 268409 294314 268461
rect 210934 268335 210986 268387
rect 271990 268335 272042 268387
rect 284854 268335 284906 268387
rect 316246 268335 316298 268387
rect 321910 268409 321962 268461
rect 324598 268409 324650 268461
rect 324694 268409 324746 268461
rect 338038 268409 338090 268461
rect 357046 268409 357098 268461
rect 451126 268409 451178 268461
rect 337846 268335 337898 268387
rect 357622 268335 357674 268387
rect 218038 268261 218090 268313
rect 272662 268261 272714 268313
rect 287062 268261 287114 268313
rect 312022 268261 312074 268313
rect 312214 268261 312266 268313
rect 330070 268261 330122 268313
rect 333430 268261 333482 268313
rect 342646 268261 342698 268313
rect 355414 268261 355466 268313
rect 360118 268261 360170 268313
rect 223702 268187 223754 268239
rect 270358 268187 270410 268239
rect 285046 268187 285098 268239
rect 312886 268187 312938 268239
rect 314806 268187 314858 268239
rect 322486 268187 322538 268239
rect 322774 268187 322826 268239
rect 326710 268187 326762 268239
rect 326806 268187 326858 268239
rect 355606 268187 355658 268239
rect 355894 268187 355946 268239
rect 360214 268187 360266 268239
rect 360886 268335 360938 268387
rect 436918 268335 436970 268387
rect 360406 268261 360458 268313
rect 380374 268261 380426 268313
rect 380470 268261 380522 268313
rect 419062 268261 419114 268313
rect 377110 268187 377162 268239
rect 378646 268187 378698 268239
rect 223222 268113 223274 268165
rect 266518 268113 266570 268165
rect 286006 268113 286058 268165
rect 315766 268113 315818 268165
rect 315862 268113 315914 268165
rect 317878 268113 317930 268165
rect 235894 268039 235946 268091
rect 222550 267965 222602 268017
rect 253462 267965 253514 268017
rect 274870 268039 274922 268091
rect 310966 268039 311018 268091
rect 317686 268039 317738 268091
rect 322198 268113 322250 268165
rect 322294 268113 322346 268165
rect 328054 268113 328106 268165
rect 328246 268113 328298 268165
rect 334966 268113 335018 268165
rect 243094 267891 243146 267943
rect 275734 267965 275786 268017
rect 296662 267965 296714 268017
rect 308278 267965 308330 268017
rect 312598 267965 312650 268017
rect 321430 268039 321482 268091
rect 326614 268039 326666 268091
rect 326710 268039 326762 268091
rect 347158 268039 347210 268091
rect 355894 268039 355946 268091
rect 357430 268113 357482 268165
rect 369238 268113 369290 268165
rect 371830 268113 371882 268165
rect 388246 268113 388298 268165
rect 388438 268187 388490 268239
rect 411286 268187 411338 268239
rect 398230 268113 398282 268165
rect 371446 268039 371498 268091
rect 372694 268039 372746 268091
rect 317878 267965 317930 268017
rect 328438 267965 328490 268017
rect 328534 267965 328586 268017
rect 345334 267965 345386 268017
rect 349846 267965 349898 268017
rect 266614 267891 266666 267943
rect 355414 267891 355466 267943
rect 358678 267965 358730 268017
rect 368854 267965 368906 268017
rect 368950 267965 369002 268017
rect 374230 267965 374282 268017
rect 374710 267965 374762 268017
rect 378838 267965 378890 268017
rect 379222 267965 379274 268017
rect 385366 267965 385418 268017
rect 368758 267891 368810 267943
rect 370966 267891 371018 267943
rect 376630 267891 376682 267943
rect 377206 267891 377258 267943
rect 380278 267891 380330 267943
rect 380374 267891 380426 267943
rect 382966 267891 383018 267943
rect 383062 267891 383114 267943
rect 388150 267891 388202 267943
rect 388918 268039 388970 268091
rect 572470 268039 572522 268091
rect 389014 267965 389066 268017
rect 397558 267965 397610 268017
rect 393814 267891 393866 267943
rect 393910 267891 393962 267943
rect 399382 267891 399434 267943
rect 65014 267817 65066 267869
rect 221974 267817 222026 267869
rect 256150 267817 256202 267869
rect 267670 267817 267722 267869
rect 357334 267817 357386 267869
rect 359062 267817 359114 267869
rect 388822 267817 388874 267869
rect 389110 267817 389162 267869
rect 401110 267817 401162 267869
rect 77782 267743 77834 267795
rect 290614 267743 290666 267795
rect 315094 267743 315146 267795
rect 315190 267743 315242 267795
rect 322294 267743 322346 267795
rect 322390 267743 322442 267795
rect 326326 267743 326378 267795
rect 326422 267743 326474 267795
rect 327574 267743 327626 267795
rect 328054 267743 328106 267795
rect 329302 267743 329354 267795
rect 329398 267743 329450 267795
rect 332566 267743 332618 267795
rect 336886 267743 336938 267795
rect 628438 267743 628490 267795
rect 255670 267669 255722 267721
rect 267766 267669 267818 267721
rect 298102 267669 298154 267721
rect 317014 267669 317066 267721
rect 317302 267669 317354 267721
rect 318454 267669 318506 267721
rect 318550 267669 318602 267721
rect 289462 267595 289514 267647
rect 267862 267521 267914 267573
rect 287926 267521 287978 267573
rect 290326 267521 290378 267573
rect 300022 267521 300074 267573
rect 300406 267595 300458 267647
rect 328726 267595 328778 267647
rect 328918 267669 328970 267721
rect 349846 267669 349898 267721
rect 352246 267669 352298 267721
rect 356854 267669 356906 267721
rect 356950 267669 357002 267721
rect 366742 267669 366794 267721
rect 366838 267669 366890 267721
rect 369334 267669 369386 267721
rect 330646 267595 330698 267647
rect 332566 267595 332618 267647
rect 337654 267595 337706 267647
rect 353686 267595 353738 267647
rect 354262 267595 354314 267647
rect 366646 267595 366698 267647
rect 366934 267595 366986 267647
rect 372886 267595 372938 267647
rect 377206 267595 377258 267647
rect 377494 267669 377546 267721
rect 379990 267669 380042 267721
rect 380086 267669 380138 267721
rect 383062 267669 383114 267721
rect 265750 267447 265802 267499
rect 317206 267447 317258 267499
rect 317686 267447 317738 267499
rect 327766 267447 327818 267499
rect 291478 267373 291530 267425
rect 299926 267373 299978 267425
rect 300022 267373 300074 267425
rect 327958 267373 328010 267425
rect 258838 267299 258890 267351
rect 321430 267299 321482 267351
rect 321526 267299 321578 267351
rect 337462 267447 337514 267499
rect 347158 267521 347210 267573
rect 347830 267521 347882 267573
rect 348982 267521 349034 267573
rect 328342 267373 328394 267425
rect 338806 267447 338858 267499
rect 348502 267447 348554 267499
rect 337942 267373 337994 267425
rect 343702 267373 343754 267425
rect 348214 267373 348266 267425
rect 349846 267447 349898 267499
rect 350710 267447 350762 267499
rect 356950 267521 357002 267573
rect 361558 267521 361610 267573
rect 377110 267521 377162 267573
rect 378742 267595 378794 267647
rect 515446 267669 515498 267721
rect 391990 267595 392042 267647
rect 396598 267595 396650 267647
rect 397174 267595 397226 267647
rect 397270 267595 397322 267647
rect 411862 267595 411914 267647
rect 384214 267521 384266 267573
rect 356854 267447 356906 267499
rect 348694 267373 348746 267425
rect 366454 267373 366506 267425
rect 328246 267299 328298 267351
rect 347830 267299 347882 267351
rect 348502 267299 348554 267351
rect 358678 267299 358730 267351
rect 267574 267225 267626 267277
rect 268054 267225 268106 267277
rect 292534 267225 292586 267277
rect 299830 267225 299882 267277
rect 299926 267225 299978 267277
rect 348694 267225 348746 267277
rect 251638 267151 251690 267203
rect 315190 267151 315242 267203
rect 317110 267151 317162 267203
rect 317782 267151 317834 267203
rect 293590 267077 293642 267129
rect 299734 267077 299786 267129
rect 299830 267077 299882 267129
rect 318166 267151 318218 267203
rect 328246 267151 328298 267203
rect 328438 267151 328490 267203
rect 337942 267151 337994 267203
rect 338038 267151 338090 267203
rect 348214 267151 348266 267203
rect 348598 267151 348650 267203
rect 359062 267225 359114 267277
rect 359158 267225 359210 267277
rect 366646 267447 366698 267499
rect 367894 267447 367946 267499
rect 368182 267447 368234 267499
rect 397750 267447 397802 267499
rect 397942 267521 397994 267573
rect 408790 267521 408842 267573
rect 406006 267447 406058 267499
rect 367414 267373 367466 267425
rect 366742 267299 366794 267351
rect 368182 267299 368234 267351
rect 368470 267299 368522 267351
rect 377398 267299 377450 267351
rect 377590 267373 377642 267425
rect 378550 267299 378602 267351
rect 378934 267373 378986 267425
rect 392950 267373 393002 267425
rect 387766 267299 387818 267351
rect 388822 267299 388874 267351
rect 399574 267373 399626 267425
rect 408982 267373 409034 267425
rect 426262 267373 426314 267425
rect 396790 267299 396842 267351
rect 413782 267299 413834 267351
rect 348982 267151 349034 267203
rect 354262 267151 354314 267203
rect 355030 267151 355082 267203
rect 366166 267151 366218 267203
rect 244246 267003 244298 267055
rect 317302 267003 317354 267055
rect 317974 267003 318026 267055
rect 326230 267003 326282 267055
rect 326326 267003 326378 267055
rect 237430 266929 237482 266981
rect 318358 266929 318410 266981
rect 318454 266929 318506 266981
rect 318838 266929 318890 266981
rect 318934 266929 318986 266981
rect 327382 266929 327434 266981
rect 327574 267003 327626 267055
rect 327958 267003 328010 267055
rect 328246 267003 328298 267055
rect 329014 267077 329066 267129
rect 331894 267077 331946 267129
rect 328342 266929 328394 266981
rect 337174 267003 337226 267055
rect 366358 267077 366410 267129
rect 367990 267225 368042 267277
rect 368374 267225 368426 267277
rect 368758 267225 368810 267277
rect 369046 267225 369098 267277
rect 374422 267225 374474 267277
rect 374230 267151 374282 267203
rect 374806 267225 374858 267277
rect 377110 267225 377162 267277
rect 409078 267225 409130 267277
rect 367894 267077 367946 267129
rect 374422 267077 374474 267129
rect 374806 267077 374858 267129
rect 377494 267077 377546 267129
rect 377686 267077 377738 267129
rect 386230 267077 386282 267129
rect 389014 267151 389066 267203
rect 412534 267151 412586 267203
rect 393046 267077 393098 267129
rect 398326 267077 398378 267129
rect 421462 267077 421514 267129
rect 329974 266929 330026 266981
rect 330070 266929 330122 266981
rect 337366 266929 337418 266981
rect 337462 266929 337514 266981
rect 348022 266929 348074 266981
rect 349846 267003 349898 267055
rect 366262 267003 366314 267055
rect 349366 266929 349418 266981
rect 353974 266929 354026 266981
rect 366550 266929 366602 266981
rect 367606 266929 367658 266981
rect 367990 267003 368042 267055
rect 397270 267003 397322 267055
rect 399286 267003 399338 267055
rect 408886 267003 408938 267055
rect 408982 266929 409034 266981
rect 293782 266855 293834 266907
rect 294262 266781 294314 266833
rect 299734 266855 299786 266907
rect 377878 266855 377930 266907
rect 377974 266855 378026 266907
rect 384214 266855 384266 266907
rect 287638 266707 287690 266759
rect 296662 266707 296714 266759
rect 369142 266781 369194 266833
rect 369334 266781 369386 266833
rect 378742 266707 378794 266759
rect 379030 266781 379082 266833
rect 385462 266781 385514 266833
rect 391030 266855 391082 266907
rect 393046 266855 393098 266907
rect 404470 266855 404522 266907
rect 406102 266855 406154 266907
rect 407158 266855 407210 266907
rect 408502 266855 408554 266907
rect 413398 266929 413450 266981
rect 397750 266781 397802 266833
rect 403222 266781 403274 266833
rect 408598 266781 408650 266833
rect 413686 266781 413738 266833
rect 230038 266633 230090 266685
rect 318166 266633 318218 266685
rect 318550 266633 318602 266685
rect 326422 266633 326474 266685
rect 326518 266633 326570 266685
rect 328054 266633 328106 266685
rect 295318 266559 295370 266611
rect 328246 266559 328298 266611
rect 215734 266485 215786 266537
rect 309814 266485 309866 266537
rect 310006 266485 310058 266537
rect 312982 266485 313034 266537
rect 315094 266485 315146 266537
rect 337270 266633 337322 266685
rect 337654 266633 337706 266685
rect 367414 266633 367466 266685
rect 367606 266633 367658 266685
rect 389590 266707 389642 266759
rect 393046 266707 393098 266759
rect 407350 266707 407402 266759
rect 408694 266707 408746 266759
rect 409654 266707 409706 266759
rect 389782 266633 389834 266685
rect 433366 266633 433418 266685
rect 328918 266559 328970 266611
rect 377686 266559 377738 266611
rect 377878 266559 377930 266611
rect 378454 266559 378506 266611
rect 378550 266559 378602 266611
rect 393046 266559 393098 266611
rect 406870 266559 406922 266611
rect 407734 266559 407786 266611
rect 409078 266559 409130 266611
rect 410326 266559 410378 266611
rect 328534 266485 328586 266537
rect 338806 266485 338858 266537
rect 347830 266485 347882 266537
rect 348598 266485 348650 266537
rect 349078 266485 349130 266537
rect 357526 266485 357578 266537
rect 358294 266485 358346 266537
rect 367414 266485 367466 266537
rect 367606 266485 367658 266537
rect 447670 266485 447722 266537
rect 270646 266411 270698 266463
rect 287926 266411 287978 266463
rect 295990 266411 296042 266463
rect 389398 266411 389450 266463
rect 399094 266411 399146 266463
rect 400246 266411 400298 266463
rect 400726 266411 400778 266463
rect 406102 266411 406154 266463
rect 406582 266411 406634 266463
rect 408598 266411 408650 266463
rect 287638 266337 287690 266389
rect 296758 266337 296810 266389
rect 296854 266337 296906 266389
rect 208534 266263 208586 266315
rect 310006 266263 310058 266315
rect 310102 266263 310154 266315
rect 317110 266263 317162 266315
rect 317206 266263 317258 266315
rect 317590 266263 317642 266315
rect 317974 266263 318026 266315
rect 318262 266263 318314 266315
rect 298006 266189 298058 266241
rect 318166 266189 318218 266241
rect 201430 266115 201482 266167
rect 310102 266115 310154 266167
rect 310198 266115 310250 266167
rect 312886 266115 312938 266167
rect 312982 266115 313034 266167
rect 318934 266263 318986 266315
rect 322486 266263 322538 266315
rect 328630 266263 328682 266315
rect 328822 266263 328874 266315
rect 346582 266263 346634 266315
rect 348022 266263 348074 266315
rect 349846 266263 349898 266315
rect 349942 266263 349994 266315
rect 357814 266263 357866 266315
rect 366454 266263 366506 266315
rect 367318 266263 367370 266315
rect 367414 266263 367466 266315
rect 393910 266263 393962 266315
rect 318454 266189 318506 266241
rect 398326 266189 398378 266241
rect 399574 266337 399626 266389
rect 413206 266337 413258 266389
rect 501622 266337 501674 266389
rect 569878 266337 569930 266389
rect 399382 266263 399434 266315
rect 461974 266263 462026 266315
rect 414358 266189 414410 266241
rect 318838 266115 318890 266167
rect 331702 266115 331754 266167
rect 331894 266115 331946 266167
rect 349942 266115 349994 266167
rect 351286 266115 351338 266167
rect 359158 266115 359210 266167
rect 360022 266115 360074 266167
rect 476182 266115 476234 266167
rect 298582 266041 298634 266093
rect 428662 266041 428714 266093
rect 299734 265967 299786 266019
rect 435670 265967 435722 266019
rect 300310 265893 300362 265945
rect 442870 265893 442922 265945
rect 288790 265819 288842 265871
rect 300406 265819 300458 265871
rect 301270 265819 301322 265871
rect 449974 265819 450026 265871
rect 287254 265745 287306 265797
rect 298102 265745 298154 265797
rect 302326 265745 302378 265797
rect 457174 265745 457226 265797
rect 302998 265671 303050 265723
rect 312214 265671 312266 265723
rect 312886 265671 312938 265723
rect 337174 265671 337226 265723
rect 337558 265671 337610 265723
rect 464278 265671 464330 265723
rect 304054 265597 304106 265649
rect 471382 265597 471434 265649
rect 257590 265523 257642 265575
rect 269878 265523 269930 265575
rect 304726 265523 304778 265575
rect 478582 265523 478634 265575
rect 306742 265449 306794 265501
rect 492886 265449 492938 265501
rect 307318 265375 307370 265427
rect 499894 265375 499946 265427
rect 308230 265301 308282 265353
rect 507094 265301 507146 265353
rect 225334 265227 225386 265279
rect 273622 265227 273674 265279
rect 308854 265227 308906 265279
rect 510646 265227 510698 265279
rect 221686 265153 221738 265205
rect 273142 265153 273194 265205
rect 309334 265153 309386 265205
rect 514294 265153 514346 265205
rect 223126 265079 223178 265131
rect 329014 265079 329066 265131
rect 329686 265079 329738 265131
rect 332374 265079 332426 265131
rect 349846 265079 349898 265131
rect 372982 265079 373034 265131
rect 376918 265079 376970 265131
rect 611830 265079 611882 265131
rect 197878 265005 197930 265057
rect 325846 265005 325898 265057
rect 326614 265005 326666 265057
rect 333142 265005 333194 265057
rect 356854 265005 356906 265057
rect 367606 265005 367658 265057
rect 81814 264931 81866 264983
rect 90646 264931 90698 264983
rect 309814 264931 309866 264983
rect 318358 264931 318410 264983
rect 318454 264931 318506 264983
rect 318742 264931 318794 264983
rect 324118 264931 324170 264983
rect 329302 264931 329354 264983
rect 347734 264931 347786 264983
rect 368566 265005 368618 265057
rect 369142 265005 369194 265057
rect 378646 265005 378698 265057
rect 379510 265005 379562 265057
rect 633142 265005 633194 265057
rect 369526 264931 369578 264983
rect 343702 264857 343754 264909
rect 382390 264857 382442 264909
rect 388630 264931 388682 264983
rect 413206 264931 413258 264983
rect 455158 264931 455210 264983
rect 475126 264931 475178 264983
rect 483862 264931 483914 264983
rect 511126 264931 511178 264983
rect 551062 264857 551114 264909
rect 158614 264487 158666 264539
rect 161206 264487 161258 264539
rect 42262 264265 42314 264317
rect 50518 264265 50570 264317
rect 77782 263599 77834 263651
rect 87766 263599 87818 263651
rect 42646 263229 42698 263281
rect 53398 263229 53450 263281
rect 42646 262267 42698 262319
rect 56182 262267 56234 262319
rect 87766 260713 87818 260765
rect 93334 260713 93386 260765
rect 90646 260639 90698 260691
rect 102550 260639 102602 260691
rect 639286 256347 639338 256399
rect 679798 256347 679850 256399
rect 93334 256273 93386 256325
rect 97846 256273 97898 256325
rect 44566 255089 44618 255141
rect 60406 255089 60458 255141
rect 625174 253387 625226 253439
rect 632086 253461 632138 253513
rect 100150 252943 100202 252995
rect 100726 252943 100778 252995
rect 191446 252425 191498 252477
rect 193270 252425 193322 252477
rect 53782 252055 53834 252107
rect 210646 252055 210698 252107
rect 45046 251981 45098 252033
rect 206806 251981 206858 252033
rect 497494 251611 497546 251663
rect 501622 251611 501674 251663
rect 674998 251611 675050 251663
rect 676918 251611 676970 251663
rect 675094 251537 675146 251589
rect 676822 251537 676874 251589
rect 674518 250945 674570 250997
rect 675382 250945 675434 250997
rect 674614 250353 674666 250405
rect 675478 250353 675530 250405
rect 42166 249835 42218 249887
rect 42646 249835 42698 249887
rect 674134 249539 674186 249591
rect 675382 249539 675434 249591
rect 613462 249095 613514 249147
rect 625174 249095 625226 249147
rect 673942 247911 673994 247963
rect 675382 247911 675434 247963
rect 205846 247393 205898 247445
rect 211606 247319 211658 247371
rect 211798 247245 211850 247297
rect 212182 247171 212234 247223
rect 211990 247097 212042 247149
rect 90742 246949 90794 247001
rect 100246 246949 100298 247001
rect 187894 246949 187946 247001
rect 201526 246949 201578 247001
rect 63286 246875 63338 246927
rect 204982 246875 205034 246927
rect 56086 246801 56138 246853
rect 204694 246801 204746 246853
rect 211606 246801 211658 246853
rect 53494 246727 53546 246779
rect 204790 246727 204842 246779
rect 56278 246653 56330 246705
rect 210166 246653 210218 246705
rect 53686 246579 53738 246631
rect 90742 246579 90794 246631
rect 100246 246579 100298 246631
rect 212662 246727 212714 246779
rect 221590 246727 221642 246779
rect 228214 246727 228266 246779
rect 229654 246727 229706 246779
rect 243094 246727 243146 246779
rect 246166 246727 246218 246779
rect 254038 246727 254090 246779
rect 211126 246653 211178 246705
rect 211030 246579 211082 246631
rect 226006 246579 226058 246631
rect 226390 246653 226442 246705
rect 243382 246653 243434 246705
rect 248278 246653 248330 246705
rect 266614 246653 266666 246705
rect 267478 246727 267530 246779
rect 269302 246727 269354 246779
rect 288310 246727 288362 246779
rect 288406 246727 288458 246779
rect 290134 246727 290186 246779
rect 291094 246727 291146 246779
rect 292630 246727 292682 246779
rect 309718 246727 309770 246779
rect 309814 246727 309866 246779
rect 310006 246727 310058 246779
rect 311158 246727 311210 246779
rect 326326 246727 326378 246779
rect 290038 246653 290090 246705
rect 292150 246653 292202 246705
rect 297142 246653 297194 246705
rect 304630 246653 304682 246705
rect 247702 246579 247754 246631
rect 247798 246579 247850 246631
rect 53302 246505 53354 246557
rect 90646 246505 90698 246557
rect 100534 246505 100586 246557
rect 212278 246505 212330 246557
rect 221590 246505 221642 246557
rect 229654 246505 229706 246557
rect 229942 246505 229994 246557
rect 243190 246505 243242 246557
rect 53206 246431 53258 246483
rect 44662 246357 44714 246409
rect 100246 246357 100298 246409
rect 100630 246357 100682 246409
rect 204886 246357 204938 246409
rect 210550 246431 210602 246483
rect 228310 246431 228362 246483
rect 228694 246431 228746 246483
rect 267478 246505 267530 246557
rect 268822 246579 268874 246631
rect 280822 246579 280874 246631
rect 288406 246579 288458 246631
rect 290134 246579 290186 246631
rect 290998 246579 291050 246631
rect 291574 246579 291626 246631
rect 291958 246579 292010 246631
rect 328534 246653 328586 246705
rect 329014 246653 329066 246705
rect 339286 246653 339338 246705
rect 307990 246579 308042 246631
rect 309430 246579 309482 246631
rect 324022 246579 324074 246631
rect 348118 246727 348170 246779
rect 348598 246727 348650 246779
rect 348886 246727 348938 246779
rect 350326 246727 350378 246779
rect 339862 246579 339914 246631
rect 340150 246579 340202 246631
rect 350134 246579 350186 246631
rect 267862 246505 267914 246557
rect 269206 246505 269258 246557
rect 287830 246505 287882 246557
rect 287926 246505 287978 246557
rect 292630 246505 292682 246557
rect 297622 246505 297674 246557
rect 297910 246505 297962 246557
rect 300214 246505 300266 246557
rect 302326 246505 302378 246557
rect 307510 246505 307562 246557
rect 248182 246431 248234 246483
rect 44758 246283 44810 246335
rect 209686 246283 209738 246335
rect 60406 246209 60458 246261
rect 161302 246209 161354 246261
rect 181558 246209 181610 246261
rect 202582 246209 202634 246261
rect 210742 246357 210794 246409
rect 266518 246357 266570 246409
rect 266614 246357 266666 246409
rect 267766 246357 267818 246409
rect 267958 246431 268010 246483
rect 288022 246431 288074 246483
rect 288310 246431 288362 246483
rect 290614 246431 290666 246483
rect 308086 246505 308138 246557
rect 326326 246505 326378 246557
rect 328918 246505 328970 246557
rect 369814 246727 369866 246779
rect 369910 246727 369962 246779
rect 378646 246727 378698 246779
rect 389494 246727 389546 246779
rect 393046 246727 393098 246779
rect 393334 246727 393386 246779
rect 352342 246653 352394 246705
rect 377206 246653 377258 246705
rect 388246 246653 388298 246705
rect 389014 246653 389066 246705
rect 392566 246653 392618 246705
rect 393430 246653 393482 246705
rect 674038 247245 674090 247297
rect 675478 247245 675530 247297
rect 403318 246727 403370 246779
rect 674326 246727 674378 246779
rect 675382 246727 675434 246779
rect 368470 246579 368522 246631
rect 369046 246579 369098 246631
rect 369814 246579 369866 246631
rect 370678 246579 370730 246631
rect 388534 246579 388586 246631
rect 350614 246505 350666 246557
rect 369430 246505 369482 246557
rect 369718 246505 369770 246557
rect 389782 246505 389834 246557
rect 287926 246357 287978 246409
rect 288118 246357 288170 246409
rect 308086 246357 308138 246409
rect 310006 246431 310058 246483
rect 347542 246431 347594 246483
rect 350326 246431 350378 246483
rect 309622 246357 309674 246409
rect 309718 246357 309770 246409
rect 368374 246357 368426 246409
rect 389494 246431 389546 246483
rect 403798 246653 403850 246705
rect 404374 246505 404426 246557
rect 405142 246431 405194 246483
rect 378646 246357 378698 246409
rect 211318 246283 211370 246335
rect 228214 246283 228266 246335
rect 228310 246283 228362 246335
rect 229942 246283 229994 246335
rect 247702 246283 247754 246335
rect 324022 246283 324074 246335
rect 327094 246283 327146 246335
rect 211894 246209 211946 246261
rect 222454 246209 222506 246261
rect 269302 246209 269354 246261
rect 271606 246209 271658 246261
rect 287350 246209 287402 246261
rect 288118 246209 288170 246261
rect 307510 246209 307562 246261
rect 308182 246209 308234 246261
rect 161398 246135 161450 246187
rect 181462 246135 181514 246187
rect 226006 246135 226058 246187
rect 228694 246135 228746 246187
rect 243094 246135 243146 246187
rect 248278 246135 248330 246187
rect 263446 246135 263498 246187
rect 277942 246135 277994 246187
rect 280822 246135 280874 246187
rect 287830 246135 287882 246187
rect 288022 246135 288074 246187
rect 307894 246135 307946 246187
rect 309814 246209 309866 246261
rect 328918 246209 328970 246261
rect 339286 246283 339338 246335
rect 339862 246283 339914 246335
rect 339958 246283 340010 246335
rect 347254 246283 347306 246335
rect 350134 246283 350186 246335
rect 352342 246209 352394 246261
rect 367606 246283 367658 246335
rect 383350 246357 383402 246409
rect 383590 246357 383642 246409
rect 391990 246209 392042 246261
rect 393046 246209 393098 246261
rect 409174 246209 409226 246261
rect 340150 246135 340202 246187
rect 340246 246135 340298 246187
rect 347350 246135 347402 246187
rect 347542 246135 347594 246187
rect 350614 246135 350666 246187
rect 367990 246135 368042 246187
rect 370198 246135 370250 246187
rect 383062 246135 383114 246187
rect 383158 246135 383210 246187
rect 393334 246135 393386 246187
rect 403894 246135 403946 246187
rect 41302 246061 41354 246113
rect 43318 246061 43370 246113
rect 504022 246061 504074 246113
rect 43414 245987 43466 246039
rect 243190 245913 243242 245965
rect 248182 245913 248234 245965
rect 263830 245913 263882 245965
rect 181366 245839 181418 245891
rect 246166 245839 246218 245891
rect 248374 245839 248426 245891
rect 263062 245839 263114 245891
rect 277750 245839 277802 245891
rect 277942 245913 277994 245965
rect 339862 245913 339914 245965
rect 347350 245987 347402 246039
rect 509782 245987 509834 246039
rect 340246 245913 340298 245965
rect 347254 245913 347306 245965
rect 368086 245913 368138 245965
rect 368374 245913 368426 245965
rect 369718 245913 369770 245965
rect 391990 245913 392042 245965
rect 400918 245913 400970 245965
rect 367510 245839 367562 245891
rect 383158 245839 383210 245891
rect 401494 245839 401546 245891
rect 251830 245765 251882 245817
rect 356662 245765 356714 245817
rect 368566 245765 368618 245817
rect 388726 245765 388778 245817
rect 202582 245691 202634 245743
rect 213142 245691 213194 245743
rect 216886 245691 216938 245743
rect 228214 245691 228266 245743
rect 243382 245691 243434 245743
rect 254038 245691 254090 245743
rect 254134 245691 254186 245743
rect 358006 245691 358058 245743
rect 383062 245691 383114 245743
rect 392950 245691 393002 245743
rect 266518 245617 266570 245669
rect 269206 245617 269258 245669
rect 277750 245617 277802 245669
rect 369238 245617 369290 245669
rect 227542 245543 227594 245595
rect 247990 245543 248042 245595
rect 262678 245543 262730 245595
rect 369814 245543 369866 245595
rect 181366 245469 181418 245521
rect 253366 245469 253418 245521
rect 357622 245469 357674 245521
rect 202198 245395 202250 245447
rect 222454 245395 222506 245447
rect 252406 245395 252458 245447
rect 357142 245395 357194 245447
rect 168598 245321 168650 245373
rect 181270 245321 181322 245373
rect 261814 245321 261866 245373
rect 372022 245321 372074 245373
rect 260854 245247 260906 245299
rect 374038 245247 374090 245299
rect 211798 245173 211850 245225
rect 247606 245173 247658 245225
rect 261238 245173 261290 245225
rect 372886 245173 372938 245225
rect 389782 245173 389834 245225
rect 407062 245173 407114 245225
rect 211990 245099 212042 245151
rect 227446 245099 227498 245151
rect 260374 245099 260426 245151
rect 375766 245099 375818 245151
rect 227062 245025 227114 245077
rect 227926 245025 227978 245077
rect 246454 245025 246506 245077
rect 248086 245025 248138 245077
rect 260470 245025 260522 245077
rect 374614 245025 374666 245077
rect 42358 244951 42410 245003
rect 214198 244951 214250 245003
rect 216502 244951 216554 245003
rect 358486 244951 358538 245003
rect 210166 244877 210218 244929
rect 214102 244877 214154 244929
rect 247702 244877 247754 244929
rect 268246 244877 268298 244929
rect 97942 244803 97994 244855
rect 193270 244803 193322 244855
rect 144598 244729 144650 244781
rect 209686 244803 209738 244855
rect 213526 244803 213578 244855
rect 247990 244803 248042 244855
rect 292342 244877 292394 244929
rect 299542 244877 299594 244929
rect 307702 244877 307754 244929
rect 307798 244877 307850 244929
rect 309142 244877 309194 244929
rect 309622 244877 309674 244929
rect 328246 244877 328298 244929
rect 328534 244877 328586 244929
rect 368470 244877 368522 244929
rect 198934 244729 198986 244781
rect 227638 244729 227690 244781
rect 228118 244729 228170 244781
rect 248086 244729 248138 244781
rect 267862 244729 267914 244781
rect 102550 244655 102602 244707
rect 142966 244655 143018 244707
rect 259222 244655 259274 244707
rect 268822 244729 268874 244781
rect 268246 244655 268298 244707
rect 308086 244803 308138 244855
rect 278038 244729 278090 244781
rect 298006 244729 298058 244781
rect 298102 244729 298154 244781
rect 328630 244803 328682 244855
rect 348214 244803 348266 244855
rect 389782 244877 389834 244929
rect 368854 244803 368906 244855
rect 388534 244803 388586 244855
rect 608182 244803 608234 244855
rect 613462 244803 613514 244855
rect 309142 244729 309194 244781
rect 327958 244729 328010 244781
rect 328054 244729 328106 244781
rect 338614 244729 338666 244781
rect 277750 244655 277802 244707
rect 318166 244655 318218 244707
rect 326806 244655 326858 244707
rect 329014 244655 329066 244707
rect 389782 244655 389834 244707
rect 404374 244655 404426 244707
rect 138166 244581 138218 244633
rect 205750 244581 205802 244633
rect 235126 244581 235178 244633
rect 267190 244581 267242 244633
rect 277846 244581 277898 244633
rect 318262 244581 318314 244633
rect 135286 244507 135338 244559
rect 206998 244507 207050 244559
rect 242230 244507 242282 244559
rect 257782 244507 257834 244559
rect 262006 244507 262058 244559
rect 338134 244507 338186 244559
rect 132406 244433 132458 244485
rect 205462 244433 205514 244485
rect 277942 244433 277994 244485
rect 328054 244433 328106 244485
rect 42070 244359 42122 244411
rect 42550 244359 42602 244411
rect 126646 244359 126698 244411
rect 205270 244359 205322 244411
rect 260566 244359 260618 244411
rect 308758 244359 308810 244411
rect 123766 244285 123818 244337
rect 205078 244285 205130 244337
rect 258934 244285 258986 244337
rect 336694 244285 336746 244337
rect 674806 244285 674858 244337
rect 675286 244285 675338 244337
rect 120886 244211 120938 244263
rect 205654 244211 205706 244263
rect 257206 244211 257258 244263
rect 335926 244211 335978 244263
rect 383062 244211 383114 244263
rect 383446 244211 383498 244263
rect 118006 244137 118058 244189
rect 204502 244137 204554 244189
rect 211510 244137 211562 244189
rect 267862 244137 267914 244189
rect 267958 244137 268010 244189
rect 297910 244137 297962 244189
rect 298006 244137 298058 244189
rect 309910 244137 309962 244189
rect 312406 244137 312458 244189
rect 368758 244137 368810 244189
rect 112246 244063 112298 244115
rect 206422 244063 206474 244115
rect 251350 244063 251402 244115
rect 356278 244063 356330 244115
rect 109366 243989 109418 244041
rect 206230 243989 206282 244041
rect 249622 243989 249674 244041
rect 355798 243989 355850 244041
rect 106486 243915 106538 243967
rect 204598 243915 204650 243967
rect 257782 243915 257834 243967
rect 352150 243915 352202 243967
rect 103606 243841 103658 243893
rect 206614 243841 206666 243893
rect 243286 243841 243338 243893
rect 352630 243841 352682 243893
rect 100150 243767 100202 243819
rect 206518 243767 206570 243819
rect 244726 243767 244778 243819
rect 353590 243767 353642 243819
rect 94966 243693 95018 243745
rect 206326 243693 206378 243745
rect 246358 243693 246410 243745
rect 299494 243693 299546 243745
rect 92086 243619 92138 243671
rect 206038 243619 206090 243671
rect 247318 243619 247370 243671
rect 307702 243693 307754 243745
rect 354358 243693 354410 243745
rect 354838 243619 354890 243671
rect 86326 243545 86378 243597
rect 206710 243545 206762 243597
rect 237142 243545 237194 243597
rect 349942 243545 349994 243597
rect 80566 243471 80618 243523
rect 206902 243471 206954 243523
rect 240502 243471 240554 243523
rect 296662 243471 296714 243523
rect 297142 243471 297194 243523
rect 351478 243471 351530 243523
rect 77686 243397 77738 243449
rect 205174 243397 205226 243449
rect 230614 243397 230666 243449
rect 346678 243397 346730 243449
rect 69046 243323 69098 243375
rect 206134 243323 206186 243375
rect 227830 243323 227882 243375
rect 296662 243323 296714 243375
rect 297142 243323 297194 243375
rect 345526 243323 345578 243375
rect 235606 243249 235658 243301
rect 266134 243249 266186 243301
rect 270166 243249 270218 243301
rect 296758 243249 296810 243301
rect 297238 243249 297290 243301
rect 323062 243249 323114 243301
rect 282166 243175 282218 243227
rect 296662 243175 296714 243227
rect 296950 243175 297002 243227
rect 308374 243175 308426 243227
rect 308758 243175 308810 243227
rect 337270 243175 337322 243227
rect 266998 243101 267050 243153
rect 279766 243101 279818 243153
rect 279958 243101 280010 243153
rect 296758 243101 296810 243153
rect 267094 243027 267146 243079
rect 277846 243027 277898 243079
rect 287350 243027 287402 243079
rect 309430 243101 309482 243153
rect 318166 243101 318218 243153
rect 339574 243101 339626 243153
rect 318262 243027 318314 243079
rect 340342 243027 340394 243079
rect 267478 242953 267530 243005
rect 304150 242953 304202 243005
rect 675190 242953 675242 243005
rect 675382 242953 675434 243005
rect 265078 242879 265130 242931
rect 277750 242879 277802 242931
rect 284662 242879 284714 242931
rect 298102 242879 298154 242931
rect 263734 242805 263786 242857
rect 277942 242805 277994 242857
rect 270838 242731 270890 242783
rect 293398 242731 293450 242783
rect 293494 242731 293546 242783
rect 301270 242805 301322 242857
rect 293878 242731 293930 242783
rect 297910 242731 297962 242783
rect 316438 242731 316490 242783
rect 320854 242657 320906 242709
rect 264886 242583 264938 242635
rect 278038 242583 278090 242635
rect 284758 242583 284810 242635
rect 317110 242583 317162 242635
rect 267862 242509 267914 242561
rect 287446 242509 287498 242561
rect 287542 242509 287594 242561
rect 293494 242509 293546 242561
rect 297910 242509 297962 242561
rect 319126 242509 319178 242561
rect 269686 242435 269738 242487
rect 274486 242361 274538 242413
rect 289462 242361 289514 242413
rect 269206 242287 269258 242339
rect 287542 242287 287594 242339
rect 293974 242435 294026 242487
rect 297526 242435 297578 242487
rect 298102 242435 298154 242487
rect 317974 242435 318026 242487
rect 290806 242361 290858 242413
rect 321334 242361 321386 242413
rect 675094 242361 675146 242413
rect 675382 242361 675434 242413
rect 299254 242287 299306 242339
rect 299638 242287 299690 242339
rect 323446 242287 323498 242339
rect 141142 242213 141194 242265
rect 161110 242213 161162 242265
rect 288982 242213 289034 242265
rect 292342 242213 292394 242265
rect 292438 242213 292490 242265
rect 321910 242213 321962 242265
rect 270454 242139 270506 242191
rect 297622 242139 297674 242191
rect 298006 242139 298058 242191
rect 305398 242139 305450 242191
rect 317974 242139 318026 242191
rect 335638 242139 335690 242191
rect 40054 242065 40106 242117
rect 42358 242065 42410 242117
rect 157942 242065 157994 242117
rect 40150 241991 40202 242043
rect 43126 241991 43178 242043
rect 161110 241991 161162 242043
rect 284278 242065 284330 242117
rect 297910 242065 297962 242117
rect 298198 242065 298250 242117
rect 316918 242065 316970 242117
rect 319606 242065 319658 242117
rect 333430 242065 333482 242117
rect 177046 241991 177098 242043
rect 37366 241917 37418 241969
rect 42934 241917 42986 241969
rect 44566 241917 44618 241969
rect 141142 241917 141194 241969
rect 205846 241991 205898 242043
rect 238486 241843 238538 241895
rect 288982 241917 289034 241969
rect 250294 241843 250346 241895
rect 273046 241843 273098 241895
rect 273142 241843 273194 241895
rect 281878 241843 281930 241895
rect 283414 241843 283466 241895
rect 292246 241991 292298 242043
rect 293590 241991 293642 242043
rect 299638 241991 299690 242043
rect 290518 241917 290570 241969
rect 291574 241917 291626 241969
rect 292342 241917 292394 241969
rect 350518 241917 350570 241969
rect 360118 241917 360170 241969
rect 371830 241917 371882 241969
rect 289174 241843 289226 241895
rect 299734 241843 299786 241895
rect 306742 241843 306794 241895
rect 309142 241843 309194 241895
rect 314230 241843 314282 241895
rect 329974 241843 330026 241895
rect 338326 241843 338378 241895
rect 378358 241843 378410 241895
rect 217558 241769 217610 241821
rect 234742 241769 234794 241821
rect 248566 241769 248618 241821
rect 273910 241769 273962 241821
rect 274006 241769 274058 241821
rect 287062 241769 287114 241821
rect 219286 241695 219338 241747
rect 233974 241695 234026 241747
rect 255094 241695 255146 241747
rect 215446 241621 215498 241673
rect 272950 241621 273002 241673
rect 273046 241621 273098 241673
rect 273814 241621 273866 241673
rect 274102 241695 274154 241747
rect 290518 241769 290570 241821
rect 290614 241769 290666 241821
rect 287350 241695 287402 241747
rect 298102 241695 298154 241747
rect 289174 241621 289226 241673
rect 289366 241621 289418 241673
rect 296470 241621 296522 241673
rect 307606 241769 307658 241821
rect 309814 241769 309866 241821
rect 305590 241695 305642 241747
rect 308470 241695 308522 241747
rect 314422 241769 314474 241821
rect 315190 241769 315242 241821
rect 374422 241769 374474 241821
rect 395830 241843 395882 241895
rect 220438 241547 220490 241599
rect 233398 241547 233450 241599
rect 237718 241547 237770 241599
rect 261622 241547 261674 241599
rect 262006 241547 262058 241599
rect 328150 241695 328202 241747
rect 328246 241695 328298 241747
rect 339766 241695 339818 241747
rect 339862 241695 339914 241747
rect 360118 241695 360170 241747
rect 314422 241621 314474 241673
rect 316054 241621 316106 241673
rect 316630 241621 316682 241673
rect 375094 241621 375146 241673
rect 223222 241473 223274 241525
rect 232150 241473 232202 241525
rect 236950 241473 237002 241525
rect 263350 241473 263402 241525
rect 264310 241473 264362 241525
rect 271990 241473 272042 241525
rect 277942 241473 277994 241525
rect 314230 241473 314282 241525
rect 213910 241399 213962 241451
rect 229174 241399 229226 241451
rect 252790 241399 252842 241451
rect 325174 241547 325226 241599
rect 325270 241547 325322 241599
rect 328246 241547 328298 241599
rect 331510 241547 331562 241599
rect 314518 241399 314570 241451
rect 336502 241473 336554 241525
rect 339190 241547 339242 241599
rect 356566 241547 356618 241599
rect 361942 241547 361994 241599
rect 373942 241547 373994 241599
rect 359350 241473 359402 241525
rect 360982 241473 361034 241525
rect 379222 241769 379274 241821
rect 409270 241769 409322 241821
rect 377014 241695 377066 241747
rect 404950 241695 405002 241747
rect 379606 241621 379658 241673
rect 409942 241621 409994 241673
rect 674230 241547 674282 241599
rect 675478 241547 675530 241599
rect 380086 241473 380138 241525
rect 383542 241473 383594 241525
rect 383638 241473 383690 241525
rect 385558 241473 385610 241525
rect 277750 241325 277802 241377
rect 314614 241325 314666 241377
rect 317782 241325 317834 241377
rect 329590 241399 329642 241451
rect 333718 241399 333770 241451
rect 362902 241399 362954 241451
rect 363190 241399 363242 241451
rect 400150 241399 400202 241451
rect 327382 241325 327434 241377
rect 332950 241325 333002 241377
rect 333334 241325 333386 241377
rect 363286 241325 363338 241377
rect 364150 241325 364202 241377
rect 401878 241325 401930 241377
rect 277846 241251 277898 241303
rect 224086 241177 224138 241229
rect 231766 241177 231818 241229
rect 233302 241177 233354 241229
rect 238678 241177 238730 241229
rect 255958 241177 256010 241229
rect 310486 241177 310538 241229
rect 317878 241251 317930 241303
rect 330166 241251 330218 241303
rect 331030 241251 331082 241303
rect 358294 241251 358346 241303
rect 362038 241251 362090 241303
rect 373558 241251 373610 241303
rect 373942 241251 373994 241303
rect 397462 241251 397514 241303
rect 331702 241177 331754 241229
rect 363766 241177 363818 241229
rect 400726 241177 400778 241229
rect 225238 241103 225290 241155
rect 231190 241103 231242 241155
rect 222550 241029 222602 241081
rect 232534 241029 232586 241081
rect 216694 240955 216746 241007
rect 236182 240955 236234 241007
rect 227350 240881 227402 240933
rect 230326 240881 230378 240933
rect 212758 240807 212810 240859
rect 233206 240807 233258 240859
rect 219286 240733 219338 240785
rect 250678 241103 250730 241155
rect 254998 241103 255050 241155
rect 314518 241103 314570 241155
rect 314614 241103 314666 241155
rect 332758 241103 332810 241155
rect 364246 241103 364298 241155
rect 402742 241103 402794 241155
rect 41782 240585 41834 240637
rect 219670 240585 219722 240637
rect 249814 241029 249866 241081
rect 254230 241029 254282 241081
rect 337846 241029 337898 241081
rect 362902 241029 362954 241081
rect 364342 241029 364394 241081
rect 373558 241029 373610 241081
rect 398422 241029 398474 241081
rect 244438 240955 244490 241007
rect 326902 240955 326954 241007
rect 326998 240955 327050 241007
rect 338326 240955 338378 241007
rect 362422 240955 362474 241007
rect 398998 240955 399050 241007
rect 237910 240881 237962 240933
rect 252886 240881 252938 240933
rect 253750 240881 253802 240933
rect 339382 240881 339434 240933
rect 339478 240881 339530 240933
rect 362230 240881 362282 240933
rect 365974 240881 366026 240933
rect 406102 240881 406154 240933
rect 237814 240807 237866 240859
rect 252022 240807 252074 240859
rect 252310 240807 252362 240859
rect 342646 240807 342698 240859
rect 366358 240807 366410 240859
rect 407158 240807 407210 240859
rect 251542 240733 251594 240785
rect 344182 240733 344234 240785
rect 365014 240733 365066 240785
rect 404470 240733 404522 240785
rect 249814 240659 249866 240711
rect 347446 240659 347498 240711
rect 367222 240659 367274 240711
rect 408886 240659 408938 240711
rect 250582 240585 250634 240637
rect 345718 240585 345770 240637
rect 364630 240585 364682 240637
rect 403414 240585 403466 240637
rect 220630 240511 220682 240563
rect 247894 240511 247946 240563
rect 248374 240511 248426 240563
rect 350422 240511 350474 240563
rect 365398 240511 365450 240563
rect 405238 240511 405290 240563
rect 674998 240511 675050 240563
rect 675478 240511 675530 240563
rect 144598 240437 144650 240489
rect 162742 240437 162794 240489
rect 220246 240437 220298 240489
rect 248662 240437 248714 240489
rect 249334 240437 249386 240489
rect 349174 240437 349226 240489
rect 366454 240437 366506 240489
rect 407734 240437 407786 240489
rect 41782 240363 41834 240415
rect 218518 240363 218570 240415
rect 237814 240363 237866 240415
rect 238966 240363 239018 240415
rect 263926 240363 263978 240415
rect 275734 240363 275786 240415
rect 283030 240363 283082 240415
rect 313366 240363 313418 240415
rect 370294 240363 370346 240415
rect 378262 240363 378314 240415
rect 408214 240363 408266 240415
rect 237334 240289 237386 240341
rect 262198 240289 262250 240341
rect 262294 240289 262346 240341
rect 277942 240289 277994 240341
rect 278038 240289 278090 240341
rect 288406 240289 288458 240341
rect 289174 240289 289226 240341
rect 306934 240289 306986 240341
rect 314614 240289 314666 240341
rect 373270 240289 373322 240341
rect 377878 240289 377930 240341
rect 407542 240289 407594 240341
rect 225430 240215 225482 240267
rect 230902 240215 230954 240267
rect 238774 240215 238826 240267
rect 259414 240215 259466 240267
rect 276790 240215 276842 240267
rect 283894 240215 283946 240267
rect 218422 240141 218474 240193
rect 237910 240141 237962 240193
rect 244150 240141 244202 240193
rect 246358 240141 246410 240193
rect 257206 240141 257258 240193
rect 277846 240141 277898 240193
rect 277942 240141 277994 240193
rect 286774 240141 286826 240193
rect 296566 240215 296618 240267
rect 298102 240215 298154 240267
rect 311638 240215 311690 240267
rect 314230 240215 314282 240267
rect 372406 240215 372458 240267
rect 376438 240215 376490 240267
rect 226294 240067 226346 240119
rect 230710 240067 230762 240119
rect 236470 240067 236522 240119
rect 264406 240067 264458 240119
rect 277654 240067 277706 240119
rect 236278 239993 236330 240045
rect 241654 239993 241706 240045
rect 256438 239993 256490 240045
rect 277750 239993 277802 240045
rect 279478 240067 279530 240119
rect 295798 240141 295850 240193
rect 295894 240141 295946 240193
rect 313174 240141 313226 240193
rect 313462 240141 313514 240193
rect 371350 240141 371402 240193
rect 373078 240141 373130 240193
rect 386806 240141 386858 240193
rect 386998 240215 387050 240267
rect 403222 240215 403274 240267
rect 404086 240141 404138 240193
rect 288214 240067 288266 240119
rect 300598 240067 300650 240119
rect 316822 240067 316874 240119
rect 326998 240067 327050 240119
rect 329302 240067 329354 240119
rect 354550 240067 354602 240119
rect 360598 240067 360650 240119
rect 378742 240067 378794 240119
rect 381814 240067 381866 240119
rect 383062 240067 383114 240119
rect 289078 239993 289130 240045
rect 292630 239993 292682 240045
rect 294262 239993 294314 240045
rect 303574 239993 303626 240045
rect 304726 239993 304778 240045
rect 308182 239993 308234 240045
rect 310486 239993 310538 240045
rect 221494 239919 221546 239971
rect 232918 239919 232970 239971
rect 238294 239919 238346 239971
rect 260662 239919 260714 239971
rect 268726 239919 268778 239971
rect 280342 239919 280394 239971
rect 286966 239919 287018 239971
rect 297622 239919 297674 239971
rect 298198 239919 298250 239971
rect 312790 239919 312842 239971
rect 313750 239919 313802 239971
rect 325270 239919 325322 239971
rect 334390 239993 334442 240045
rect 334486 239993 334538 240045
rect 365878 239993 365930 240045
rect 377206 239993 377258 240045
rect 405526 239993 405578 240045
rect 327862 239919 327914 239971
rect 351766 239919 351818 239971
rect 360214 239919 360266 239971
rect 378646 239919 378698 239971
rect 234550 239845 234602 239897
rect 238582 239845 238634 239897
rect 277078 239845 277130 239897
rect 283798 239845 283850 239897
rect 283894 239845 283946 239897
rect 295222 239845 295274 239897
rect 295702 239845 295754 239897
rect 218710 239771 218762 239823
rect 234358 239771 234410 239823
rect 274870 239771 274922 239823
rect 228022 239697 228074 239749
rect 229942 239697 229994 239749
rect 241078 239697 241130 239749
rect 244630 239697 244682 239749
rect 269398 239697 269450 239749
rect 276310 239697 276362 239749
rect 277654 239771 277706 239823
rect 282934 239771 282986 239823
rect 283030 239771 283082 239823
rect 294742 239771 294794 239823
rect 299062 239771 299114 239823
rect 305782 239771 305834 239823
rect 278038 239697 278090 239749
rect 278230 239697 278282 239749
rect 281782 239697 281834 239749
rect 281878 239697 281930 239749
rect 292150 239697 292202 239749
rect 292246 239697 292298 239749
rect 297910 239697 297962 239749
rect 302998 239697 303050 239749
rect 307606 239697 307658 239749
rect 326614 239845 326666 239897
rect 348694 239845 348746 239897
rect 375670 239845 375722 239897
rect 383062 239919 383114 239971
rect 380854 239845 380906 239897
rect 388150 239845 388202 239897
rect 314806 239771 314858 239823
rect 327094 239771 327146 239823
rect 350038 239771 350090 239823
rect 380566 239771 380618 239823
rect 384886 239771 384938 239823
rect 308854 239697 308906 239749
rect 310198 239697 310250 239749
rect 311638 239697 311690 239749
rect 323638 239697 323690 239749
rect 214486 239623 214538 239675
rect 225142 239623 225194 239675
rect 229078 239623 229130 239675
rect 230230 239623 230282 239675
rect 238198 239623 238250 239675
rect 241846 239623 241898 239675
rect 265654 239623 265706 239675
rect 270166 239623 270218 239675
rect 270262 239623 270314 239675
rect 272278 239623 272330 239675
rect 226294 239549 226346 239601
rect 235798 239549 235850 239601
rect 271414 239549 271466 239601
rect 277942 239623 277994 239675
rect 278902 239623 278954 239675
rect 279670 239623 279722 239675
rect 280534 239623 280586 239675
rect 275350 239549 275402 239601
rect 281110 239549 281162 239601
rect 273526 239475 273578 239527
rect 281590 239475 281642 239527
rect 285046 239475 285098 239527
rect 287062 239623 287114 239675
rect 290806 239623 290858 239675
rect 304054 239623 304106 239675
rect 307990 239623 308042 239675
rect 309526 239623 309578 239675
rect 310294 239623 310346 239675
rect 315670 239623 315722 239675
rect 328822 239697 328874 239749
rect 330070 239697 330122 239749
rect 339190 239697 339242 239749
rect 376054 239697 376106 239749
rect 386998 239697 387050 239749
rect 325654 239623 325706 239675
rect 328630 239623 328682 239675
rect 328726 239623 328778 239675
rect 353494 239623 353546 239675
rect 374806 239623 374858 239675
rect 382678 239623 382730 239675
rect 383254 239623 383306 239675
rect 396406 239623 396458 239675
rect 286678 239549 286730 239601
rect 292534 239549 292586 239601
rect 292630 239549 292682 239601
rect 298006 239549 298058 239601
rect 301846 239549 301898 239601
rect 306838 239549 306890 239601
rect 306934 239549 306986 239601
rect 313846 239549 313898 239601
rect 324406 239549 324458 239601
rect 343702 239549 343754 239601
rect 373846 239549 373898 239601
rect 398614 239549 398666 239601
rect 275926 239401 275978 239453
rect 286006 239401 286058 239453
rect 296950 239475 297002 239527
rect 297622 239475 297674 239527
rect 312598 239475 312650 239527
rect 321622 239475 321674 239527
rect 338902 239475 338954 239527
rect 291862 239401 291914 239453
rect 42550 239327 42602 239379
rect 275446 239327 275498 239379
rect 287734 239327 287786 239379
rect 287830 239327 287882 239379
rect 288982 239327 289034 239379
rect 42358 239253 42410 239305
rect 215926 239253 215978 239305
rect 218902 239253 218954 239305
rect 272470 239253 272522 239305
rect 285526 239253 285578 239305
rect 287254 239253 287306 239305
rect 297526 239401 297578 239453
rect 297814 239401 297866 239453
rect 305014 239401 305066 239453
rect 323062 239401 323114 239453
rect 292054 239327 292106 239379
rect 302422 239327 302474 239379
rect 302518 239327 302570 239379
rect 307222 239327 307274 239379
rect 320854 239327 320906 239379
rect 324694 239327 324746 239379
rect 324886 239401 324938 239453
rect 331318 239401 331370 239453
rect 361558 239401 361610 239453
rect 383062 239475 383114 239527
rect 378646 239401 378698 239453
rect 392086 239401 392138 239453
rect 341302 239327 341354 239379
rect 380086 239327 380138 239379
rect 386614 239327 386666 239379
rect 386710 239327 386762 239379
rect 406678 239327 406730 239379
rect 293206 239253 293258 239305
rect 302806 239253 302858 239305
rect 323446 239253 323498 239305
rect 341974 239253 342026 239305
rect 378742 239253 378794 239305
rect 394102 239253 394154 239305
rect 42550 239179 42602 239231
rect 43222 239179 43274 239231
rect 240502 239179 240554 239231
rect 255670 239179 255722 239231
rect 276214 239179 276266 239231
rect 280438 239179 280490 239231
rect 291478 239179 291530 239231
rect 301846 239179 301898 239231
rect 318262 239179 318314 239231
rect 324886 239179 324938 239231
rect 328630 239179 328682 239231
rect 346966 239179 347018 239231
rect 378646 239179 378698 239231
rect 383830 239179 383882 239231
rect 386806 239179 386858 239231
rect 396886 239179 396938 239231
rect 273238 239105 273290 239157
rect 286678 239105 286730 239157
rect 286774 239105 286826 239157
rect 289366 239105 289418 239157
rect 291862 239105 291914 239157
rect 299158 239105 299210 239157
rect 322678 239105 322730 239157
rect 340918 239105 340970 239157
rect 377494 239105 377546 239157
rect 386710 239105 386762 239157
rect 236182 239031 236234 239083
rect 238390 239031 238442 239083
rect 271894 239031 271946 239083
rect 287830 239031 287882 239083
rect 288982 239031 289034 239083
rect 294454 239031 294506 239083
rect 295990 239031 296042 239083
rect 304054 239031 304106 239083
rect 321238 239031 321290 239083
rect 337174 239031 337226 239083
rect 339862 239031 339914 239083
rect 340246 239031 340298 239083
rect 375190 239031 375242 239083
rect 400630 239031 400682 239083
rect 142966 238957 143018 239009
rect 211030 238957 211082 239009
rect 216694 238957 216746 239009
rect 228118 238957 228170 239009
rect 231958 238957 232010 239009
rect 237526 238957 237578 239009
rect 268150 238957 268202 239009
rect 268246 238957 268298 239009
rect 270934 238957 270986 239009
rect 278518 238957 278570 239009
rect 280726 238957 280778 239009
rect 290902 238957 290954 239009
rect 293302 238957 293354 239009
rect 294070 238957 294122 239009
rect 303190 238957 303242 239009
rect 316438 238957 316490 239009
rect 377302 238957 377354 239009
rect 380470 238957 380522 239009
rect 387574 238957 387626 239009
rect 240118 238883 240170 238935
rect 256822 238883 256874 238935
rect 258262 238883 258314 238935
rect 226870 238809 226922 238861
rect 235030 238809 235082 238861
rect 239158 238809 239210 238861
rect 258550 238809 258602 238861
rect 317686 238883 317738 238935
rect 325942 238883 325994 238935
rect 326710 238883 326762 238935
rect 328918 238883 328970 238935
rect 331894 238883 331946 238935
rect 360502 238883 360554 238935
rect 366838 238883 366890 238935
rect 224566 238735 224618 238787
rect 239542 238735 239594 238787
rect 257782 238735 257834 238787
rect 256054 238661 256106 238713
rect 308950 238735 309002 238787
rect 329110 238809 329162 238861
rect 330646 238809 330698 238861
rect 357238 238809 357290 238861
rect 368182 238809 368234 238861
rect 375958 238809 376010 238861
rect 381430 238883 381482 238935
rect 389206 238883 389258 238935
rect 383350 238809 383402 238861
rect 318166 238735 318218 238787
rect 318646 238735 318698 238787
rect 332182 238735 332234 238787
rect 332278 238735 332330 238787
rect 345910 238735 345962 238787
rect 258838 238661 258890 238713
rect 325846 238661 325898 238713
rect 325942 238661 325994 238713
rect 327574 238661 327626 238713
rect 331126 238661 331178 238713
rect 358774 238735 358826 238787
rect 368566 238735 368618 238787
rect 379030 238735 379082 238787
rect 379702 238735 379754 238787
rect 385366 238735 385418 238787
rect 217078 238587 217130 238639
rect 255190 238587 255242 238639
rect 255574 238587 255626 238639
rect 317974 238587 318026 238639
rect 320086 238587 320138 238639
rect 322102 238587 322154 238639
rect 322294 238587 322346 238639
rect 42166 238513 42218 238565
rect 42358 238513 42410 238565
rect 253846 238513 253898 238565
rect 318070 238513 318122 238565
rect 318166 238513 318218 238565
rect 322390 238513 322442 238565
rect 322486 238513 322538 238565
rect 331606 238513 331658 238565
rect 331798 238587 331850 238639
rect 332086 238587 332138 238639
rect 351382 238661 351434 238713
rect 358870 238661 358922 238713
rect 372598 238661 372650 238713
rect 383062 238661 383114 238713
rect 334102 238587 334154 238639
rect 365302 238587 365354 238639
rect 368662 238587 368714 238639
rect 387094 238587 387146 238639
rect 334966 238513 335018 238565
rect 218038 238439 218090 238491
rect 253462 238439 253514 238491
rect 254614 238439 254666 238491
rect 335350 238513 335402 238565
rect 348022 238513 348074 238565
rect 375958 238513 376010 238565
rect 384598 238513 384650 238565
rect 336982 238439 337034 238491
rect 369430 238439 369482 238491
rect 388822 238439 388874 238491
rect 216310 238365 216362 238417
rect 237526 238365 237578 238417
rect 240598 238365 240650 238417
rect 317686 238365 317738 238417
rect 318070 238365 318122 238417
rect 253366 238291 253418 238343
rect 322486 238365 322538 238417
rect 330742 238365 330794 238417
rect 335254 238365 335306 238417
rect 367030 238365 367082 238417
rect 371638 238365 371690 238417
rect 393622 238365 393674 238417
rect 252406 238217 252458 238269
rect 321910 238217 321962 238269
rect 338710 238291 338762 238343
rect 370390 238291 370442 238343
rect 390358 238291 390410 238343
rect 639766 238291 639818 238343
rect 649942 238291 649994 238343
rect 251638 238143 251690 238195
rect 331606 238217 331658 238269
rect 341494 238217 341546 238269
rect 369814 238217 369866 238269
rect 389686 238217 389738 238269
rect 228214 238069 228266 238121
rect 245878 238069 245930 238121
rect 251158 238069 251210 238121
rect 340438 238143 340490 238195
rect 370870 238143 370922 238195
rect 391894 238143 391946 238195
rect 222838 237995 222890 238047
rect 243766 237995 243818 238047
rect 249430 237995 249482 238047
rect 321910 237995 321962 238047
rect 322102 237995 322154 238047
rect 223318 237921 223370 237973
rect 242422 237921 242474 237973
rect 250198 237921 250250 237973
rect 315862 237921 315914 237973
rect 42166 237847 42218 237899
rect 47542 237847 47594 237899
rect 222934 237847 222986 237899
rect 221878 237773 221930 237825
rect 228502 237847 228554 237899
rect 230806 237847 230858 237899
rect 247990 237847 248042 237899
rect 322294 237921 322346 237973
rect 322486 237995 322538 238047
rect 326806 237995 326858 238047
rect 343510 238069 343562 238121
rect 372022 238069 372074 238121
rect 394198 238069 394250 238121
rect 345238 237995 345290 238047
rect 371254 237995 371306 238047
rect 392470 237995 392522 238047
rect 346294 237921 346346 237973
rect 375286 237921 375338 237973
rect 401206 237921 401258 237973
rect 639382 237921 639434 237973
rect 649750 237921 649802 237973
rect 316054 237847 316106 237899
rect 221494 237699 221546 237751
rect 228214 237699 228266 237751
rect 242614 237773 242666 237825
rect 247222 237773 247274 237825
rect 315766 237773 315818 237825
rect 315862 237773 315914 237825
rect 322006 237773 322058 237825
rect 326806 237847 326858 237899
rect 351286 237847 351338 237899
rect 362806 237847 362858 237899
rect 382294 237847 382346 237899
rect 384118 237847 384170 237899
rect 410422 237847 410474 237899
rect 637942 237847 637994 237899
rect 650422 237847 650474 237899
rect 353014 237773 353066 237825
rect 359830 237773 359882 237825
rect 380950 237773 381002 237825
rect 384502 237773 384554 237825
rect 410998 237773 411050 237825
rect 638902 237773 638954 237825
rect 649558 237773 649610 237825
rect 244822 237699 244874 237751
rect 245782 237699 245834 237751
rect 356182 237699 356234 237751
rect 637366 237699 637418 237751
rect 650134 237699 650186 237751
rect 224086 237625 224138 237677
rect 240694 237625 240746 237677
rect 246742 237625 246794 237677
rect 315574 237625 315626 237677
rect 322390 237625 322442 237677
rect 354454 237625 354506 237677
rect 549238 237625 549290 237677
rect 650998 237625 651050 237677
rect 148342 237551 148394 237603
rect 207094 237551 207146 237603
rect 221974 237551 222026 237603
rect 223702 237551 223754 237603
rect 241558 237551 241610 237603
rect 245014 237551 245066 237603
rect 357814 237551 357866 237603
rect 374230 237551 374282 237603
rect 399670 237551 399722 237603
rect 420598 237551 420650 237603
rect 608182 237551 608234 237603
rect 637846 237551 637898 237603
rect 650230 237551 650282 237603
rect 256822 237477 256874 237529
rect 310006 237477 310058 237529
rect 248950 237403 249002 237455
rect 258838 237403 258890 237455
rect 268150 237403 268202 237455
rect 282262 237403 282314 237455
rect 286486 237403 286538 237455
rect 287158 237403 287210 237455
rect 292534 237403 292586 237455
rect 293686 237403 293738 237455
rect 293782 237403 293834 237455
rect 295414 237403 295466 237455
rect 304726 237403 304778 237455
rect 315382 237403 315434 237455
rect 239542 237329 239594 237381
rect 257398 237329 257450 237381
rect 274198 237329 274250 237381
rect 281494 237329 281546 237381
rect 281686 237329 281738 237381
rect 286774 237329 286826 237381
rect 291286 237329 291338 237381
rect 317590 237477 317642 237529
rect 319030 237477 319082 237529
rect 332374 237477 332426 237529
rect 332758 237477 332810 237529
rect 347926 237477 347978 237529
rect 373462 237477 373514 237529
rect 397942 237477 397994 237529
rect 315574 237403 315626 237455
rect 322390 237403 322442 237455
rect 322486 237403 322538 237455
rect 317398 237329 317450 237381
rect 368566 237329 368618 237381
rect 372982 237403 373034 237455
rect 396214 237403 396266 237455
rect 376630 237329 376682 237381
rect 225526 237255 225578 237307
rect 237430 237255 237482 237307
rect 276694 237255 276746 237307
rect 284470 237255 284522 237307
rect 287158 237255 287210 237307
rect 299638 237255 299690 237307
rect 299734 237255 299786 237307
rect 322294 237255 322346 237307
rect 322774 237255 322826 237307
rect 358390 237255 358442 237307
rect 369046 237255 369098 237307
rect 227350 237181 227402 237233
rect 233494 237181 233546 237233
rect 275830 237181 275882 237233
rect 286582 237181 286634 237233
rect 273526 237107 273578 237159
rect 291670 237181 291722 237233
rect 291382 237107 291434 237159
rect 302326 237107 302378 237159
rect 305878 237107 305930 237159
rect 315574 237181 315626 237233
rect 316630 237181 316682 237233
rect 339862 237181 339914 237233
rect 380182 237255 380234 237307
rect 385942 237255 385994 237307
rect 387670 237181 387722 237233
rect 318454 237107 318506 237159
rect 322486 237107 322538 237159
rect 329686 237107 329738 237159
rect 355702 237107 355754 237159
rect 379990 237107 380042 237159
rect 380182 237107 380234 237159
rect 221110 237033 221162 237085
rect 246550 237033 246602 237085
rect 282742 237033 282794 237085
rect 227254 236959 227306 237011
rect 234070 236959 234122 237011
rect 277270 236959 277322 237011
rect 279766 236959 279818 237011
rect 220726 236885 220778 236937
rect 246934 236885 246986 236937
rect 271030 236885 271082 236937
rect 288982 236959 289034 237011
rect 289270 237033 289322 237085
rect 300982 237033 301034 237085
rect 310006 237033 310058 237085
rect 324118 237033 324170 237085
rect 327478 237033 327530 237085
rect 350710 237033 350762 237085
rect 298006 236959 298058 237011
rect 300790 236959 300842 237011
rect 306262 236959 306314 237011
rect 326710 236959 326762 237011
rect 349558 236959 349610 237011
rect 284374 236885 284426 236937
rect 298774 236885 298826 236937
rect 326230 236885 326282 236937
rect 332758 236885 332810 236937
rect 332854 236885 332906 236937
rect 339478 236885 339530 236937
rect 217462 236811 217514 236863
rect 254326 236811 254378 236863
rect 278806 236811 278858 236863
rect 274678 236737 274730 236789
rect 294358 236737 294410 236789
rect 295318 236811 295370 236863
rect 303670 236811 303722 236863
rect 308950 236811 309002 236863
rect 333910 236811 333962 236863
rect 370774 236811 370826 236863
rect 381142 236811 381194 236863
rect 296182 236737 296234 236789
rect 328246 236737 328298 236789
rect 352438 236737 352490 236789
rect 42166 236663 42218 236715
rect 42934 236663 42986 236715
rect 278422 236663 278474 236715
rect 279382 236663 279434 236715
rect 285814 236663 285866 236715
rect 299254 236663 299306 236715
rect 324502 236663 324554 236715
rect 344758 236663 344810 236715
rect 381910 236663 381962 236715
rect 390934 236663 390986 236715
rect 258166 236589 258218 236641
rect 262294 236589 262346 236641
rect 268342 236589 268394 236641
rect 281398 236589 281450 236641
rect 288694 236589 288746 236641
rect 312118 236589 312170 236641
rect 325270 236589 325322 236641
rect 331702 236589 331754 236641
rect 274102 236515 274154 236567
rect 289654 236515 289706 236567
rect 289942 236515 289994 236567
rect 304726 236515 304778 236567
rect 324022 236515 324074 236567
rect 343030 236589 343082 236641
rect 225046 236441 225098 236493
rect 238870 236441 238922 236493
rect 276406 236441 276458 236493
rect 294838 236441 294890 236493
rect 321814 236441 321866 236493
rect 338230 236515 338282 236567
rect 205942 236367 205994 236419
rect 272662 236367 272714 236419
rect 146806 236219 146858 236271
rect 168406 236219 168458 236271
rect 271510 236293 271562 236345
rect 227734 236219 227786 236271
rect 232822 236219 232874 236271
rect 236566 236219 236618 236271
rect 238966 236219 239018 236271
rect 278134 236219 278186 236271
rect 281206 236219 281258 236271
rect 281398 236293 281450 236345
rect 288118 236293 288170 236345
rect 288982 236367 289034 236419
rect 297334 236367 297386 236419
rect 289366 236219 289418 236271
rect 145558 236145 145610 236197
rect 146422 236145 146474 236197
rect 146710 236145 146762 236197
rect 174166 236145 174218 236197
rect 205942 236145 205994 236197
rect 210262 236145 210314 236197
rect 210646 236145 210698 236197
rect 213046 236145 213098 236197
rect 225910 236145 225962 236197
rect 236758 236145 236810 236197
rect 290326 236293 290378 236345
rect 301462 236293 301514 236345
rect 332278 236293 332330 236345
rect 361078 236293 361130 236345
rect 290806 236219 290858 236271
rect 293974 236219 294026 236271
rect 297526 236219 297578 236271
rect 300214 236219 300266 236271
rect 319990 236219 320042 236271
rect 334198 236219 334250 236271
rect 335062 236219 335114 236271
rect 335254 236219 335306 236271
rect 290902 236145 290954 236197
rect 291766 236145 291818 236197
rect 319318 236145 319370 236197
rect 320470 236145 320522 236197
rect 336118 236145 336170 236197
rect 541462 236145 541514 236197
rect 549238 236145 549290 236197
rect 638710 236145 638762 236197
rect 639190 236145 639242 236197
rect 265942 236071 265994 236123
rect 339958 236071 340010 236123
rect 264790 235997 264842 236049
rect 310774 235997 310826 236049
rect 312982 235997 313034 236049
rect 369622 235997 369674 236049
rect 267670 235923 267722 235975
rect 340726 235923 340778 235975
rect 262870 235849 262922 235901
rect 338518 235849 338570 235901
rect 258358 235775 258410 235827
rect 336310 235775 336362 235827
rect 261142 235701 261194 235753
rect 337750 235701 337802 235753
rect 256342 235627 256394 235679
rect 335542 235627 335594 235679
rect 260086 235553 260138 235605
rect 336982 235553 337034 235605
rect 273910 235479 273962 235531
rect 355414 235479 355466 235531
rect 42166 235405 42218 235457
rect 43030 235405 43082 235457
rect 236086 235405 236138 235457
rect 265462 235405 265514 235457
rect 273814 235405 273866 235457
rect 356182 235405 356234 235457
rect 245686 235331 245738 235383
rect 353974 235331 354026 235383
rect 239350 235257 239402 235309
rect 350998 235257 351050 235309
rect 146134 235183 146186 235235
rect 146422 235183 146474 235235
rect 246358 235183 246410 235235
rect 353206 235183 353258 235235
rect 241846 235109 241898 235161
rect 350038 235109 350090 235161
rect 238678 235035 238730 235087
rect 347830 235035 347882 235087
rect 241654 234961 241706 235013
rect 349558 234961 349610 235013
rect 244630 234887 244682 234939
rect 351766 234887 351818 234939
rect 42166 234813 42218 234865
rect 42358 234813 42410 234865
rect 238582 234813 238634 234865
rect 348790 234813 348842 234865
rect 231670 234739 231722 234791
rect 347350 234739 347402 234791
rect 226966 234665 227018 234717
rect 345142 234665 345194 234717
rect 265270 234591 265322 234643
rect 308854 234591 308906 234643
rect 312022 234591 312074 234643
rect 367702 234591 367754 234643
rect 266614 234517 266666 234569
rect 306742 234517 306794 234569
rect 316054 234517 316106 234569
rect 322390 234517 322442 234569
rect 266038 234443 266090 234495
rect 307318 234443 307370 234495
rect 368566 234443 368618 234495
rect 379990 234443 380042 234495
rect 283318 234369 283370 234421
rect 320374 234369 320426 234421
rect 283702 234295 283754 234347
rect 319702 234295 319754 234347
rect 383062 234295 383114 234347
rect 384406 234295 384458 234347
rect 267094 234221 267146 234273
rect 305110 234221 305162 234273
rect 42070 234147 42122 234199
rect 43126 234147 43178 234199
rect 267862 234147 267914 234199
rect 303382 234147 303434 234199
rect 268822 234073 268874 234125
rect 301942 234073 301994 234125
rect 269302 233999 269354 234051
rect 300310 233999 300362 234051
rect 293494 233925 293546 233977
rect 322582 233925 322634 233977
rect 269878 233851 269930 233903
rect 301366 233851 301418 233903
rect 286486 233777 286538 233829
rect 314326 233777 314378 233829
rect 292870 233703 292922 233755
rect 321430 233703 321482 233755
rect 210358 233629 210410 233681
rect 212374 233629 212426 233681
rect 286102 233629 286154 233681
rect 315094 233629 315146 233681
rect 208054 233555 208106 233607
rect 213526 233555 213578 233607
rect 269110 233555 269162 233607
rect 270262 233555 270314 233607
rect 298582 233555 298634 233607
rect 210070 233481 210122 233533
rect 213142 233481 213194 233533
rect 213910 233481 213962 233533
rect 209974 233407 210026 233459
rect 289846 233481 289898 233533
rect 295702 233481 295754 233533
rect 297046 233481 297098 233533
rect 146806 233259 146858 233311
rect 171286 233259 171338 233311
rect 645718 232889 645770 232941
rect 649846 232889 649898 232941
rect 42262 232519 42314 232571
rect 43222 232519 43274 232571
rect 645142 232297 645194 232349
rect 645526 232297 645578 232349
rect 649654 232297 649706 232349
rect 204982 232075 205034 232127
rect 205558 232075 205610 232127
rect 645142 231557 645194 231609
rect 650518 231557 650570 231609
rect 645142 231113 645194 231165
rect 645334 231113 645386 231165
rect 650326 231113 650378 231165
rect 645142 230669 645194 230721
rect 650038 230669 650090 230721
rect 146806 230521 146858 230573
rect 151126 230521 151178 230573
rect 144406 230447 144458 230499
rect 165526 230447 165578 230499
rect 666646 229485 666698 229537
rect 674422 229485 674474 229537
rect 669622 228893 669674 228945
rect 674710 228893 674762 228945
rect 146806 228745 146858 228797
rect 159766 228745 159818 228797
rect 669718 227857 669770 227909
rect 674422 227857 674474 227909
rect 146710 227635 146762 227687
rect 162646 227635 162698 227687
rect 43222 227561 43274 227613
rect 43510 227561 43562 227613
rect 146806 227561 146858 227613
rect 202966 227561 203018 227613
rect 146326 227487 146378 227539
rect 146518 227487 146570 227539
rect 205078 227413 205130 227465
rect 207382 227413 207434 227465
rect 144022 226377 144074 226429
rect 156886 226377 156938 226429
rect 673366 225785 673418 225837
rect 674710 225785 674762 225837
rect 679798 225785 679850 225837
rect 206134 224823 206186 224875
rect 144022 224675 144074 224727
rect 200086 224675 200138 224727
rect 673846 224675 673898 224727
rect 679990 224675 680042 224727
rect 141046 224601 141098 224653
rect 204502 224601 204554 224653
rect 206134 224601 206186 224653
rect 146614 224527 146666 224579
rect 205462 224527 205514 224579
rect 206422 224527 206474 224579
rect 206806 224527 206858 224579
rect 149686 224453 149738 224505
rect 204598 224453 204650 224505
rect 152566 224379 152618 224431
rect 206422 224379 206474 224431
rect 144022 221863 144074 221915
rect 179926 221863 179978 221915
rect 144118 221789 144170 221841
rect 182806 221789 182858 221841
rect 146134 221715 146186 221767
rect 146230 221715 146282 221767
rect 155446 221715 155498 221767
rect 204502 221715 204554 221767
rect 161206 221641 161258 221693
rect 204982 221641 205034 221693
rect 164086 221567 164138 221619
rect 205366 221567 205418 221619
rect 166966 221493 167018 221545
rect 206902 221493 206954 221545
rect 169846 221419 169898 221471
rect 204598 221419 204650 221471
rect 42358 221049 42410 221101
rect 44950 221049 45002 221101
rect 42358 220309 42410 220361
rect 45142 220309 45194 220361
rect 42358 219421 42410 219473
rect 44854 219421 44906 219473
rect 144022 218903 144074 218955
rect 177142 218903 177194 218955
rect 175606 218829 175658 218881
rect 204502 218829 204554 218881
rect 178486 218755 178538 218807
rect 204598 218755 204650 218807
rect 181366 218681 181418 218733
rect 204694 218681 204746 218733
rect 184246 218607 184298 218659
rect 205366 218607 205418 218659
rect 146518 217719 146570 217771
rect 146518 217571 146570 217623
rect 144022 216017 144074 216069
rect 174262 216017 174314 216069
rect 187126 215943 187178 215995
rect 204790 215943 204842 215995
rect 192886 215869 192938 215921
rect 204502 215869 204554 215921
rect 146422 213427 146474 213479
rect 146710 213427 146762 213479
rect 146422 213279 146474 213331
rect 171382 213279 171434 213331
rect 144118 213205 144170 213257
rect 154006 213205 154058 213257
rect 144022 213131 144074 213183
rect 148246 213131 148298 213183
rect 205558 213131 205610 213183
rect 207190 213131 207242 213183
rect 679798 212243 679850 212295
rect 680086 212243 680138 212295
rect 146230 211577 146282 211629
rect 146518 211577 146570 211629
rect 647926 210245 647978 210297
rect 679798 210245 679850 210297
rect 144022 207433 144074 207485
rect 165622 207433 165674 207485
rect 144118 207359 144170 207411
rect 168502 207359 168554 207411
rect 674614 207359 674666 207411
rect 676822 207359 676874 207411
rect 674422 205731 674474 205783
rect 675478 205731 675530 205783
rect 675190 205139 675242 205191
rect 675478 205139 675530 205191
rect 42358 204473 42410 204525
rect 43030 204473 43082 204525
rect 144022 204473 144074 204525
rect 148438 204473 148490 204525
rect 673942 204399 673994 204451
rect 675382 204399 675434 204451
rect 42358 204325 42410 204377
rect 44566 204325 44618 204377
rect 674998 202179 675050 202231
rect 675286 202179 675338 202231
rect 675094 202031 675146 202083
rect 675286 202031 675338 202083
rect 144022 201587 144074 201639
rect 197206 201587 197258 201639
rect 40246 201513 40298 201565
rect 41782 201513 41834 201565
rect 40054 201439 40106 201491
rect 42166 201439 42218 201491
rect 674038 201291 674090 201343
rect 675382 201291 675434 201343
rect 41974 201069 42026 201121
rect 42358 201069 42410 201121
rect 674902 200847 674954 200899
rect 675382 200847 675434 200899
rect 144118 198849 144170 198901
rect 188566 198849 188618 198901
rect 37366 198775 37418 198827
rect 43222 198775 43274 198827
rect 144022 198775 144074 198827
rect 191446 198775 191498 198827
rect 40150 198701 40202 198753
rect 40918 198701 40970 198753
rect 146230 198701 146282 198753
rect 194326 198701 194378 198753
rect 674806 197591 674858 197643
rect 675382 197591 675434 197643
rect 42070 197443 42122 197495
rect 42934 197443 42986 197495
rect 41782 197369 41834 197421
rect 41782 197147 41834 197199
rect 674614 196999 674666 197051
rect 675478 196999 675530 197051
rect 674710 196555 674762 196607
rect 675382 196555 675434 196607
rect 144022 195815 144074 195867
rect 185686 195815 185738 195867
rect 42550 195741 42602 195793
rect 42838 195741 42890 195793
rect 42838 195593 42890 195645
rect 43222 195593 43274 195645
rect 42166 195297 42218 195349
rect 42358 195297 42410 195349
rect 42070 194483 42122 194535
rect 50422 194483 50474 194535
rect 42070 193447 42122 193499
rect 43030 193447 43082 193499
rect 42166 192189 42218 192241
rect 43126 192189 43178 192241
rect 42070 191449 42122 191501
rect 42358 191449 42410 191501
rect 144022 190117 144074 190169
rect 151222 190117 151274 190169
rect 204886 190117 204938 190169
rect 205078 190117 205130 190169
rect 42166 187675 42218 187727
rect 42838 187675 42890 187727
rect 42262 187157 42314 187209
rect 42934 187231 42986 187283
rect 146422 187231 146474 187283
rect 197302 187231 197354 187283
rect 204886 187157 204938 187209
rect 205078 187157 205130 187209
rect 206998 187157 207050 187209
rect 207286 187157 207338 187209
rect 42166 187083 42218 187135
rect 42550 187083 42602 187135
rect 144502 184419 144554 184471
rect 148534 184419 148586 184471
rect 146806 184345 146858 184397
rect 194422 184345 194474 184397
rect 655318 184345 655370 184397
rect 674422 184345 674474 184397
rect 660982 183901 661034 183953
rect 674710 183901 674762 183953
rect 666742 182865 666794 182917
rect 674422 182865 674474 182917
rect 146806 181459 146858 181511
rect 188662 181459 188714 181511
rect 145270 178647 145322 178699
rect 148630 178647 148682 178699
rect 146806 178573 146858 178625
rect 191542 178573 191594 178625
rect 146806 175687 146858 175739
rect 185782 175687 185834 175739
rect 144022 175613 144074 175665
rect 146518 175613 146570 175665
rect 146806 172801 146858 172853
rect 162742 172801 162794 172853
rect 146806 171247 146858 171299
rect 159862 171247 159914 171299
rect 146806 167251 146858 167303
rect 156982 167251 157034 167303
rect 647062 167177 647114 167229
rect 674710 167177 674762 167229
rect 144022 166659 144074 166711
rect 146518 166659 146570 166711
rect 646294 164217 646346 164269
rect 674614 164217 674666 164269
rect 144022 164143 144074 164195
rect 208726 164143 208778 164195
rect 647926 164143 647978 164195
rect 674710 164143 674762 164195
rect 144694 163699 144746 163751
rect 146806 163699 146858 163751
rect 674710 163625 674762 163677
rect 677110 163625 677162 163677
rect 674806 163255 674858 163307
rect 676822 163255 676874 163307
rect 206998 162885 207050 162937
rect 207382 162885 207434 162937
rect 144022 161257 144074 161309
rect 148726 161257 148778 161309
rect 674902 160739 674954 160791
rect 675382 160739 675434 160791
rect 674998 159999 675050 160051
rect 675478 159999 675530 160051
rect 144022 158445 144074 158497
rect 148822 158445 148874 158497
rect 674518 157705 674570 157757
rect 675190 157705 675242 157757
rect 674614 156891 674666 156943
rect 675478 156891 675530 156943
rect 144022 155707 144074 155759
rect 148918 155707 148970 155759
rect 144118 155633 144170 155685
rect 200182 155633 200234 155685
rect 144214 155559 144266 155611
rect 203062 155559 203114 155611
rect 144022 152747 144074 152799
rect 180022 152747 180074 152799
rect 144118 152673 144170 152725
rect 182902 152673 182954 152725
rect 674230 152599 674282 152651
rect 675382 152599 675434 152651
rect 674806 152155 674858 152207
rect 675478 152155 675530 152207
rect 674134 151415 674186 151467
rect 675382 151415 675434 151467
rect 674710 150305 674762 150357
rect 675478 150305 675530 150357
rect 144118 149861 144170 149913
rect 149014 149861 149066 149913
rect 144022 149787 144074 149839
rect 177238 149787 177290 149839
rect 144022 149639 144074 149691
rect 144502 149639 144554 149691
rect 144694 147197 144746 147249
rect 144022 147123 144074 147175
rect 144694 147049 144746 147101
rect 144118 146901 144170 146953
rect 144502 146901 144554 146953
rect 174358 146901 174410 146953
rect 144502 146235 144554 146287
rect 146326 146235 146378 146287
rect 144214 146087 144266 146139
rect 146326 146087 146378 146139
rect 144214 144311 144266 144363
rect 154102 144311 154154 144363
rect 144214 144015 144266 144067
rect 208822 144015 208874 144067
rect 144214 142535 144266 142587
rect 149206 142535 149258 142587
rect 144214 141129 144266 141181
rect 171478 141129 171530 141181
rect 144214 140833 144266 140885
rect 144502 140833 144554 140885
rect 655222 138539 655274 138591
rect 674710 138539 674762 138591
rect 655126 138391 655178 138443
rect 674422 138391 674474 138443
rect 144502 138317 144554 138369
rect 168598 138317 168650 138369
rect 143830 138243 143882 138295
rect 208918 138243 208970 138295
rect 143926 138169 143978 138221
rect 144502 138169 144554 138221
rect 144694 136911 144746 136963
rect 144790 136689 144842 136741
rect 146902 136245 146954 136297
rect 149302 136245 149354 136297
rect 146902 135949 146954 136001
rect 149398 135949 149450 136001
rect 655414 135579 655466 135631
rect 674614 135579 674666 135631
rect 646486 135357 646538 135409
rect 674710 135357 674762 135409
rect 144214 134839 144266 134891
rect 146998 134839 147050 134891
rect 146710 134543 146762 134595
rect 146806 134321 146858 134373
rect 144214 134173 144266 134225
rect 146806 134173 146858 134225
rect 144502 132915 144554 132967
rect 144214 132693 144266 132745
rect 209110 132693 209162 132745
rect 146806 132619 146858 132671
rect 165718 132619 165770 132671
rect 144214 132545 144266 132597
rect 144502 132545 144554 132597
rect 209014 132545 209066 132597
rect 143926 130103 143978 130155
rect 144214 130103 144266 130155
rect 144502 129659 144554 129711
rect 151414 129659 151466 129711
rect 144214 129585 144266 129637
rect 209206 129585 209258 129637
rect 144502 129511 144554 129563
rect 146326 129511 146378 129563
rect 147094 126847 147146 126899
rect 149494 126847 149546 126899
rect 146710 126773 146762 126825
rect 203158 126773 203210 126825
rect 143926 126699 143978 126751
rect 144214 126699 144266 126751
rect 146326 126699 146378 126751
rect 208630 126699 208682 126751
rect 204790 126625 204842 126677
rect 204886 126625 204938 126677
rect 39862 125293 39914 125345
rect 42454 125293 42506 125345
rect 146710 124035 146762 124087
rect 197398 124035 197450 124087
rect 146326 123887 146378 123939
rect 200278 123887 200330 123939
rect 146326 123739 146378 123791
rect 146902 123739 146954 123791
rect 647830 121223 647882 121275
rect 674710 121223 674762 121275
rect 647734 121149 647786 121201
rect 674422 121149 674474 121201
rect 146902 121075 146954 121127
rect 149590 121075 149642 121127
rect 647926 121075 647978 121127
rect 674614 121075 674666 121127
rect 146710 121001 146762 121053
rect 208534 121001 208586 121053
rect 146326 119151 146378 119203
rect 146710 118559 146762 118611
rect 194518 118559 194570 118611
rect 146710 118263 146762 118315
rect 188758 118263 188810 118315
rect 146326 118115 146378 118167
rect 208438 118115 208490 118167
rect 674806 118041 674858 118093
rect 676822 118041 676874 118093
rect 146326 117967 146378 118019
rect 674710 117967 674762 118019
rect 676918 117967 676970 118019
rect 675478 115747 675530 115799
rect 146902 115525 146954 115577
rect 149686 115525 149738 115577
rect 675478 115525 675530 115577
rect 146710 115229 146762 115281
rect 208342 115229 208394 115281
rect 143830 115155 143882 115207
rect 144310 115155 144362 115207
rect 144406 115155 144458 115207
rect 144502 115155 144554 115207
rect 143734 115081 143786 115133
rect 144118 115081 144170 115133
rect 144118 114933 144170 114985
rect 146326 115155 146378 115207
rect 146326 115007 146378 115059
rect 146998 115007 147050 115059
rect 144502 114933 144554 114985
rect 144598 114933 144650 114985
rect 674614 114785 674666 114837
rect 675382 114785 675434 114837
rect 146710 112639 146762 112691
rect 191638 112639 191690 112691
rect 144406 112417 144458 112469
rect 148150 112417 148202 112469
rect 146710 112343 146762 112395
rect 148054 112343 148106 112395
rect 207190 112343 207242 112395
rect 207382 112343 207434 112395
rect 674518 110937 674570 110989
rect 675094 110937 675146 110989
rect 144406 109531 144458 109583
rect 147958 109531 148010 109583
rect 146710 109457 146762 109509
rect 185878 109457 185930 109509
rect 674326 107311 674378 107363
rect 675382 107311 675434 107363
rect 674806 106941 674858 106993
rect 675478 106941 675530 106993
rect 144406 106645 144458 106697
rect 147862 106645 147914 106697
rect 146710 106571 146762 106623
rect 162838 106571 162890 106623
rect 204790 106571 204842 106623
rect 204982 106571 205034 106623
rect 143830 106497 143882 106549
rect 146710 106423 146762 106475
rect 674134 106127 674186 106179
rect 675382 106127 675434 106179
rect 674710 105165 674762 105217
rect 675382 105165 675434 105217
rect 144022 104869 144074 104921
rect 146518 104795 146570 104847
rect 146902 104795 146954 104847
rect 146518 104647 146570 104699
rect 647926 104499 647978 104551
rect 665206 104499 665258 104551
rect 144790 104203 144842 104255
rect 159958 104203 160010 104255
rect 144310 103759 144362 103811
rect 151318 103759 151370 103811
rect 144118 103685 144170 103737
rect 208246 103685 208298 103737
rect 146902 103611 146954 103663
rect 206710 103611 206762 103663
rect 146326 103537 146378 103589
rect 204502 103537 204554 103589
rect 144598 103463 144650 103515
rect 206230 103463 206282 103515
rect 143734 103315 143786 103367
rect 144598 103315 144650 103367
rect 144022 101539 144074 101591
rect 157078 101539 157130 101591
rect 144118 100799 144170 100851
rect 147766 100799 147818 100851
rect 146710 100725 146762 100777
rect 204694 100725 204746 100777
rect 144022 100651 144074 100703
rect 206902 100651 206954 100703
rect 144406 100577 144458 100629
rect 204598 100577 204650 100629
rect 151126 100503 151178 100555
rect 204502 100503 204554 100555
rect 191446 100429 191498 100481
rect 204790 100429 204842 100481
rect 143926 99985 143978 100037
rect 144310 99985 144362 100037
rect 640726 99319 640778 99371
rect 668182 99319 668234 99371
rect 144022 98061 144074 98113
rect 180118 98061 180170 98113
rect 144118 97987 144170 98039
rect 182998 97987 183050 98039
rect 144310 97913 144362 97965
rect 208150 97913 208202 97965
rect 154006 97839 154058 97891
rect 206518 97839 206570 97891
rect 156886 97765 156938 97817
rect 204502 97765 204554 97817
rect 174262 97691 174314 97743
rect 205270 97691 205322 97743
rect 177142 97617 177194 97669
rect 206134 97617 206186 97669
rect 182806 97543 182858 97595
rect 204502 97543 204554 97595
rect 144022 95101 144074 95153
rect 174454 95101 174506 95153
rect 144118 95027 144170 95079
rect 177334 95027 177386 95079
rect 146518 94953 146570 95005
rect 206326 94953 206378 95005
rect 144598 94879 144650 94931
rect 206902 94879 206954 94931
rect 151222 94805 151274 94857
rect 204598 94805 204650 94857
rect 165622 94731 165674 94783
rect 205846 94731 205898 94783
rect 168502 94657 168554 94709
rect 205750 94657 205802 94709
rect 171382 94583 171434 94635
rect 204502 94583 204554 94635
rect 647350 92733 647402 92785
rect 660694 92733 660746 92785
rect 646678 92659 646730 92711
rect 659830 92659 659882 92711
rect 647542 92585 647594 92637
rect 661750 92585 661802 92637
rect 647254 92437 647306 92489
rect 659734 92437 659786 92489
rect 647830 92363 647882 92415
rect 663094 92363 663146 92415
rect 647734 92289 647786 92341
rect 662518 92289 662570 92341
rect 144118 92215 144170 92267
rect 154006 92215 154058 92267
rect 646198 92215 646250 92267
rect 661174 92215 661226 92267
rect 144022 92141 144074 92193
rect 171574 92141 171626 92193
rect 646582 92141 646634 92193
rect 658870 92141 658922 92193
rect 203062 92067 203114 92119
rect 204598 92067 204650 92119
rect 200182 91993 200234 92045
rect 204502 91993 204554 92045
rect 197302 91919 197354 91971
rect 204694 91919 204746 91971
rect 194422 91845 194474 91897
rect 204598 91845 204650 91897
rect 188662 91771 188714 91823
rect 204790 91771 204842 91823
rect 144022 89403 144074 89455
rect 151222 89403 151274 89455
rect 144310 89329 144362 89381
rect 165622 89329 165674 89381
rect 204982 89329 205034 89381
rect 144118 89255 144170 89307
rect 168502 89255 168554 89307
rect 205078 89255 205130 89307
rect 156982 89181 157034 89233
rect 204694 89181 204746 89233
rect 206998 89181 207050 89233
rect 207190 89181 207242 89233
rect 159862 89107 159914 89159
rect 205270 89107 205322 89159
rect 162742 89033 162794 89085
rect 204598 89033 204650 89085
rect 185782 88959 185834 89011
rect 204502 88959 204554 89011
rect 191542 88885 191594 88937
rect 204790 88885 204842 88937
rect 646870 87997 646922 88049
rect 650902 87997 650954 88049
rect 658006 87257 658058 87309
rect 657046 87109 657098 87161
rect 647926 87035 647978 87087
rect 663286 87035 663338 87087
rect 144502 86443 144554 86495
rect 647926 86443 647978 86495
rect 651094 86443 651146 86495
rect 154102 86369 154154 86421
rect 204694 86369 204746 86421
rect 144502 86295 144554 86347
rect 174358 86295 174410 86347
rect 206614 86295 206666 86347
rect 177238 86221 177290 86273
rect 204598 86221 204650 86273
rect 180022 86147 180074 86199
rect 205558 86147 205610 86199
rect 182902 86073 182954 86125
rect 204502 86073 204554 86125
rect 646870 85111 646922 85163
rect 650998 85111 651050 85163
rect 146710 84963 146762 85015
rect 204502 84963 204554 85015
rect 151414 83483 151466 83535
rect 206230 83483 206282 83535
rect 165718 83409 165770 83461
rect 206710 83409 206762 83461
rect 647926 83409 647978 83461
rect 657046 83409 657098 83461
rect 168598 83335 168650 83387
rect 205750 83335 205802 83387
rect 171478 83261 171530 83313
rect 204502 83261 204554 83313
rect 146710 82077 146762 82129
rect 204502 82077 204554 82129
rect 647926 81855 647978 81907
rect 663286 81855 663338 81907
rect 645910 81781 645962 81833
rect 663382 81781 663434 81833
rect 647638 81633 647690 81685
rect 661078 81633 661130 81685
rect 647926 81263 647978 81315
rect 657526 81263 657578 81315
rect 143926 80671 143978 80723
rect 144694 80671 144746 80723
rect 659446 80671 659498 80723
rect 659542 80671 659594 80723
rect 203158 80597 203210 80649
rect 205270 80597 205322 80649
rect 200278 80523 200330 80575
rect 204502 80523 204554 80575
rect 197398 80449 197450 80501
rect 204598 80449 204650 80501
rect 194518 80375 194570 80427
rect 204694 80375 204746 80427
rect 188758 80301 188810 80353
rect 210166 80301 210218 80353
rect 647926 80153 647978 80205
rect 656950 80153 657002 80205
rect 645430 79635 645482 79687
rect 651190 79635 651242 79687
rect 647734 79265 647786 79317
rect 658870 79265 658922 79317
rect 647830 78821 647882 78873
rect 660694 78821 660746 78873
rect 647926 78303 647978 78355
rect 662518 78303 662570 78355
rect 144310 77859 144362 77911
rect 151126 77859 151178 77911
rect 146710 77785 146762 77837
rect 146614 77711 146666 77763
rect 157078 77711 157130 77763
rect 189910 77711 189962 77763
rect 204598 77711 204650 77763
rect 647446 77711 647498 77763
rect 659446 77711 659498 77763
rect 159958 77637 160010 77689
rect 206518 77637 206570 77689
rect 647926 77637 647978 77689
rect 650998 77637 651050 77689
rect 162838 77563 162890 77615
rect 204502 77563 204554 77615
rect 185878 77489 185930 77541
rect 205942 77489 205994 77541
rect 146614 77415 146666 77467
rect 189910 77415 189962 77467
rect 204694 77415 204746 77467
rect 191638 77341 191690 77393
rect 204790 77341 204842 77393
rect 647926 77267 647978 77319
rect 662902 77267 662954 77319
rect 646486 76897 646538 76949
rect 658294 76897 658346 76949
rect 646486 76749 646538 76801
rect 650902 76749 650954 76801
rect 646102 75787 646154 75839
rect 661750 75787 661802 75839
rect 646486 75417 646538 75469
rect 656854 75417 656906 75469
rect 146518 75047 146570 75099
rect 160150 75047 160202 75099
rect 144022 74973 144074 75025
rect 156982 74973 157034 75025
rect 144310 74899 144362 74951
rect 161494 74899 161546 74951
rect 154006 74825 154058 74877
rect 204694 74825 204746 74877
rect 174454 74751 174506 74803
rect 206806 74751 206858 74803
rect 177334 74677 177386 74729
rect 204598 74677 204650 74729
rect 180118 74603 180170 74655
rect 205750 74603 205802 74655
rect 182998 74529 183050 74581
rect 204502 74529 204554 74581
rect 144310 74159 144362 74211
rect 145462 74159 145514 74211
rect 144118 74085 144170 74137
rect 148342 74085 148394 74137
rect 145462 74011 145514 74063
rect 146038 74011 146090 74063
rect 647254 72531 647306 72583
rect 663190 72531 663242 72583
rect 646870 72457 646922 72509
rect 660118 72457 660170 72509
rect 646102 72235 646154 72287
rect 663382 72235 663434 72287
rect 146038 72013 146090 72065
rect 154678 72013 154730 72065
rect 151222 71939 151274 71991
rect 206806 71939 206858 71991
rect 161494 71865 161546 71917
rect 204982 71865 205034 71917
rect 165622 71791 165674 71843
rect 205462 71791 205514 71843
rect 168502 71717 168554 71769
rect 204598 71717 204650 71769
rect 171574 71643 171626 71695
rect 204502 71643 204554 71695
rect 144022 70237 144074 70289
rect 149782 70237 149834 70289
rect 146038 69201 146090 69253
rect 146326 69201 146378 69253
rect 144022 69127 144074 69179
rect 206998 69127 207050 69179
rect 207286 69127 207338 69179
rect 206518 69053 206570 69105
rect 149782 68979 149834 69031
rect 204118 68979 204170 69031
rect 205174 68979 205226 69031
rect 207478 68979 207530 69031
rect 154678 68905 154730 68957
rect 204598 68905 204650 68957
rect 156982 68831 157034 68883
rect 206422 68831 206474 68883
rect 160150 68757 160202 68809
rect 204502 68757 204554 68809
rect 144118 67203 144170 67255
rect 152662 67203 152714 67255
rect 146326 66389 146378 66441
rect 158326 66389 158378 66441
rect 146806 66241 146858 66293
rect 144022 66167 144074 66219
rect 144694 66167 144746 66219
rect 205462 66167 205514 66219
rect 152662 66093 152714 66145
rect 206326 66093 206378 66145
rect 158326 66019 158378 66071
rect 204502 66019 204554 66071
rect 145462 65871 145514 65923
rect 146326 65871 146378 65923
rect 145078 65723 145130 65775
rect 145462 65723 145514 65775
rect 144118 64983 144170 65035
rect 144310 64983 144362 65035
rect 144310 64835 144362 64887
rect 204598 64835 204650 64887
rect 144982 64761 145034 64813
rect 204502 64761 204554 64813
rect 146902 63355 146954 63407
rect 204502 63355 204554 63407
rect 144022 62911 144074 62963
rect 144310 62911 144362 62963
rect 144022 62467 144074 62519
rect 149782 62467 149834 62519
rect 160534 60765 160586 60817
rect 204598 60765 204650 60817
rect 156310 60691 156362 60743
rect 204694 60691 204746 60743
rect 152662 60617 152714 60669
rect 204502 60617 204554 60669
rect 151222 60543 151274 60595
rect 204886 60543 204938 60595
rect 148342 60469 148394 60521
rect 204790 60469 204842 60521
rect 146902 60395 146954 60447
rect 206806 60395 206858 60447
rect 149782 60321 149834 60373
rect 204598 60321 204650 60373
rect 207766 60321 207818 60373
rect 208726 60321 208778 60373
rect 207862 60247 207914 60299
rect 208822 60247 208874 60299
rect 208822 59951 208874 60003
rect 209110 59951 209162 60003
rect 209494 59951 209546 60003
rect 209974 59951 210026 60003
rect 144022 59581 144074 59633
rect 160534 59581 160586 59633
rect 144022 58989 144074 59041
rect 204502 58989 204554 59041
rect 144022 57065 144074 57117
rect 156310 57065 156362 57117
rect 144022 56473 144074 56525
rect 152662 56473 152714 56525
rect 209974 54845 210026 54897
rect 144022 54623 144074 54675
rect 151222 54623 151274 54675
rect 210166 54253 210218 54305
rect 218998 54253 219050 54305
rect 221014 54253 221066 54305
rect 207478 54179 207530 54231
rect 216310 54179 216362 54231
rect 144022 54105 144074 54157
rect 148342 54105 148394 54157
rect 210070 54105 210122 54157
rect 219190 54105 219242 54157
rect 209206 54031 209258 54083
rect 218998 54031 219050 54083
rect 209302 53957 209354 54009
rect 218806 53957 218858 54009
rect 208438 53883 208490 53935
rect 219190 53883 219242 53935
rect 208054 53809 208106 53861
rect 216790 53809 216842 53861
rect 212374 53735 212426 53787
rect 221206 53735 221258 53787
rect 210262 53661 210314 53713
rect 293782 53661 293834 53713
rect 209974 53587 210026 53639
rect 330934 53587 330986 53639
rect 211558 53513 211610 53565
rect 216598 53513 216650 53565
rect 219190 53513 219242 53565
rect 219814 53513 219866 53565
rect 221014 53513 221066 53565
rect 403126 53513 403178 53565
rect 210358 53439 210410 53491
rect 217798 53439 217850 53491
rect 218998 53439 219050 53491
rect 452182 53439 452234 53491
rect 209590 53365 209642 53417
rect 217462 53365 217514 53417
rect 218806 53365 218858 53417
rect 466486 53365 466538 53417
rect 209398 53291 209450 53343
rect 219670 53291 219722 53343
rect 219862 53291 219914 53343
rect 517846 53291 517898 53343
rect 207190 53217 207242 53269
rect 215542 53217 215594 53269
rect 209782 53143 209834 53195
rect 213334 53143 213386 53195
rect 208150 53069 208202 53121
rect 215734 53069 215786 53121
rect 216022 53069 216074 53121
rect 308086 53217 308138 53269
rect 308182 53143 308234 53195
rect 348406 53217 348458 53269
rect 348502 53143 348554 53195
rect 207958 52995 208010 53047
rect 218134 52995 218186 53047
rect 420502 53217 420554 53269
rect 443542 53217 443594 53269
rect 463702 53217 463754 53269
rect 483862 53217 483914 53269
rect 463606 53143 463658 53195
rect 420598 53069 420650 53121
rect 443446 53069 443498 53121
rect 483862 52995 483914 53047
rect 514006 52995 514058 53047
rect 207286 52847 207338 52899
rect 219862 52847 219914 52899
rect 212182 52625 212234 52677
rect 220918 52625 220970 52677
rect 151318 52551 151370 52603
rect 217270 52551 217322 52603
rect 151126 52403 151178 52455
rect 216118 52403 216170 52455
rect 211222 52329 211274 52381
rect 227446 52329 227498 52381
rect 137494 52255 137546 52307
rect 221782 52255 221834 52307
rect 146710 52107 146762 52159
rect 161302 52107 161354 52159
rect 181366 52107 181418 52159
rect 227158 52181 227210 52233
rect 144406 52033 144458 52085
rect 212182 52033 212234 52085
rect 144598 51959 144650 52011
rect 225718 52107 225770 52159
rect 212374 52033 212426 52085
rect 213430 52033 213482 52085
rect 146518 51885 146570 51937
rect 227542 51885 227594 51937
rect 423382 51885 423434 51937
rect 432790 51885 432842 51937
rect 483862 51885 483914 51937
rect 493846 51885 493898 51937
rect 544342 51885 544394 51937
rect 552790 51885 552842 51937
rect 625750 51885 625802 51937
rect 639670 51885 639722 51937
rect 213430 51811 213482 51863
rect 645526 51811 645578 51863
rect 209686 51737 209738 51789
rect 213718 51737 213770 51789
rect 216598 51737 216650 51789
rect 645718 51737 645770 51789
rect 209878 51663 209930 51715
rect 214102 51663 214154 51715
rect 221782 51589 221834 51641
rect 243862 51589 243914 51641
rect 145366 51515 145418 51567
rect 237622 51515 237674 51567
rect 145558 51441 145610 51493
rect 236374 51441 236426 51493
rect 145942 51367 145994 51419
rect 237142 51367 237194 51419
rect 287926 51663 287978 51715
rect 288022 51663 288074 51715
rect 292054 51663 292106 51715
rect 292054 51515 292106 51567
rect 302422 51515 302474 51567
rect 302518 51515 302570 51567
rect 322582 51515 322634 51567
rect 144310 51293 144362 51345
rect 145654 51219 145706 51271
rect 227446 51293 227498 51345
rect 145750 51145 145802 51197
rect 217270 51145 217322 51197
rect 233782 51219 233834 51271
rect 322582 51367 322634 51419
rect 348406 51663 348458 51715
rect 403318 51663 403370 51715
rect 423382 51663 423434 51715
rect 469558 51663 469610 51715
rect 483862 51663 483914 51715
rect 330934 51589 330986 51641
rect 348310 51589 348362 51641
rect 348502 51589 348554 51641
rect 372022 51589 372074 51641
rect 372118 51515 372170 51567
rect 432790 51589 432842 51641
rect 452662 51589 452714 51641
rect 403126 51515 403178 51567
rect 452758 51515 452810 51567
rect 469366 51589 469418 51641
rect 493846 51515 493898 51567
rect 552790 51663 552842 51715
rect 544342 51589 544394 51641
rect 610486 51663 610538 51715
rect 610678 51589 610730 51641
rect 625750 51589 625802 51641
rect 235414 51145 235466 51197
rect 146134 51071 146186 51123
rect 232342 51071 232394 51123
rect 146230 50997 146282 51049
rect 232726 50997 232778 51049
rect 146422 50923 146474 50975
rect 231958 50923 232010 50975
rect 146614 50849 146666 50901
rect 230998 50849 231050 50901
rect 146806 50775 146858 50827
rect 230614 50775 230666 50827
rect 144886 50701 144938 50753
rect 228790 50701 228842 50753
rect 145078 50627 145130 50679
rect 228310 50627 228362 50679
rect 145270 50553 145322 50605
rect 229750 50553 229802 50605
rect 145174 50479 145226 50531
rect 229366 50479 229418 50531
rect 145462 50405 145514 50457
rect 228406 50405 228458 50457
rect 144502 50331 144554 50383
rect 208150 50331 208202 50383
rect 208246 50331 208298 50383
rect 216886 50331 216938 50383
rect 146038 50257 146090 50309
rect 207958 50257 208010 50309
rect 144214 50183 144266 50235
rect 224278 50257 224330 50309
rect 217270 50183 217322 50235
rect 235990 50183 236042 50235
rect 144982 50109 145034 50161
rect 234550 50109 234602 50161
rect 145846 50035 145898 50087
rect 234934 50035 234986 50087
rect 144118 49961 144170 50013
rect 237238 49961 237290 50013
rect 146326 49887 146378 49939
rect 232822 49887 232874 49939
rect 209110 49813 209162 49865
rect 221494 49813 221546 49865
rect 208150 49739 208202 49791
rect 225334 49739 225386 49791
rect 207958 49665 208010 49717
rect 226582 49665 226634 49717
rect 208342 49591 208394 49643
rect 219478 49591 219530 49643
rect 223702 48925 223754 48977
rect 229654 48925 229706 48977
rect 208534 48851 208586 48903
rect 220534 48851 220586 48903
rect 222934 48851 222986 48903
rect 645334 48851 645386 48903
rect 209014 48777 209066 48829
rect 222070 48777 222122 48829
rect 222262 48777 222314 48829
rect 645238 48777 645290 48829
rect 208630 48703 208682 48755
rect 221686 48703 221738 48755
rect 224086 48703 224138 48755
rect 645142 48703 645194 48755
rect 208918 48629 208970 48681
rect 222358 48629 222410 48681
rect 148438 48555 148490 48607
rect 235030 48555 235082 48607
rect 208822 48481 208874 48533
rect 222742 48481 222794 48533
rect 188566 48407 188618 48459
rect 241174 48407 241226 48459
rect 208726 48333 208778 48385
rect 223894 48333 223946 48385
rect 197206 48259 197258 48311
rect 241558 48259 241610 48311
rect 149110 48185 149162 48237
rect 226102 48185 226154 48237
rect 149206 48111 149258 48163
rect 224566 48111 224618 48163
rect 149398 48037 149450 48089
rect 223126 48037 223178 48089
rect 149302 47963 149354 48015
rect 223510 47963 223562 48015
rect 149590 47889 149642 47941
rect 220150 47889 220202 47941
rect 149494 47815 149546 47867
rect 221302 47815 221354 47867
rect 149686 47741 149738 47793
rect 219094 47741 219146 47793
rect 147766 47667 147818 47719
rect 216502 47667 216554 47719
rect 147862 47593 147914 47645
rect 217654 47593 217706 47645
rect 147958 47519 148010 47571
rect 217942 47519 217994 47571
rect 514006 47519 514058 47571
rect 525910 47519 525962 47571
rect 148054 47445 148106 47497
rect 218326 47445 218378 47497
rect 148150 47371 148202 47423
rect 218710 47371 218762 47423
rect 179926 47297 179978 47349
rect 238582 47297 238634 47349
rect 185686 47223 185738 47275
rect 240406 47223 240458 47275
rect 202966 47149 203018 47201
rect 239350 47149 239402 47201
rect 148822 47075 148874 47127
rect 233302 47075 233354 47127
rect 200086 47001 200138 47053
rect 238966 47001 239018 47053
rect 194326 46927 194378 46979
rect 240790 46927 240842 46979
rect 148918 46853 148970 46905
rect 230134 46853 230186 46905
rect 148534 46779 148586 46831
rect 231574 46779 231626 46831
rect 207862 46705 207914 46757
rect 224950 46705 225002 46757
rect 225046 46705 225098 46757
rect 227926 46705 227978 46757
rect 149014 46631 149066 46683
rect 226486 46631 226538 46683
rect 148726 46557 148778 46609
rect 234166 46557 234218 46609
rect 148630 46483 148682 46535
rect 230518 46483 230570 46535
rect 218518 46409 218570 46461
rect 645622 46409 645674 46461
rect 159766 46335 159818 46387
rect 239446 46335 239498 46387
rect 207766 46261 207818 46313
rect 225046 46261 225098 46313
rect 148246 46187 148298 46239
rect 236758 46187 236810 46239
rect 162646 46113 162698 46165
rect 239830 46113 239882 46165
rect 293782 45817 293834 45869
rect 302326 45817 302378 45869
rect 211702 45299 211754 45351
rect 327286 45299 327338 45351
rect 211414 45225 211466 45277
rect 328054 45225 328106 45277
rect 213910 45151 213962 45203
rect 446902 45151 446954 45203
rect 214678 45077 214730 45129
rect 506806 45077 506858 45129
rect 215062 45003 215114 45055
rect 506710 45003 506762 45055
rect 215446 44929 215498 44981
rect 526966 44929 527018 44981
rect 452182 43523 452234 43575
rect 461110 43523 461162 43575
rect 213238 43227 213290 43279
rect 410998 43227 411050 43279
rect 446902 43153 446954 43205
rect 454966 43153 455018 43205
rect 348310 42857 348362 42909
rect 357430 42857 357482 42909
rect 133654 42783 133706 42835
rect 136534 42783 136586 42835
rect 212470 42339 212522 42391
rect 310102 42339 310154 42391
rect 206902 42117 206954 42169
rect 405238 42117 405290 42169
rect 213622 42043 213674 42095
rect 460054 42043 460106 42095
rect 214294 41969 214346 42021
rect 514870 41969 514922 42021
rect 506806 41895 506858 41947
rect 521590 41969 521642 42021
rect 403414 41821 403466 41873
rect 506710 41747 506762 41799
rect 518518 41747 518570 41799
<< metal2 >>
rect 93910 1010977 93962 1010983
rect 93910 1010919 93962 1010925
rect 97078 1010977 97130 1010983
rect 97078 1010919 97130 1010925
rect 93718 1005575 93770 1005581
rect 93718 1005517 93770 1005523
rect 92566 1005427 92618 1005433
rect 92566 1005369 92618 1005375
rect 92470 1005205 92522 1005211
rect 92470 1005147 92522 1005153
rect 92374 1003725 92426 1003731
rect 92374 1003667 92426 1003673
rect 87860 995846 87916 995855
rect 81408 995813 81662 995832
rect 81408 995807 81674 995813
rect 81408 995804 81622 995807
rect 87552 995804 87860 995832
rect 88752 995813 89054 995832
rect 91248 995813 91550 995832
rect 88752 995807 89066 995813
rect 88752 995804 89014 995807
rect 87860 995781 87916 995790
rect 81622 995749 81674 995755
rect 91248 995807 91562 995813
rect 91248 995804 91510 995807
rect 89014 995749 89066 995755
rect 91510 995749 91562 995755
rect 92386 995739 92414 1003667
rect 92482 995813 92510 1005147
rect 92578 995855 92606 1005369
rect 92662 1005353 92714 1005359
rect 92662 1005295 92714 1005301
rect 92564 995846 92620 995855
rect 92470 995807 92522 995813
rect 92564 995781 92620 995790
rect 92470 995749 92522 995755
rect 89782 995733 89834 995739
rect 85940 995698 85996 995707
rect 85728 995656 85940 995684
rect 89424 995681 89782 995684
rect 89424 995675 89834 995681
rect 92374 995733 92426 995739
rect 92674 995707 92702 1005295
rect 92950 1005279 93002 1005285
rect 92950 1005221 93002 1005227
rect 92758 999507 92810 999513
rect 92758 999449 92810 999455
rect 92374 995675 92426 995681
rect 92660 995698 92716 995707
rect 89424 995656 89822 995675
rect 85940 995633 85996 995642
rect 92660 995633 92716 995642
rect 86516 995550 86572 995559
rect 77088 995508 77342 995536
rect 69142 995141 69194 995147
rect 69142 995083 69194 995089
rect 61846 993883 61898 993889
rect 61846 993825 61898 993831
rect 47638 988333 47690 988339
rect 47638 988275 47690 988281
rect 44758 988259 44810 988265
rect 44758 988201 44810 988207
rect 43126 987889 43178 987895
rect 43126 987831 43178 987837
rect 41794 968771 41822 969252
rect 41780 968762 41836 968771
rect 41780 968697 41836 968706
rect 41794 967143 41822 967402
rect 43138 967323 43166 987831
rect 42166 967317 42218 967323
rect 42166 967259 42218 967265
rect 43126 967317 43178 967323
rect 43126 967259 43178 967265
rect 41780 967134 41836 967143
rect 41780 967069 41836 967078
rect 42178 966736 42206 967259
rect 41794 965071 41822 965552
rect 41780 965062 41836 965071
rect 41780 964997 41836 965006
rect 41794 964035 41822 964368
rect 41780 964026 41836 964035
rect 41780 963961 41836 963970
rect 41794 963295 41822 963702
rect 41780 963286 41836 963295
rect 41780 963221 41836 963230
rect 42178 962851 42206 963081
rect 42164 962842 42220 962851
rect 42164 962777 42220 962786
rect 42082 962259 42110 962518
rect 42068 962250 42124 962259
rect 42068 962185 42124 962194
rect 42164 962102 42220 962111
rect 42452 962102 42508 962111
rect 42220 962060 42302 962088
rect 42164 962037 42220 962046
rect 42178 961200 42206 961260
rect 42274 961200 42302 962060
rect 42452 962037 42508 962046
rect 42178 961172 42302 961200
rect 42466 961033 42494 962037
rect 42166 961027 42218 961033
rect 42166 960969 42218 960975
rect 42454 961027 42506 961033
rect 42454 960969 42506 960975
rect 42178 960594 42206 960969
rect 42178 959595 42206 960045
rect 42164 959586 42220 959595
rect 42164 959521 42220 959530
rect 41794 959151 41822 959410
rect 41780 959142 41836 959151
rect 41780 959077 41836 959086
rect 41986 958411 42014 958744
rect 41972 958402 42028 958411
rect 41972 958337 42028 958346
rect 42178 957819 42206 958226
rect 42164 957810 42220 957819
rect 42164 957745 42220 957754
rect 41780 956626 41836 956635
rect 41780 956561 41836 956570
rect 41794 956376 41822 956561
rect 42082 955261 42110 955710
rect 42070 955255 42122 955261
rect 42070 955197 42122 955203
rect 42838 955255 42890 955261
rect 42838 955197 42890 955203
rect 41794 954669 41822 955077
rect 41782 954663 41834 954669
rect 41782 954605 41834 954611
rect 41782 954441 41834 954447
rect 41782 954383 41834 954389
rect 41794 952227 41822 954383
rect 37366 952221 37418 952227
rect 37366 952163 37418 952169
rect 41782 952221 41834 952227
rect 41782 952163 41834 952169
rect 37378 942871 37406 952163
rect 42452 949374 42508 949383
rect 42452 949309 42508 949318
rect 42356 948486 42412 948495
rect 42356 948421 42358 948430
rect 42410 948421 42412 948430
rect 42358 948389 42410 948395
rect 42466 947491 42494 949309
rect 42646 947929 42698 947935
rect 42644 947894 42646 947903
rect 42698 947894 42700 947903
rect 42644 947829 42700 947838
rect 42454 947485 42506 947491
rect 42454 947427 42506 947433
rect 40628 946562 40684 946571
rect 40628 946497 40684 946506
rect 40244 945082 40300 945091
rect 40244 945017 40300 945026
rect 37364 942862 37420 942871
rect 37364 942797 37420 942806
rect 40258 927437 40286 945017
rect 40436 944934 40492 944943
rect 40436 944869 40492 944878
rect 40054 927431 40106 927437
rect 40054 927373 40106 927379
rect 40246 927431 40298 927437
rect 40246 927373 40298 927379
rect 40066 908216 40094 927373
rect 39970 908188 40094 908216
rect 39970 892879 39998 908188
rect 39958 892873 40010 892879
rect 39958 892815 40010 892821
rect 40150 892873 40202 892879
rect 40150 892815 40202 892821
rect 40162 877728 40190 892815
rect 40066 877700 40190 877728
rect 40066 864019 40094 877700
rect 40054 864013 40106 864019
rect 40054 863955 40106 863961
rect 40246 864013 40298 864019
rect 40246 863955 40298 863961
rect 40258 832421 40286 863955
rect 40246 832415 40298 832421
rect 40246 832357 40298 832363
rect 40054 832341 40106 832347
rect 40054 832283 40106 832289
rect 40066 826649 40094 832283
rect 40054 826643 40106 826649
rect 40054 826585 40106 826591
rect 40246 826643 40298 826649
rect 40246 826585 40298 826591
rect 40258 820031 40286 826585
rect 40244 820022 40300 820031
rect 40244 819957 40300 819966
rect 40450 819587 40478 944869
rect 40642 820771 40670 946497
rect 42850 939171 42878 955197
rect 42836 939162 42892 939171
rect 42836 939097 42892 939106
rect 42356 932502 42412 932511
rect 42356 932437 42412 932446
rect 42370 931031 42398 932437
rect 42356 931022 42412 931031
rect 42356 930957 42358 930966
rect 42410 930957 42412 930966
rect 44662 930983 44714 930989
rect 42358 930925 42410 930931
rect 44662 930925 44714 930931
rect 42166 823905 42218 823911
rect 42164 823870 42166 823879
rect 42218 823870 42220 823879
rect 42164 823805 42220 823814
rect 42166 823165 42218 823171
rect 42164 823130 42166 823139
rect 42218 823130 42220 823139
rect 42164 823065 42220 823074
rect 42166 822277 42218 822283
rect 42164 822242 42166 822251
rect 42218 822242 42220 822251
rect 42164 822177 42220 822186
rect 43220 821206 43276 821215
rect 43220 821141 43276 821150
rect 40628 820762 40684 820771
rect 40628 820697 40684 820706
rect 40436 819578 40492 819587
rect 40436 819513 40492 819522
rect 37268 819134 37324 819143
rect 37268 819069 37324 819078
rect 37282 802123 37310 819069
rect 41684 817950 41740 817959
rect 41684 817885 41740 817894
rect 40148 816766 40204 816775
rect 40148 816701 40204 816710
rect 37364 812770 37420 812779
rect 37364 812705 37420 812714
rect 37378 802271 37406 812705
rect 40162 803487 40190 816701
rect 40244 815878 40300 815887
rect 40244 815813 40300 815822
rect 40150 803481 40202 803487
rect 40150 803423 40202 803429
rect 37364 802262 37420 802271
rect 37364 802197 37420 802206
rect 37268 802114 37324 802123
rect 37268 802049 37324 802058
rect 40258 801975 40286 815813
rect 41492 811142 41548 811151
rect 41492 811077 41548 811086
rect 40244 801966 40300 801975
rect 40244 801901 40300 801910
rect 41506 800601 41534 811077
rect 41588 809218 41644 809227
rect 41588 809153 41644 809162
rect 41494 800595 41546 800601
rect 41494 800537 41546 800543
rect 41602 800527 41630 809153
rect 41590 800521 41642 800527
rect 41698 800495 41726 817885
rect 42836 815730 42892 815739
rect 42836 815665 42892 815674
rect 41876 813658 41932 813667
rect 41876 813593 41932 813602
rect 41780 809662 41836 809671
rect 41780 809597 41836 809606
rect 41590 800463 41642 800469
rect 41684 800486 41740 800495
rect 41684 800421 41740 800430
rect 41794 800347 41822 809597
rect 41780 800338 41836 800347
rect 41780 800273 41836 800282
rect 41890 800231 41918 813593
rect 41972 812326 42028 812335
rect 41972 812261 42028 812270
rect 41986 802081 42014 812261
rect 42166 810511 42218 810517
rect 42166 810453 42218 810459
rect 42068 808330 42124 808339
rect 42068 808265 42124 808274
rect 41974 802075 42026 802081
rect 41974 802017 42026 802023
rect 42082 800347 42110 808265
rect 42068 800338 42124 800347
rect 42068 800273 42124 800282
rect 42178 800231 42206 810453
rect 42850 807113 42878 815665
rect 43028 814990 43084 814999
rect 43028 814925 43084 814934
rect 43042 810517 43070 814925
rect 43030 810511 43082 810517
rect 43030 810453 43082 810459
rect 43028 810402 43084 810411
rect 43028 810337 43084 810346
rect 42454 807107 42506 807113
rect 42454 807049 42506 807055
rect 42838 807107 42890 807113
rect 42838 807049 42890 807055
rect 42466 802271 42494 807049
rect 42836 806998 42892 807007
rect 42836 806933 42892 806942
rect 42850 805527 42878 806933
rect 42836 805518 42892 805527
rect 42836 805453 42838 805462
rect 42890 805453 42892 805462
rect 42838 805421 42890 805427
rect 42838 803481 42890 803487
rect 42838 803423 42890 803429
rect 42452 802262 42508 802271
rect 42452 802197 42508 802206
rect 42454 802075 42506 802081
rect 42454 802017 42506 802023
rect 41878 800225 41930 800231
rect 41878 800167 41930 800173
rect 42166 800225 42218 800231
rect 42166 800167 42218 800173
rect 41878 800003 41930 800009
rect 41878 799945 41930 799951
rect 41890 799422 41918 799945
rect 42466 799755 42494 802017
rect 42452 799746 42508 799755
rect 42452 799681 42508 799690
rect 42850 798381 42878 803423
rect 43042 798529 43070 810337
rect 43124 807738 43180 807747
rect 43124 807673 43180 807682
rect 43030 798523 43082 798529
rect 43030 798465 43082 798471
rect 43028 798414 43084 798423
rect 42838 798375 42890 798381
rect 43028 798349 43084 798358
rect 42838 798317 42890 798323
rect 42166 798153 42218 798159
rect 42166 798095 42218 798101
rect 42178 797605 42206 798095
rect 42742 798079 42794 798085
rect 42742 798021 42794 798027
rect 42070 797339 42122 797345
rect 42070 797281 42122 797287
rect 42082 796980 42110 797281
rect 42754 796309 42782 798021
rect 42166 796303 42218 796309
rect 42166 796245 42218 796251
rect 42742 796303 42794 796309
rect 42742 796245 42794 796251
rect 42178 795765 42206 796245
rect 42742 796155 42794 796161
rect 42742 796097 42794 796103
rect 42166 795045 42218 795051
rect 42166 794987 42218 794993
rect 42178 794569 42206 794987
rect 41876 794270 41932 794279
rect 41876 794205 41932 794214
rect 41890 793946 41918 794205
rect 42068 793826 42124 793835
rect 42068 793761 42124 793770
rect 42082 793280 42110 793761
rect 42754 793053 42782 796097
rect 42166 793047 42218 793053
rect 42166 792989 42218 792995
rect 42742 793047 42794 793053
rect 42742 792989 42794 792995
rect 42178 792729 42206 792989
rect 42742 792899 42794 792905
rect 42742 792841 42794 792847
rect 42452 792494 42508 792503
rect 42452 792429 42508 792438
rect 42082 791171 42110 791430
rect 42068 791162 42124 791171
rect 42068 791097 42124 791106
rect 42164 791014 42220 791023
rect 42164 790949 42220 790958
rect 42178 790797 42206 790949
rect 42166 790679 42218 790685
rect 42166 790621 42218 790627
rect 42178 790246 42206 790621
rect 42166 789939 42218 789945
rect 42166 789881 42218 789887
rect 42178 789580 42206 789881
rect 42466 789501 42494 792429
rect 42754 790685 42782 792841
rect 43042 792355 43070 798349
rect 43138 795051 43166 807673
rect 43126 795045 43178 795051
rect 43126 794987 43178 794993
rect 43126 794897 43178 794903
rect 43126 794839 43178 794845
rect 43138 792905 43166 794839
rect 43126 792899 43178 792905
rect 43126 792841 43178 792847
rect 43028 792346 43084 792355
rect 43028 792281 43084 792290
rect 42836 791902 42892 791911
rect 42836 791837 42892 791846
rect 42742 790679 42794 790685
rect 42742 790621 42794 790627
rect 42740 790570 42796 790579
rect 42740 790505 42796 790514
rect 42166 789495 42218 789501
rect 42166 789437 42218 789443
rect 42454 789495 42506 789501
rect 42454 789437 42506 789443
rect 42178 788957 42206 789437
rect 42164 788646 42220 788655
rect 42164 788581 42220 788590
rect 42178 788396 42206 788581
rect 42166 787053 42218 787059
rect 42166 786995 42218 787001
rect 42178 786546 42206 786995
rect 42166 786461 42218 786467
rect 42166 786403 42218 786409
rect 42178 785921 42206 786403
rect 42754 785801 42782 790505
rect 42850 786467 42878 791837
rect 42932 791754 42988 791763
rect 42932 791689 42988 791698
rect 42946 787059 42974 791689
rect 42934 787053 42986 787059
rect 42934 786995 42986 787001
rect 42838 786461 42890 786467
rect 42838 786403 42890 786409
rect 42070 785795 42122 785801
rect 42070 785737 42122 785743
rect 42742 785795 42794 785801
rect 42742 785737 42794 785743
rect 42082 785288 42110 785737
rect 42740 780506 42796 780515
rect 42740 780441 42742 780450
rect 42794 780441 42796 780450
rect 42742 780409 42794 780415
rect 42742 779727 42794 779733
rect 42740 779692 42742 779701
rect 42794 779692 42796 779701
rect 42740 779627 42796 779636
rect 42742 778913 42794 778919
rect 42740 778878 42742 778887
rect 42794 778878 42796 778887
rect 42740 778813 42796 778822
rect 43234 777259 43262 821141
rect 43414 800669 43466 800675
rect 43414 800611 43466 800617
rect 43318 800225 43370 800231
rect 43318 800167 43370 800173
rect 43330 796161 43358 800167
rect 43426 797345 43454 800611
rect 43606 800595 43658 800601
rect 43606 800537 43658 800543
rect 43510 800521 43562 800527
rect 43510 800463 43562 800469
rect 43414 797339 43466 797345
rect 43414 797281 43466 797287
rect 43318 796155 43370 796161
rect 43318 796097 43370 796103
rect 43522 794903 43550 800463
rect 43510 794897 43562 794903
rect 43510 794839 43562 794845
rect 43618 789945 43646 800537
rect 43606 789939 43658 789945
rect 43606 789881 43658 789887
rect 43316 777990 43372 777999
rect 43316 777925 43372 777934
rect 43220 777250 43276 777259
rect 43220 777185 43276 777194
rect 42932 774882 42988 774891
rect 42932 774817 42988 774826
rect 38996 773550 39052 773559
rect 38996 773485 39052 773494
rect 38804 772662 38860 772671
rect 38804 772597 38860 772606
rect 37364 769554 37420 769563
rect 37364 769489 37420 769498
rect 37378 758759 37406 769489
rect 38818 760239 38846 772597
rect 39010 760345 39038 773485
rect 41492 771182 41548 771191
rect 41492 771117 41548 771126
rect 41396 769110 41452 769119
rect 41396 769045 41452 769054
rect 38998 760339 39050 760345
rect 38998 760281 39050 760287
rect 38804 760230 38860 760239
rect 38804 760165 38860 760174
rect 37364 758750 37420 758759
rect 37364 758685 37420 758694
rect 41410 757385 41438 769045
rect 41506 757459 41534 771117
rect 41876 770442 41932 770451
rect 41876 770377 41932 770386
rect 41588 767926 41644 767935
rect 41588 767861 41644 767870
rect 41494 757453 41546 757459
rect 41602 757427 41630 767861
rect 41780 766002 41836 766011
rect 41780 765937 41836 765946
rect 41684 765262 41740 765271
rect 41684 765197 41740 765206
rect 41494 757395 41546 757401
rect 41588 757418 41644 757427
rect 41398 757379 41450 757385
rect 41588 757353 41644 757362
rect 41398 757321 41450 757327
rect 41698 757311 41726 765197
rect 41686 757305 41738 757311
rect 41686 757247 41738 757253
rect 41794 757131 41822 765937
rect 41780 757122 41836 757131
rect 41780 757057 41836 757066
rect 41890 757015 41918 770377
rect 42068 767334 42124 767343
rect 42068 767269 42124 767278
rect 41972 766446 42028 766455
rect 41972 766381 42028 766390
rect 41986 758463 42014 766381
rect 41972 758454 42028 758463
rect 41972 758389 42028 758398
rect 42082 757131 42110 767269
rect 42946 766043 42974 774817
rect 43028 772514 43084 772523
rect 43028 772449 43084 772458
rect 42934 766037 42986 766043
rect 42934 765979 42986 765985
rect 42164 763486 42220 763495
rect 42164 763421 42220 763430
rect 42178 762015 42206 763421
rect 42164 762006 42220 762015
rect 42164 761941 42166 761950
rect 42218 761941 42220 761950
rect 42166 761909 42218 761915
rect 43042 760535 43070 772449
rect 43028 760526 43084 760535
rect 43028 760461 43084 760470
rect 43030 760339 43082 760345
rect 43030 760281 43082 760287
rect 42068 757122 42124 757131
rect 42068 757057 42124 757066
rect 41878 757009 41930 757015
rect 41878 756951 41930 756957
rect 41878 756787 41930 756793
rect 41878 756729 41930 756735
rect 41890 756245 41918 756729
rect 43042 754943 43070 760281
rect 43222 757527 43274 757533
rect 43222 757469 43274 757475
rect 42070 754937 42122 754943
rect 42070 754879 42122 754885
rect 43030 754937 43082 754943
rect 43030 754879 43082 754885
rect 42082 754430 42110 754879
rect 43234 754129 43262 757469
rect 42166 754123 42218 754129
rect 42166 754065 42218 754071
rect 43222 754123 43274 754129
rect 43222 754065 43274 754071
rect 42178 753764 42206 754065
rect 42068 753126 42124 753135
rect 42068 753061 42124 753070
rect 42082 752580 42110 753061
rect 43126 751829 43178 751835
rect 42068 751794 42124 751803
rect 43126 751771 43178 751777
rect 43220 751794 43276 751803
rect 42068 751729 42124 751738
rect 43030 751755 43082 751761
rect 42082 751396 42110 751729
rect 43030 751697 43082 751703
rect 42934 751681 42986 751687
rect 42934 751623 42986 751629
rect 42068 751054 42124 751063
rect 42068 750989 42124 750998
rect 42082 750730 42110 750989
rect 42166 750423 42218 750429
rect 42166 750365 42218 750371
rect 42178 750064 42206 750365
rect 42070 749831 42122 749837
rect 42070 749773 42122 749779
rect 42082 749546 42110 749773
rect 42454 749313 42506 749319
rect 42454 749255 42506 749261
rect 41780 748686 41836 748695
rect 41780 748621 41836 748630
rect 41794 748214 41822 748621
rect 41780 747502 41836 747511
rect 41780 747437 41836 747446
rect 41794 747030 41822 747437
rect 41890 747363 41918 747622
rect 41876 747354 41932 747363
rect 41876 747289 41932 747298
rect 42166 746945 42218 746951
rect 42166 746887 42218 746893
rect 42178 746401 42206 746887
rect 42466 746137 42494 749255
rect 42946 746951 42974 751623
rect 43042 749837 43070 751697
rect 43138 750429 43166 751771
rect 43220 751729 43276 751738
rect 43234 751687 43262 751729
rect 43222 751681 43274 751687
rect 43222 751623 43274 751629
rect 43126 750423 43178 750429
rect 43126 750365 43178 750371
rect 43126 750275 43178 750281
rect 43126 750217 43178 750223
rect 43030 749831 43082 749837
rect 43030 749773 43082 749779
rect 43028 747206 43084 747215
rect 43028 747141 43084 747150
rect 42934 746945 42986 746951
rect 42934 746887 42986 746893
rect 42932 746762 42988 746771
rect 42932 746697 42988 746706
rect 42070 746131 42122 746137
rect 42070 746073 42122 746079
rect 42454 746131 42506 746137
rect 42454 746073 42506 746079
rect 42082 745772 42110 746073
rect 42452 746022 42508 746031
rect 42508 745980 42590 746008
rect 42452 745957 42508 745966
rect 42562 745564 42590 745980
rect 42466 745545 42590 745564
rect 42166 745539 42218 745545
rect 42166 745481 42218 745487
rect 42454 745539 42590 745545
rect 42506 745536 42590 745539
rect 42454 745481 42506 745487
rect 42178 745180 42206 745481
rect 42166 743837 42218 743843
rect 42166 743779 42218 743785
rect 42178 743365 42206 743779
rect 42070 743097 42122 743103
rect 42070 743039 42122 743045
rect 42082 742738 42110 743039
rect 42946 742659 42974 746697
rect 43042 743103 43070 747141
rect 43138 743843 43166 750217
rect 43126 743837 43178 743843
rect 43126 743779 43178 743785
rect 43030 743097 43082 743103
rect 43030 743039 43082 743045
rect 42166 742653 42218 742659
rect 42166 742595 42218 742601
rect 42934 742653 42986 742659
rect 42934 742595 42986 742601
rect 42178 742072 42206 742595
rect 42836 737290 42892 737299
rect 42836 737225 42838 737234
rect 42890 737225 42892 737234
rect 42838 737193 42890 737199
rect 42166 736733 42218 736739
rect 42164 736698 42166 736707
rect 42218 736698 42220 736707
rect 42164 736633 42220 736642
rect 42838 735697 42890 735703
rect 42836 735662 42838 735671
rect 42890 735662 42892 735671
rect 42836 735597 42892 735606
rect 43220 734922 43276 734931
rect 43220 734857 43276 734866
rect 43124 731666 43180 731675
rect 43124 731601 43180 731610
rect 40244 730334 40300 730343
rect 40244 730269 40300 730278
rect 40258 717129 40286 730269
rect 41684 728854 41740 728863
rect 41684 728789 41740 728798
rect 41588 725894 41644 725903
rect 41588 725829 41644 725838
rect 41492 723230 41548 723239
rect 41492 723165 41548 723174
rect 41396 722786 41452 722795
rect 41396 722721 41452 722730
rect 40246 717123 40298 717129
rect 40246 717065 40298 717071
rect 41410 714211 41438 722721
rect 41506 714359 41534 723165
rect 41492 714350 41548 714359
rect 41492 714285 41548 714294
rect 41396 714202 41452 714211
rect 41396 714137 41452 714146
rect 41602 714095 41630 725829
rect 41698 714211 41726 728789
rect 41780 727966 41836 727975
rect 41780 727901 41836 727910
rect 41684 714202 41740 714211
rect 41684 714137 41740 714146
rect 41590 714089 41642 714095
rect 41590 714031 41642 714037
rect 41794 713915 41822 727901
rect 41876 727226 41932 727235
rect 41876 727161 41932 727170
rect 41780 713906 41836 713915
rect 41890 713873 41918 727161
rect 42164 724710 42220 724719
rect 42164 724645 42220 724654
rect 41972 724118 42028 724127
rect 41972 724053 42028 724062
rect 41986 713947 42014 724053
rect 42068 722046 42124 722055
rect 42068 721981 42124 721990
rect 41974 713941 42026 713947
rect 41974 713883 42026 713889
rect 42082 713873 42110 721981
rect 42178 713915 42206 724645
rect 42452 720418 42508 720427
rect 42452 720353 42508 720362
rect 42466 718799 42494 720353
rect 42452 718790 42508 718799
rect 42452 718725 42454 718734
rect 42506 718725 42508 718734
rect 42454 718693 42506 718699
rect 42454 717123 42506 717129
rect 42454 717065 42506 717071
rect 42164 713906 42220 713915
rect 41780 713841 41836 713850
rect 41878 713867 41930 713873
rect 41878 713809 41930 713815
rect 42070 713867 42122 713873
rect 42164 713841 42220 713850
rect 42070 713809 42122 713815
rect 41878 713571 41930 713577
rect 41878 713513 41930 713519
rect 41890 713064 41918 713513
rect 42466 713281 42494 717065
rect 42454 713275 42506 713281
rect 42454 713217 42506 713223
rect 41878 711721 41930 711727
rect 41878 711663 41930 711669
rect 41890 711214 41918 711663
rect 43138 711505 43166 731601
rect 43126 711499 43178 711505
rect 43126 711441 43178 711447
rect 43124 711390 43180 711399
rect 43124 711325 43180 711334
rect 43028 711094 43084 711103
rect 43028 711029 43084 711038
rect 42166 710907 42218 710913
rect 42166 710849 42218 710855
rect 42178 710548 42206 710849
rect 42166 709945 42218 709951
rect 42166 709887 42218 709893
rect 42178 709364 42206 709887
rect 42068 708578 42124 708587
rect 42068 708513 42124 708522
rect 42082 708180 42110 708513
rect 41876 707986 41932 707995
rect 41876 707921 41932 707930
rect 42740 707986 42796 707995
rect 42740 707921 42796 707930
rect 41890 707514 41918 707921
rect 42166 707429 42218 707435
rect 42166 707371 42218 707377
rect 42178 706881 42206 707371
rect 41780 706802 41836 706811
rect 41780 706737 41836 706746
rect 41794 706330 41822 706737
rect 42452 705470 42508 705479
rect 42452 705405 42508 705414
rect 42082 704739 42110 705041
rect 42068 704730 42124 704739
rect 42068 704665 42124 704674
rect 41794 704147 41822 704406
rect 42166 704321 42218 704327
rect 42166 704263 42218 704269
rect 41780 704138 41836 704147
rect 41780 704073 41836 704082
rect 42178 703845 42206 704263
rect 42070 703581 42122 703587
rect 42070 703523 42122 703529
rect 42082 703222 42110 703523
rect 42166 702915 42218 702921
rect 42166 702857 42218 702863
rect 42178 702556 42206 702857
rect 42166 702471 42218 702477
rect 42166 702413 42218 702419
rect 42178 702005 42206 702413
rect 42070 700473 42122 700479
rect 42070 700415 42122 700421
rect 42082 700188 42110 700415
rect 42466 700109 42494 705405
rect 42754 702477 42782 707921
rect 43042 704327 43070 711029
rect 43138 709951 43166 711325
rect 43126 709945 43178 709951
rect 43126 709887 43178 709893
rect 43124 709762 43180 709771
rect 43124 709697 43180 709706
rect 43030 704321 43082 704327
rect 43030 704263 43082 704269
rect 43030 704173 43082 704179
rect 43030 704115 43082 704121
rect 43042 702921 43070 704115
rect 43138 703587 43166 709697
rect 43126 703581 43178 703587
rect 43126 703523 43178 703529
rect 43126 703433 43178 703439
rect 43126 703375 43178 703381
rect 43030 702915 43082 702921
rect 43030 702857 43082 702863
rect 43028 702806 43084 702815
rect 43028 702741 43084 702750
rect 42742 702471 42794 702477
rect 42742 702413 42794 702419
rect 42166 700103 42218 700109
rect 42166 700045 42218 700051
rect 42454 700103 42506 700109
rect 42454 700045 42506 700051
rect 42178 699522 42206 700045
rect 42454 699881 42506 699887
rect 42454 699823 42506 699829
rect 42166 699215 42218 699221
rect 42166 699157 42218 699163
rect 42178 698856 42206 699157
rect 42466 693491 42494 699823
rect 43042 699221 43070 702741
rect 43138 700479 43166 703375
rect 43126 700473 43178 700479
rect 43126 700415 43178 700421
rect 43030 699215 43082 699221
rect 43030 699157 43082 699163
rect 42836 694074 42892 694083
rect 42836 694009 42838 694018
rect 42890 694009 42892 694018
rect 42838 693977 42890 693983
rect 42452 693482 42508 693491
rect 42452 693417 42508 693426
rect 42454 692777 42506 692783
rect 42452 692742 42454 692751
rect 42506 692742 42508 692751
rect 42452 692677 42508 692686
rect 43234 690827 43262 734857
rect 43330 734043 43358 777925
rect 43798 766037 43850 766043
rect 43798 765979 43850 765985
rect 43702 757453 43754 757459
rect 43702 757395 43754 757401
rect 43606 757379 43658 757385
rect 43606 757321 43658 757327
rect 43510 757305 43562 757311
rect 43510 757247 43562 757253
rect 43522 752076 43550 757247
rect 43426 752048 43550 752076
rect 43426 751835 43454 752048
rect 43414 751829 43466 751835
rect 43414 751771 43466 751777
rect 43618 749319 43646 757321
rect 43714 751909 43742 757395
rect 43702 751903 43754 751909
rect 43702 751845 43754 751851
rect 43810 750281 43838 765979
rect 43798 750275 43850 750281
rect 43798 750217 43850 750223
rect 43606 749313 43658 749319
rect 43606 749255 43658 749261
rect 43316 734034 43372 734043
rect 43316 733969 43372 733978
rect 43510 714311 43562 714317
rect 43510 714253 43562 714259
rect 43414 713941 43466 713947
rect 43414 713883 43466 713889
rect 43318 713867 43370 713873
rect 43318 713809 43370 713815
rect 43330 707435 43358 713809
rect 43426 711547 43454 713883
rect 43412 711538 43468 711547
rect 43412 711473 43468 711482
rect 43414 711425 43466 711431
rect 43414 711367 43466 711373
rect 43318 707429 43370 707435
rect 43318 707371 43370 707377
rect 43426 704179 43454 711367
rect 43522 710913 43550 714253
rect 43702 714089 43754 714095
rect 43702 714031 43754 714037
rect 43606 711499 43658 711505
rect 43606 711441 43658 711447
rect 43510 710907 43562 710913
rect 43510 710849 43562 710855
rect 43414 704173 43466 704179
rect 43414 704115 43466 704121
rect 43618 703439 43646 711441
rect 43714 711431 43742 714031
rect 43702 711425 43754 711431
rect 43702 711367 43754 711373
rect 43606 703433 43658 703439
rect 43606 703375 43658 703381
rect 43508 691706 43564 691715
rect 43508 691641 43564 691650
rect 43220 690818 43276 690827
rect 43220 690753 43276 690762
rect 41684 688302 41740 688311
rect 41684 688237 41740 688246
rect 40148 687118 40204 687127
rect 40148 687053 40204 687062
rect 37364 683270 37420 683279
rect 37364 683205 37420 683214
rect 37378 672623 37406 683205
rect 37364 672614 37420 672623
rect 37364 672549 37420 672558
rect 40162 672285 40190 687053
rect 40244 686378 40300 686387
rect 40244 686313 40300 686322
rect 40258 673955 40286 686313
rect 40916 684898 40972 684907
rect 40916 684833 40972 684842
rect 40244 673946 40300 673955
rect 40244 673881 40300 673890
rect 40150 672279 40202 672285
rect 40150 672221 40202 672227
rect 40930 670953 40958 684833
rect 41300 681494 41356 681503
rect 41300 681429 41356 681438
rect 41314 670995 41342 681429
rect 41300 670986 41356 670995
rect 40918 670947 40970 670953
rect 41300 670921 41356 670930
rect 40918 670889 40970 670895
rect 41698 670879 41726 688237
rect 41780 685638 41836 685647
rect 41780 685573 41836 685582
rect 41794 674579 41822 685573
rect 41972 684010 42028 684019
rect 41972 683945 42028 683954
rect 41876 679570 41932 679579
rect 41876 679505 41932 679514
rect 41782 674573 41834 674579
rect 41782 674515 41834 674521
rect 41782 672279 41834 672285
rect 41782 672221 41834 672227
rect 41686 670873 41738 670879
rect 41686 670815 41738 670821
rect 41794 670657 41822 672221
rect 41890 670731 41918 679505
rect 41986 674672 42014 683945
rect 42068 682678 42124 682687
rect 42068 682613 42124 682622
rect 42082 674820 42110 682613
rect 43028 681346 43084 681355
rect 43028 681281 43084 681290
rect 42164 678830 42220 678839
rect 42164 678765 42220 678774
rect 42178 675023 42206 678765
rect 42452 676758 42508 676767
rect 42452 676693 42508 676702
rect 42466 675837 42494 676693
rect 42454 675831 42506 675837
rect 42454 675773 42506 675779
rect 42466 675731 42494 675773
rect 42452 675722 42508 675731
rect 42452 675657 42508 675666
rect 42166 675017 42218 675023
rect 42166 674959 42218 674965
rect 42454 675017 42506 675023
rect 42454 674959 42506 674965
rect 42082 674792 42206 674820
rect 41986 674644 42110 674672
rect 41974 674573 42026 674579
rect 41974 674515 42026 674521
rect 41986 670847 42014 674515
rect 41972 670838 42028 670847
rect 41972 670773 42028 670782
rect 41878 670725 41930 670731
rect 42082 670699 42110 674644
rect 42178 670995 42206 674792
rect 42164 670986 42220 670995
rect 42164 670921 42220 670930
rect 42166 670873 42218 670879
rect 42164 670838 42166 670847
rect 42218 670838 42220 670847
rect 42164 670773 42220 670782
rect 41878 670667 41930 670673
rect 42068 670690 42124 670699
rect 41782 670651 41834 670657
rect 42068 670625 42124 670634
rect 41782 670593 41834 670599
rect 42164 670394 42220 670403
rect 42164 670329 42220 670338
rect 42178 669848 42206 670329
rect 42466 670139 42494 674959
rect 43042 670824 43070 681281
rect 43124 678238 43180 678247
rect 43124 678173 43180 678182
rect 43138 670995 43166 678173
rect 43124 670986 43180 670995
rect 43124 670921 43180 670930
rect 43318 670947 43370 670953
rect 43318 670889 43370 670895
rect 43042 670796 43262 670824
rect 43030 670725 43082 670731
rect 43030 670667 43082 670673
rect 42454 670133 42506 670139
rect 42454 670075 42506 670081
rect 43042 668955 43070 670667
rect 43126 670651 43178 670657
rect 43126 670593 43178 670599
rect 43030 668949 43082 668955
rect 43030 668891 43082 668897
rect 42742 668727 42794 668733
rect 42742 668669 42794 668675
rect 42838 668727 42890 668733
rect 42838 668669 42890 668675
rect 42166 668579 42218 668585
rect 42166 668521 42218 668527
rect 42178 667998 42206 668521
rect 42166 667913 42218 667919
rect 42166 667855 42218 667861
rect 42178 667361 42206 667855
rect 42166 666729 42218 666735
rect 42166 666671 42218 666677
rect 42178 666148 42206 666671
rect 42164 665362 42220 665371
rect 42164 665297 42220 665306
rect 42178 664964 42206 665297
rect 42166 664879 42218 664885
rect 42166 664821 42218 664827
rect 42178 664298 42206 664821
rect 42070 664213 42122 664219
rect 42070 664155 42122 664161
rect 42082 663706 42110 664155
rect 42166 663547 42218 663553
rect 42166 663489 42218 663495
rect 42178 663114 42206 663489
rect 42452 662846 42508 662855
rect 42452 662781 42508 662790
rect 42178 661523 42206 661856
rect 42164 661514 42220 661523
rect 42164 661449 42220 661458
rect 42082 661056 42110 661190
rect 42082 661028 42206 661056
rect 42070 660883 42122 660889
rect 42070 660825 42122 660831
rect 42082 660672 42110 660825
rect 42178 660783 42206 661028
rect 42164 660774 42220 660783
rect 42164 660709 42220 660718
rect 41780 660330 41836 660339
rect 41780 660265 41836 660274
rect 41794 660006 41822 660265
rect 42166 659699 42218 659705
rect 42166 659641 42218 659647
rect 42178 659340 42206 659641
rect 41876 659146 41932 659155
rect 41876 659081 41932 659090
rect 41890 658822 41918 659081
rect 42466 657411 42494 662781
rect 42754 660889 42782 668669
rect 42850 663553 42878 668669
rect 43138 668585 43166 670593
rect 43126 668579 43178 668585
rect 43126 668521 43178 668527
rect 43234 668456 43262 670796
rect 43330 668733 43358 670889
rect 43414 670133 43466 670139
rect 43414 670075 43466 670081
rect 43318 668727 43370 668733
rect 43318 668669 43370 668675
rect 43138 668428 43262 668456
rect 43138 666735 43166 668428
rect 43126 666729 43178 666735
rect 43426 666680 43454 670075
rect 43126 666671 43178 666677
rect 43234 666652 43454 666680
rect 43234 666532 43262 666652
rect 43138 666504 43262 666532
rect 43138 664219 43166 666504
rect 43126 664213 43178 664219
rect 43126 664155 43178 664161
rect 42838 663547 42890 663553
rect 42838 663489 42890 663495
rect 42836 663438 42892 663447
rect 42836 663373 42892 663382
rect 42742 660883 42794 660889
rect 42742 660825 42794 660831
rect 42850 659705 42878 663373
rect 43124 662402 43180 662411
rect 43124 662337 43180 662346
rect 42838 659699 42890 659705
rect 42838 659641 42890 659647
rect 42070 657405 42122 657411
rect 42070 657347 42122 657353
rect 42454 657405 42506 657411
rect 42454 657347 42506 657353
rect 42082 656972 42110 657347
rect 42454 656739 42506 656745
rect 42454 656681 42506 656687
rect 41780 656630 41836 656639
rect 41780 656565 41836 656574
rect 41794 656306 41822 656565
rect 42166 656221 42218 656227
rect 42166 656163 42218 656169
rect 42178 655677 42206 656163
rect 42466 651163 42494 656681
rect 43138 656227 43166 662337
rect 43126 656221 43178 656227
rect 43126 656163 43178 656169
rect 42452 651154 42508 651163
rect 42452 651089 42508 651098
rect 42452 649822 42508 649831
rect 42452 649757 42454 649766
rect 42506 649757 42508 649766
rect 42454 649725 42506 649731
rect 42454 649561 42506 649567
rect 42452 649526 42454 649535
rect 42506 649526 42508 649535
rect 42452 649461 42508 649470
rect 43220 648490 43276 648499
rect 43220 648425 43276 648434
rect 43124 645382 43180 645391
rect 43124 645317 43180 645326
rect 39860 643902 39916 643911
rect 39860 643837 39916 643846
rect 37364 640054 37420 640063
rect 37364 639989 37420 639998
rect 37378 628223 37406 639989
rect 37364 628214 37420 628223
rect 37364 628149 37420 628158
rect 39874 627885 39902 643837
rect 39956 643162 40012 643171
rect 39956 643097 40012 643106
rect 39970 627927 39998 643097
rect 41492 642422 41548 642431
rect 41492 642357 41548 642366
rect 41300 639462 41356 639471
rect 41300 639397 41356 639406
rect 39956 627918 40012 627927
rect 39862 627879 39914 627885
rect 39956 627853 40012 627862
rect 39862 627821 39914 627827
rect 41314 627779 41342 639397
rect 41506 627811 41534 642357
rect 41684 641682 41740 641691
rect 41684 641617 41740 641626
rect 41588 636354 41644 636363
rect 41588 636289 41644 636298
rect 41494 627805 41546 627811
rect 41300 627770 41356 627779
rect 41602 627779 41630 636289
rect 41494 627747 41546 627753
rect 41588 627770 41644 627779
rect 41300 627705 41356 627714
rect 41698 627737 41726 641617
rect 41876 640794 41932 640803
rect 41876 640729 41932 640738
rect 41588 627705 41644 627714
rect 41686 627731 41738 627737
rect 41686 627673 41738 627679
rect 41890 627441 41918 640729
rect 41972 637686 42028 637695
rect 41972 637621 42028 637630
rect 41986 627441 42014 637621
rect 42068 636798 42124 636807
rect 42068 636733 42124 636742
rect 42082 627483 42110 636733
rect 42164 635614 42220 635623
rect 42164 635549 42220 635558
rect 42178 627631 42206 635549
rect 43028 635022 43084 635031
rect 43028 634957 43084 634966
rect 42452 633542 42508 633551
rect 42452 633477 42508 633486
rect 42466 632367 42494 633477
rect 42452 632358 42508 632367
rect 42452 632293 42508 632302
rect 42466 630771 42494 632293
rect 42454 630765 42506 630771
rect 42454 630707 42506 630713
rect 43042 628052 43070 634957
rect 43138 630845 43166 645317
rect 43126 630839 43178 630845
rect 43126 630781 43178 630787
rect 43042 628024 43166 628052
rect 43138 627885 43166 628024
rect 43030 627879 43082 627885
rect 43030 627821 43082 627827
rect 43126 627879 43178 627885
rect 43126 627821 43178 627827
rect 42164 627622 42220 627631
rect 42164 627557 42220 627566
rect 42068 627474 42124 627483
rect 41878 627435 41930 627441
rect 41878 627377 41930 627383
rect 41974 627435 42026 627441
rect 42068 627409 42124 627418
rect 42934 627435 42986 627441
rect 41974 627377 42026 627383
rect 42934 627377 42986 627383
rect 41878 627213 41930 627219
rect 41878 627155 41930 627161
rect 41890 626632 41918 627155
rect 42166 625363 42218 625369
rect 42166 625305 42218 625311
rect 42178 624782 42206 625305
rect 42166 624697 42218 624703
rect 42166 624639 42218 624645
rect 42178 624161 42206 624639
rect 42946 623519 42974 627377
rect 43042 625369 43070 627821
rect 43126 627731 43178 627737
rect 43126 627673 43178 627679
rect 43030 625363 43082 625369
rect 43030 625305 43082 625311
rect 43030 625215 43082 625221
rect 43030 625157 43082 625163
rect 42166 623513 42218 623519
rect 42166 623455 42218 623461
rect 42934 623513 42986 623519
rect 42934 623455 42986 623461
rect 42178 622965 42206 623455
rect 42934 623365 42986 623371
rect 42934 623307 42986 623313
rect 42166 622255 42218 622261
rect 42166 622197 42218 622203
rect 42178 621748 42206 622197
rect 42068 621702 42124 621711
rect 42068 621637 42124 621646
rect 42082 621125 42110 621637
rect 41972 620814 42028 620823
rect 41972 620749 42028 620758
rect 41986 620490 42014 620749
rect 42166 620405 42218 620411
rect 42166 620347 42218 620353
rect 42178 619929 42206 620347
rect 42946 620060 42974 623307
rect 43042 622261 43070 625157
rect 43030 622255 43082 622261
rect 43030 622197 43082 622203
rect 43138 620411 43166 627673
rect 43126 620405 43178 620411
rect 43126 620347 43178 620353
rect 42946 620032 43166 620060
rect 41780 618298 41836 618307
rect 41780 618233 41836 618242
rect 41794 617974 41822 618233
rect 41986 618159 42014 618640
rect 41972 618150 42028 618159
rect 41972 618085 42028 618094
rect 41780 617854 41836 617863
rect 41780 617789 41836 617798
rect 41794 617456 41822 617789
rect 42166 617371 42218 617377
rect 42166 617313 42218 617319
rect 42178 616790 42206 617313
rect 41780 616522 41836 616531
rect 41780 616457 41836 616466
rect 41794 616157 41822 616457
rect 43138 615897 43166 620032
rect 42166 615891 42218 615897
rect 42166 615833 42218 615839
rect 43126 615891 43178 615897
rect 43126 615833 43178 615839
rect 42178 615606 42206 615833
rect 42166 614189 42218 614195
rect 42166 614131 42218 614137
rect 42178 613756 42206 614131
rect 42742 613523 42794 613529
rect 42742 613465 42794 613471
rect 41780 613414 41836 613423
rect 41780 613349 41836 613358
rect 41794 613121 41822 613349
rect 41780 612822 41836 612831
rect 41780 612757 41836 612766
rect 41794 612498 41822 612757
rect 42754 607905 42782 613465
rect 42166 607899 42218 607905
rect 42166 607841 42218 607847
rect 42742 607899 42794 607905
rect 42742 607841 42794 607847
rect 42178 606319 42206 607841
rect 42742 607751 42794 607757
rect 42740 607716 42742 607725
rect 42794 607716 42796 607725
rect 42740 607651 42796 607660
rect 42740 606902 42796 606911
rect 42740 606837 42742 606846
rect 42794 606837 42796 606846
rect 42742 606805 42794 606811
rect 42164 606310 42220 606319
rect 42164 606245 42220 606254
rect 43234 604691 43262 648425
rect 43522 647611 43550 691641
rect 43892 680606 43948 680615
rect 43892 680541 43948 680550
rect 43606 673759 43658 673765
rect 43606 673701 43658 673707
rect 43618 669344 43646 673701
rect 43618 669316 43742 669344
rect 43714 667919 43742 669316
rect 43702 667913 43754 667919
rect 43702 667855 43754 667861
rect 43906 665329 43934 680541
rect 43606 665323 43658 665329
rect 43606 665265 43658 665271
rect 43894 665323 43946 665329
rect 43894 665265 43946 665271
rect 43618 664885 43646 665265
rect 43606 664879 43658 664885
rect 43606 664821 43658 664827
rect 43508 647602 43564 647611
rect 43508 647537 43564 647546
rect 43604 647010 43660 647019
rect 43604 646945 43660 646954
rect 43414 627953 43466 627959
rect 43414 627895 43466 627901
rect 43318 627879 43370 627885
rect 43318 627821 43370 627827
rect 43330 625221 43358 627821
rect 43318 625215 43370 625221
rect 43318 625157 43370 625163
rect 43316 625106 43372 625115
rect 43316 625041 43372 625050
rect 43330 617377 43358 625041
rect 43426 624703 43454 627895
rect 43510 627805 43562 627811
rect 43510 627747 43562 627753
rect 43414 624697 43466 624703
rect 43414 624639 43466 624645
rect 43522 623371 43550 627747
rect 43510 623365 43562 623371
rect 43510 623307 43562 623313
rect 43318 617371 43370 617377
rect 43318 617313 43370 617319
rect 43508 605274 43564 605283
rect 43508 605209 43564 605218
rect 43220 604682 43276 604691
rect 43220 604617 43276 604626
rect 43412 602906 43468 602915
rect 43412 602841 43468 602850
rect 41588 601870 41644 601879
rect 41588 601805 41644 601814
rect 40052 600686 40108 600695
rect 40052 600621 40108 600630
rect 40066 586001 40094 600621
rect 41396 598466 41452 598475
rect 41396 598401 41452 598410
rect 40054 585995 40106 586001
rect 40054 585937 40106 585943
rect 41410 584563 41438 598401
rect 41492 596246 41548 596255
rect 41492 596181 41548 596190
rect 41506 584711 41534 596181
rect 41602 584859 41630 601805
rect 41876 599206 41932 599215
rect 41876 599141 41932 599150
rect 41780 595210 41836 595219
rect 41780 595145 41836 595154
rect 41588 584850 41644 584859
rect 41588 584785 41644 584794
rect 41492 584702 41548 584711
rect 41492 584637 41548 584646
rect 41396 584554 41452 584563
rect 41396 584489 41452 584498
rect 41794 584299 41822 595145
rect 41890 586149 41918 599141
rect 41972 597578 42028 597587
rect 41972 597513 42028 597522
rect 41878 586143 41930 586149
rect 41878 586085 41930 586091
rect 41878 585995 41930 586001
rect 41878 585937 41930 585943
rect 41890 584415 41918 585937
rect 41876 584406 41932 584415
rect 41876 584341 41932 584350
rect 41782 584293 41834 584299
rect 41782 584235 41834 584241
rect 41986 584225 42014 597513
rect 42068 593138 42124 593147
rect 42068 593073 42124 593082
rect 42082 584267 42110 593073
rect 42164 592398 42220 592407
rect 42164 592333 42220 592342
rect 42068 584258 42124 584267
rect 41974 584219 42026 584225
rect 42178 584225 42206 592333
rect 42836 591806 42892 591815
rect 42836 591741 42892 591750
rect 42740 590474 42796 590483
rect 42740 590409 42796 590418
rect 42754 589447 42782 590409
rect 42740 589438 42796 589447
rect 42740 589373 42796 589382
rect 42742 586143 42794 586149
rect 42742 586085 42794 586091
rect 42754 584711 42782 586085
rect 42740 584702 42796 584711
rect 42740 584637 42796 584646
rect 42068 584193 42124 584202
rect 42166 584219 42218 584225
rect 41974 584161 42026 584167
rect 42166 584161 42218 584167
rect 41974 583997 42026 584003
rect 41974 583939 42026 583945
rect 41986 583445 42014 583939
rect 42850 583823 42878 591741
rect 43126 584737 43178 584743
rect 43126 584679 43178 584685
rect 42836 583814 42892 583823
rect 42836 583749 42892 583758
rect 41972 582038 42028 582047
rect 41972 581973 42028 581982
rect 41986 581605 42014 581973
rect 43030 581555 43082 581561
rect 43030 581497 43082 581503
rect 42070 581481 42122 581487
rect 42070 581423 42122 581429
rect 42932 581446 42988 581455
rect 42082 580974 42110 581423
rect 42932 581381 42988 581390
rect 41780 580262 41836 580271
rect 41780 580197 41836 580206
rect 41794 579790 41822 580197
rect 42164 578930 42220 578939
rect 42164 578865 42220 578874
rect 42178 578569 42206 578865
rect 42946 578453 42974 581381
rect 42934 578447 42986 578453
rect 42934 578389 42986 578395
rect 42932 578338 42988 578347
rect 42070 578299 42122 578305
rect 42932 578273 42988 578282
rect 42070 578241 42122 578247
rect 42082 577940 42110 578241
rect 42166 577707 42218 577713
rect 42166 577649 42218 577655
rect 42178 577274 42206 577649
rect 41780 577006 41836 577015
rect 41780 576941 41836 576950
rect 41794 576756 41822 576941
rect 42452 576414 42508 576423
rect 42452 576349 42508 576358
rect 41780 575970 41836 575979
rect 41780 575905 41836 575914
rect 41794 575424 41822 575905
rect 41780 575082 41836 575091
rect 41780 575017 41836 575026
rect 41794 574797 41822 575017
rect 42164 574638 42220 574647
rect 42164 574573 42220 574582
rect 42178 574240 42206 574573
rect 42166 574155 42218 574161
rect 42166 574097 42218 574103
rect 42178 573574 42206 574097
rect 42466 573273 42494 576349
rect 42070 573267 42122 573273
rect 42070 573209 42122 573215
rect 42454 573267 42506 573273
rect 42454 573209 42506 573215
rect 42082 572982 42110 573209
rect 42452 573158 42508 573167
rect 42452 573093 42508 573102
rect 42166 572823 42218 572829
rect 42166 572765 42218 572771
rect 42178 572390 42206 572765
rect 42466 572681 42494 573093
rect 42946 572829 42974 578273
rect 43042 577713 43070 581497
rect 43138 581487 43166 584679
rect 43222 584293 43274 584299
rect 43222 584235 43274 584241
rect 43126 581481 43178 581487
rect 43126 581423 43178 581429
rect 43234 581284 43262 584235
rect 43318 584219 43370 584225
rect 43318 584161 43370 584167
rect 43330 581561 43358 584161
rect 43318 581555 43370 581561
rect 43318 581497 43370 581503
rect 43138 581256 43262 581284
rect 43030 577707 43082 577713
rect 43030 577649 43082 577655
rect 43028 577598 43084 577607
rect 43028 577533 43084 577542
rect 42934 572823 42986 572829
rect 42934 572765 42986 572771
rect 42454 572675 42506 572681
rect 42454 572617 42506 572623
rect 42934 572675 42986 572681
rect 42934 572617 42986 572623
rect 42166 571047 42218 571053
rect 42166 570989 42218 570995
rect 42178 570540 42206 570989
rect 42166 570381 42218 570387
rect 42082 570329 42166 570332
rect 42082 570323 42218 570329
rect 42082 570304 42206 570323
rect 42838 570307 42890 570313
rect 42082 569948 42110 570304
rect 42838 570249 42890 570255
rect 42070 569789 42122 569795
rect 42070 569731 42122 569737
rect 42082 569282 42110 569731
rect 34484 564722 34540 564731
rect 34484 564657 34540 564666
rect 34498 564541 34526 564657
rect 34486 564535 34538 564541
rect 34486 564477 34538 564483
rect 42164 563538 42220 563547
rect 42164 563473 42166 563482
rect 42218 563473 42220 563482
rect 42166 563441 42218 563447
rect 42850 562881 42878 570249
rect 42946 569795 42974 572617
rect 43042 571053 43070 577533
rect 43138 574161 43166 581256
rect 43126 574155 43178 574161
rect 43126 574097 43178 574103
rect 43124 574046 43180 574055
rect 43124 573981 43180 573990
rect 43030 571047 43082 571053
rect 43030 570989 43082 570995
rect 43138 570387 43166 573981
rect 43126 570381 43178 570387
rect 43126 570323 43178 570329
rect 42934 569789 42986 569795
rect 42934 569731 42986 569737
rect 42836 562872 42892 562881
rect 42836 562807 42892 562816
rect 43220 562058 43276 562067
rect 43220 561993 43276 562002
rect 42932 558950 42988 558959
rect 42932 558885 42988 558894
rect 40244 557470 40300 557479
rect 40244 557405 40300 557414
rect 40258 544265 40286 557405
rect 41396 555990 41452 555999
rect 41396 555925 41452 555934
rect 41684 555990 41740 555999
rect 41684 555925 41740 555934
rect 41410 553039 41438 555925
rect 41396 553030 41452 553039
rect 41396 552965 41452 552974
rect 41588 551994 41644 552003
rect 41588 551929 41644 551938
rect 41602 544728 41630 551929
rect 41410 544700 41630 544728
rect 40246 544259 40298 544265
rect 40246 544201 40298 544207
rect 41014 544259 41066 544265
rect 41014 544201 41066 544207
rect 41026 544159 41054 544201
rect 41012 544150 41068 544159
rect 41012 544085 41068 544094
rect 41410 541379 41438 544700
rect 41698 544580 41726 555925
rect 42164 555250 42220 555259
rect 42164 555185 42220 555194
rect 41972 554362 42028 554371
rect 41972 554297 42028 554306
rect 41780 553030 41836 553039
rect 41780 552965 41836 552974
rect 41506 544552 41726 544580
rect 41398 541373 41450 541379
rect 41506 541347 41534 544552
rect 41794 544432 41822 552965
rect 41878 544555 41930 544561
rect 41878 544497 41930 544503
rect 41698 544404 41822 544432
rect 41698 541347 41726 544404
rect 41398 541315 41450 541321
rect 41492 541338 41548 541347
rect 41492 541273 41548 541282
rect 41684 541338 41740 541347
rect 41684 541273 41740 541282
rect 41890 541051 41918 544497
rect 41876 541042 41932 541051
rect 41986 541009 42014 554297
rect 42068 550070 42124 550079
rect 42068 550005 42124 550014
rect 42082 541009 42110 550005
rect 42178 544561 42206 555185
rect 42452 551402 42508 551411
rect 42508 551360 42590 551388
rect 42452 551337 42508 551346
rect 42452 551254 42508 551263
rect 42452 551189 42508 551198
rect 42166 544555 42218 544561
rect 42166 544497 42218 544503
rect 42466 544413 42494 551189
rect 42166 544407 42218 544413
rect 42166 544349 42218 544355
rect 42454 544407 42506 544413
rect 42454 544349 42506 544355
rect 42178 541051 42206 544349
rect 42452 541190 42508 541199
rect 42562 541176 42590 551360
rect 42946 549464 42974 558885
rect 42946 549436 43070 549464
rect 43042 549390 43070 549436
rect 43042 549362 43166 549390
rect 42932 549330 42988 549339
rect 42932 549265 42988 549274
rect 42946 541675 42974 549265
rect 43028 548590 43084 548599
rect 43028 548525 43084 548534
rect 42934 541669 42986 541675
rect 42934 541611 42986 541617
rect 42934 541521 42986 541527
rect 42934 541463 42986 541469
rect 42508 541148 42590 541176
rect 42452 541125 42508 541134
rect 42164 541042 42220 541051
rect 41876 540977 41932 540986
rect 41974 541003 42026 541009
rect 41974 540945 42026 540951
rect 42070 541003 42122 541009
rect 42164 540977 42220 540986
rect 42454 541003 42506 541009
rect 42070 540945 42122 540951
rect 42506 540963 42590 540991
rect 42454 540945 42506 540951
rect 41974 540781 42026 540787
rect 41974 540723 42026 540729
rect 41986 540245 42014 540723
rect 41876 538970 41932 538979
rect 41876 538905 41932 538914
rect 41890 538424 41918 538905
rect 42166 538339 42218 538345
rect 42166 538281 42218 538287
rect 42178 537758 42206 538281
rect 42068 537046 42124 537055
rect 42068 536981 42124 536990
rect 42082 536574 42110 536981
rect 42070 535823 42122 535829
rect 42070 535765 42122 535771
rect 42082 535390 42110 535765
rect 42164 535270 42220 535279
rect 42164 535205 42220 535214
rect 42178 534724 42206 535205
rect 42166 534639 42218 534645
rect 42166 534581 42218 534587
rect 42178 534058 42206 534581
rect 41972 533790 42028 533799
rect 41972 533725 42028 533734
rect 41986 533540 42014 533725
rect 42164 532754 42220 532763
rect 42164 532689 42220 532698
rect 42178 532241 42206 532689
rect 41780 531866 41836 531875
rect 41780 531801 41836 531810
rect 41794 531616 41822 531801
rect 42166 531531 42218 531537
rect 42166 531473 42218 531479
rect 42454 531531 42506 531537
rect 42562 531519 42590 540963
rect 42946 538345 42974 541463
rect 42934 538339 42986 538345
rect 42934 538281 42986 538287
rect 42934 538191 42986 538197
rect 42934 538133 42986 538139
rect 42946 534645 42974 538133
rect 43042 535829 43070 548525
rect 43030 535823 43082 535829
rect 43030 535765 43082 535771
rect 43030 535675 43082 535681
rect 43030 535617 43082 535623
rect 42934 534639 42986 534645
rect 42934 534581 42986 534587
rect 42932 534530 42988 534539
rect 42932 534465 42988 534474
rect 42506 531491 42590 531519
rect 42454 531473 42506 531479
rect 42178 531024 42206 531473
rect 42452 531422 42508 531431
rect 42452 531357 42508 531366
rect 42166 530939 42218 530945
rect 42166 530881 42218 530887
rect 42178 530401 42206 530881
rect 42070 530199 42122 530205
rect 42070 530141 42122 530147
rect 42082 529766 42110 530141
rect 42466 529465 42494 531357
rect 42946 530205 42974 534465
rect 43042 530945 43070 535617
rect 43030 530939 43082 530945
rect 43030 530881 43082 530887
rect 42934 530199 42986 530205
rect 42934 530141 42986 530147
rect 42932 530090 42988 530099
rect 42932 530025 42988 530034
rect 42166 529459 42218 529465
rect 42166 529401 42218 529407
rect 42454 529459 42506 529465
rect 42454 529401 42506 529407
rect 42178 529205 42206 529401
rect 42166 527683 42218 527689
rect 42166 527625 42218 527631
rect 42178 527365 42206 527625
rect 42946 527245 42974 530025
rect 43030 529977 43082 529983
rect 43030 529919 43082 529925
rect 42070 527239 42122 527245
rect 42070 527181 42122 527187
rect 42934 527239 42986 527245
rect 42934 527181 42986 527187
rect 42082 526732 42110 527181
rect 41780 526538 41836 526547
rect 41780 526473 41836 526482
rect 41794 526066 41822 526473
rect 41588 524170 41644 524179
rect 41588 524105 41644 524114
rect 41602 504051 41630 524105
rect 43042 519845 43070 529919
rect 43138 527689 43166 549362
rect 43126 527683 43178 527689
rect 43126 527625 43178 527631
rect 41878 519839 41930 519845
rect 41878 519781 41930 519787
rect 43030 519839 43082 519845
rect 43030 519781 43082 519787
rect 41588 504042 41644 504051
rect 41588 503977 41644 503986
rect 41780 491018 41836 491027
rect 41780 490953 41836 490962
rect 41794 481111 41822 490953
rect 41780 481102 41836 481111
rect 41780 481037 41836 481046
rect 41890 435527 41918 519781
rect 42164 510110 42220 510119
rect 42164 510045 42220 510054
rect 42178 504051 42206 510045
rect 42164 504042 42220 504051
rect 42164 503977 42220 503986
rect 42262 437181 42314 437187
rect 42260 437146 42262 437155
rect 42314 437146 42316 437155
rect 42260 437081 42316 437090
rect 42262 436293 42314 436299
rect 42260 436258 42262 436267
rect 42314 436258 42316 436267
rect 42260 436193 42316 436202
rect 41876 435518 41932 435527
rect 41876 435453 41932 435462
rect 43234 433603 43262 561993
rect 43426 559847 43454 602841
rect 43522 561623 43550 605209
rect 43618 603803 43646 646945
rect 43796 646122 43852 646131
rect 43796 646057 43852 646066
rect 43702 630839 43754 630845
rect 43702 630781 43754 630787
rect 43714 614195 43742 630781
rect 43702 614189 43754 614195
rect 43702 614131 43754 614137
rect 43604 603794 43660 603803
rect 43604 603729 43660 603738
rect 43508 561614 43564 561623
rect 43508 561549 43564 561558
rect 43618 560587 43646 603729
rect 43810 602915 43838 646057
rect 43796 602906 43852 602915
rect 43796 602841 43852 602850
rect 43604 560578 43660 560587
rect 43604 560513 43660 560522
rect 43412 559838 43468 559847
rect 43412 559773 43468 559782
rect 43316 547702 43372 547711
rect 43316 547637 43372 547646
rect 43330 546231 43358 547637
rect 43316 546222 43372 546231
rect 43316 546157 43372 546166
rect 43330 544857 43358 546157
rect 43318 544851 43370 544857
rect 43318 544793 43370 544799
rect 43318 541669 43370 541675
rect 43318 541611 43370 541617
rect 43330 538197 43358 541611
rect 43318 538191 43370 538197
rect 43318 538133 43370 538139
rect 43316 434482 43372 434491
rect 43316 434417 43372 434426
rect 43220 433594 43276 433603
rect 43220 433529 43276 433538
rect 41972 429894 42028 429903
rect 41972 429829 42028 429838
rect 41780 426934 41836 426943
rect 41780 426869 41836 426878
rect 37364 423678 37420 423687
rect 37364 423613 37420 423622
rect 37268 422050 37324 422059
rect 37268 421985 37324 421994
rect 37282 414765 37310 421985
rect 37378 416541 37406 423613
rect 40148 423234 40204 423243
rect 40148 423169 40204 423178
rect 37366 416535 37418 416541
rect 37366 416477 37418 416483
rect 40162 415209 40190 423169
rect 40244 421310 40300 421319
rect 40244 421245 40300 421254
rect 40258 415431 40286 421245
rect 40246 415425 40298 415431
rect 40246 415367 40298 415373
rect 40150 415203 40202 415209
rect 40150 415145 40202 415151
rect 37270 414759 37322 414765
rect 37270 414701 37322 414707
rect 41794 413433 41822 426869
rect 41986 418336 42014 429829
rect 43330 429140 43358 434417
rect 43426 432123 43454 559773
rect 43510 541373 43562 541379
rect 43510 541315 43562 541321
rect 43522 535681 43550 541315
rect 43510 535675 43562 535681
rect 43510 535617 43562 535623
rect 43618 433011 43646 560513
rect 44566 544851 44618 544857
rect 44566 544793 44618 544799
rect 43604 433002 43660 433011
rect 43604 432937 43660 432946
rect 43412 432114 43468 432123
rect 43412 432049 43468 432058
rect 43234 429112 43358 429140
rect 42548 424418 42604 424427
rect 42604 424376 42686 424404
rect 42548 424353 42604 424362
rect 42356 419978 42412 419987
rect 42356 419913 42412 419922
rect 42370 418507 42398 419913
rect 42356 418498 42412 418507
rect 42356 418433 42358 418442
rect 42410 418433 42412 418442
rect 42358 418401 42410 418407
rect 41986 418308 42398 418336
rect 41782 413427 41834 413433
rect 41782 413369 41834 413375
rect 41782 413205 41834 413211
rect 41782 413147 41834 413153
rect 41794 412624 41822 413147
rect 42370 411509 42398 418308
rect 42454 416535 42506 416541
rect 42454 416477 42506 416483
rect 42358 411503 42410 411509
rect 42358 411445 42410 411451
rect 42466 411380 42494 416477
rect 42166 411355 42218 411361
rect 42166 411297 42218 411303
rect 42370 411352 42494 411380
rect 42178 410805 42206 411297
rect 42178 409733 42206 410182
rect 42166 409727 42218 409733
rect 42166 409669 42218 409675
rect 42370 409511 42398 411352
rect 42658 411232 42686 424376
rect 43124 421014 43180 421023
rect 43124 420949 43180 420958
rect 42934 415425 42986 415431
rect 42934 415367 42986 415373
rect 42562 411204 42686 411232
rect 42562 409881 42590 411204
rect 42550 409875 42602 409881
rect 42550 409817 42602 409823
rect 42550 409727 42602 409733
rect 42550 409669 42602 409675
rect 42166 409505 42218 409511
rect 42166 409447 42218 409453
rect 42358 409505 42410 409511
rect 42358 409447 42410 409453
rect 42178 408965 42206 409447
rect 42358 409357 42410 409363
rect 42358 409299 42410 409305
rect 42166 408247 42218 408253
rect 42166 408189 42218 408195
rect 42178 407769 42206 408189
rect 42070 407507 42122 407513
rect 42070 407449 42122 407455
rect 42082 407148 42110 407449
rect 42370 407069 42398 409299
rect 42166 407063 42218 407069
rect 42166 407005 42218 407011
rect 42358 407063 42410 407069
rect 42358 407005 42410 407011
rect 42178 406482 42206 407005
rect 42068 406362 42124 406371
rect 42068 406297 42124 406306
rect 42082 405929 42110 406297
rect 42562 406107 42590 409669
rect 42946 409363 42974 415367
rect 43030 415203 43082 415209
rect 43030 415145 43082 415151
rect 42934 409357 42986 409363
rect 42934 409299 42986 409305
rect 42934 409209 42986 409215
rect 42934 409151 42986 409157
rect 42550 406101 42602 406107
rect 42550 406043 42602 406049
rect 42164 405178 42220 405187
rect 42164 405113 42220 405122
rect 42178 404646 42206 405113
rect 42178 404632 42302 404646
rect 42192 404618 42302 404632
rect 41794 403707 41822 403997
rect 42166 403881 42218 403887
rect 42166 403823 42218 403829
rect 41780 403698 41836 403707
rect 41780 403633 41836 403642
rect 42178 403448 42206 403823
rect 42166 403363 42218 403369
rect 42166 403305 42218 403311
rect 42178 402782 42206 403305
rect 42274 403263 42302 404618
rect 42946 403369 42974 409151
rect 43042 407513 43070 415145
rect 43138 408253 43166 420949
rect 43234 414913 43262 429112
rect 43222 414907 43274 414913
rect 43222 414849 43274 414855
rect 43702 414907 43754 414913
rect 43702 414849 43754 414855
rect 43222 414759 43274 414765
rect 43222 414701 43274 414707
rect 43126 408247 43178 408253
rect 43126 408189 43178 408195
rect 43030 407507 43082 407513
rect 43030 407449 43082 407455
rect 43234 403887 43262 414701
rect 43222 403881 43274 403887
rect 43222 403823 43274 403829
rect 42934 403363 42986 403369
rect 42934 403305 42986 403311
rect 43714 403263 43742 414849
rect 42260 403254 42316 403263
rect 42260 403189 42316 403198
rect 43508 403254 43564 403263
rect 43508 403189 43564 403198
rect 43700 403254 43756 403263
rect 43700 403189 43756 403198
rect 41780 402662 41836 402671
rect 41780 402597 41836 402606
rect 41794 402157 41822 402597
rect 41780 401922 41836 401931
rect 41780 401857 41836 401866
rect 41794 401598 41822 401857
rect 41780 400146 41836 400155
rect 41780 400081 41836 400090
rect 41794 399748 41822 400081
rect 41780 399554 41836 399563
rect 41780 399489 41836 399498
rect 41794 399121 41822 399489
rect 41780 398814 41836 398823
rect 41780 398749 41836 398758
rect 41794 398490 41822 398749
rect 42358 393965 42410 393971
rect 42356 393930 42358 393939
rect 42410 393930 42412 393939
rect 42356 393865 42412 393874
rect 42646 392929 42698 392935
rect 42644 392894 42646 392903
rect 42698 392894 42700 392903
rect 42644 392829 42700 392838
rect 42358 392337 42410 392343
rect 42356 392302 42358 392311
rect 42410 392302 42412 392311
rect 42356 392237 42412 392246
rect 43220 391266 43276 391275
rect 43220 391201 43276 391210
rect 41972 386678 42028 386687
rect 41972 386613 42028 386622
rect 37268 381202 37324 381211
rect 37268 381137 37324 381146
rect 37282 371623 37310 381137
rect 40148 380462 40204 380471
rect 40148 380397 40204 380406
rect 40052 380018 40108 380027
rect 40052 379953 40108 379962
rect 37364 378834 37420 378843
rect 37364 378769 37420 378778
rect 37378 373251 37406 378769
rect 37366 373245 37418 373251
rect 37366 373187 37418 373193
rect 40066 373103 40094 379953
rect 40054 373097 40106 373103
rect 40054 373039 40106 373045
rect 40162 372585 40190 380397
rect 40244 378094 40300 378103
rect 40244 378029 40300 378038
rect 40150 372579 40202 372585
rect 40150 372521 40202 372527
rect 40258 372289 40286 378029
rect 40246 372283 40298 372289
rect 40246 372225 40298 372231
rect 37270 371617 37322 371623
rect 37270 371559 37322 371565
rect 38326 371617 38378 371623
rect 38326 371559 38378 371565
rect 38338 370555 38366 371559
rect 38324 370546 38380 370555
rect 38324 370481 38380 370490
rect 41986 370217 42014 386613
rect 42356 383570 42412 383579
rect 42356 383505 42412 383514
rect 42260 376614 42316 376623
rect 42260 376549 42316 376558
rect 42274 375291 42302 376549
rect 42260 375282 42316 375291
rect 42260 375217 42262 375226
rect 42314 375217 42316 375226
rect 42262 375185 42314 375191
rect 41974 370211 42026 370217
rect 41974 370153 42026 370159
rect 42370 369995 42398 383505
rect 43124 377798 43180 377807
rect 43124 377733 43180 377742
rect 43030 373097 43082 373103
rect 43030 373039 43082 373045
rect 42838 372579 42890 372585
rect 42838 372521 42890 372527
rect 42166 369989 42218 369995
rect 42166 369931 42218 369937
rect 42358 369989 42410 369995
rect 42358 369931 42410 369937
rect 42178 369445 42206 369931
rect 42358 369841 42410 369847
rect 42358 369783 42410 369789
rect 42370 368145 42398 369783
rect 42070 368139 42122 368145
rect 42070 368081 42122 368087
rect 42358 368139 42410 368145
rect 42358 368081 42410 368087
rect 42082 367632 42110 368081
rect 42070 367399 42122 367405
rect 42070 367341 42122 367347
rect 42082 366966 42110 367341
rect 42850 366295 42878 372521
rect 42934 372283 42986 372289
rect 42934 372225 42986 372231
rect 42070 366289 42122 366295
rect 42070 366231 42122 366237
rect 42838 366289 42890 366295
rect 42838 366231 42890 366237
rect 42082 365782 42110 366231
rect 42166 365031 42218 365037
rect 42166 364973 42218 364979
rect 42178 364569 42206 364973
rect 42070 364291 42122 364297
rect 42070 364233 42122 364239
rect 42082 363932 42110 364233
rect 42946 363705 42974 372225
rect 43042 364297 43070 373039
rect 43138 365037 43166 377733
rect 43126 365031 43178 365037
rect 43126 364973 43178 364979
rect 43030 364291 43082 364297
rect 43030 364233 43082 364239
rect 42166 363699 42218 363705
rect 42166 363641 42218 363647
rect 42934 363699 42986 363705
rect 42934 363641 42986 363647
rect 42178 363266 42206 363641
rect 42068 362850 42124 362859
rect 42068 362785 42124 362794
rect 42082 362748 42110 362785
rect 41876 361962 41932 361971
rect 41876 361897 41932 361906
rect 41890 361416 41918 361897
rect 41794 360639 41822 360824
rect 42166 360665 42218 360671
rect 41780 360630 41836 360639
rect 42166 360607 42218 360613
rect 41780 360565 41836 360574
rect 42178 360232 42206 360607
rect 42260 360186 42316 360195
rect 42260 360121 42316 360130
rect 42274 359615 42302 360121
rect 42192 359587 42302 359615
rect 41780 359446 41836 359455
rect 41780 359381 41836 359390
rect 41794 358974 41822 359381
rect 41780 358706 41836 358715
rect 41780 358641 41836 358650
rect 41794 358382 41822 358641
rect 41780 356930 41836 356939
rect 41780 356865 41836 356874
rect 41794 356565 41822 356865
rect 41780 356486 41836 356495
rect 41780 356421 41836 356430
rect 41794 355940 41822 356421
rect 41780 355598 41836 355607
rect 41780 355533 41836 355542
rect 41794 355274 41822 355533
rect 42358 350749 42410 350755
rect 42356 350714 42358 350723
rect 42410 350714 42412 350723
rect 42356 350649 42412 350658
rect 42358 350009 42410 350015
rect 42356 349974 42358 349983
rect 42410 349974 42412 349983
rect 42356 349909 42412 349918
rect 42358 349121 42410 349127
rect 42356 349086 42358 349095
rect 42410 349086 42412 349095
rect 42356 349021 42412 349030
rect 43234 347763 43262 391201
rect 43522 390979 43550 403189
rect 43508 390970 43564 390979
rect 43508 390905 43564 390914
rect 43318 373245 43370 373251
rect 43318 373187 43370 373193
rect 43330 360671 43358 373187
rect 43318 360665 43370 360671
rect 43318 360607 43370 360613
rect 43220 347754 43276 347763
rect 43220 347689 43276 347698
rect 43220 347606 43276 347615
rect 43220 347541 43276 347550
rect 41876 343610 41932 343619
rect 41876 343545 41932 343554
rect 41780 340354 41836 340363
rect 41780 340289 41836 340298
rect 37364 339910 37420 339919
rect 37364 339845 37420 339854
rect 37172 337394 37228 337403
rect 37172 337329 37228 337338
rect 37186 329813 37214 337329
rect 37378 336515 37406 339845
rect 39956 337986 40012 337995
rect 39956 337921 40012 337930
rect 37364 336506 37420 336515
rect 37364 336441 37420 336450
rect 37364 335618 37420 335627
rect 37364 335553 37420 335562
rect 37174 329807 37226 329813
rect 37174 329749 37226 329755
rect 37378 328481 37406 335553
rect 39970 328555 39998 337921
rect 40052 337246 40108 337255
rect 40052 337181 40108 337190
rect 40066 328851 40094 337181
rect 40244 334878 40300 334887
rect 40244 334813 40300 334822
rect 40054 328845 40106 328851
rect 40054 328787 40106 328793
rect 39958 328549 40010 328555
rect 39958 328491 40010 328497
rect 37366 328475 37418 328481
rect 37366 328417 37418 328423
rect 40258 328407 40286 334813
rect 40246 328401 40298 328407
rect 40246 328343 40298 328349
rect 41794 327075 41822 340289
rect 41890 330701 41918 343545
rect 42548 334434 42604 334443
rect 42548 334369 42604 334378
rect 42260 333546 42316 333555
rect 42260 333481 42316 333490
rect 42274 332075 42302 333481
rect 42260 332066 42316 332075
rect 42260 332001 42262 332010
rect 42314 332001 42316 332010
rect 42262 331969 42314 331975
rect 42562 330868 42590 334369
rect 42562 330840 42686 330868
rect 41878 330695 41930 330701
rect 41878 330637 41930 330643
rect 42550 330695 42602 330701
rect 42550 330637 42602 330643
rect 41782 327069 41834 327075
rect 41782 327011 41834 327017
rect 41782 326773 41834 326779
rect 41782 326715 41834 326721
rect 41794 326266 41822 326715
rect 42562 324929 42590 330637
rect 42070 324923 42122 324929
rect 42070 324865 42122 324871
rect 42550 324923 42602 324929
rect 42550 324865 42602 324871
rect 42082 324416 42110 324865
rect 42658 324652 42686 330840
rect 43126 329807 43178 329813
rect 43126 329749 43178 329755
rect 42934 328845 42986 328851
rect 42934 328787 42986 328793
rect 42838 328401 42890 328407
rect 42838 328343 42890 328349
rect 42562 324624 42686 324652
rect 42166 324183 42218 324189
rect 42166 324125 42218 324131
rect 42178 323750 42206 324125
rect 42166 323147 42218 323153
rect 42166 323089 42218 323095
rect 42178 322566 42206 323089
rect 42562 321821 42590 324624
rect 42070 321815 42122 321821
rect 42070 321757 42122 321763
rect 42550 321815 42602 321821
rect 42550 321757 42602 321763
rect 42082 321382 42110 321757
rect 42166 321075 42218 321081
rect 42166 321017 42218 321023
rect 42178 320716 42206 321017
rect 42850 320637 42878 328343
rect 42946 321081 42974 328787
rect 43030 328475 43082 328481
rect 43030 328417 43082 328423
rect 42934 321075 42986 321081
rect 42934 321017 42986 321023
rect 42934 320927 42986 320933
rect 42934 320869 42986 320875
rect 42166 320631 42218 320637
rect 42166 320573 42218 320579
rect 42838 320631 42890 320637
rect 42838 320573 42890 320579
rect 42178 320081 42206 320573
rect 42068 319782 42124 319791
rect 42068 319717 42124 319726
rect 42082 319532 42110 319717
rect 42262 318781 42314 318787
rect 41876 318746 41932 318755
rect 42262 318723 42314 318729
rect 41876 318681 41932 318690
rect 41890 318241 41918 318681
rect 41780 317858 41836 317867
rect 41780 317793 41836 317802
rect 41794 317608 41822 317793
rect 42274 317059 42302 318723
rect 42192 317031 42302 317059
rect 42946 316641 42974 320869
rect 43042 318787 43070 328417
rect 43138 323153 43166 329749
rect 43126 323147 43178 323153
rect 43126 323089 43178 323095
rect 43030 318781 43082 318787
rect 43030 318723 43082 318729
rect 42070 316635 42122 316641
rect 42070 316577 42122 316583
rect 42934 316635 42986 316641
rect 42934 316577 42986 316583
rect 42082 316424 42110 316577
rect 41780 316082 41836 316091
rect 41780 316017 41836 316026
rect 41794 315758 41822 316017
rect 41780 315490 41836 315499
rect 41780 315425 41836 315434
rect 41794 315205 41822 315425
rect 41876 313714 41932 313723
rect 41876 313649 41932 313658
rect 41890 313390 41918 313649
rect 41780 313270 41836 313279
rect 41780 313205 41836 313214
rect 41794 312724 41822 313205
rect 41780 312382 41836 312391
rect 41780 312317 41836 312326
rect 41794 312058 41822 312317
rect 42358 307533 42410 307539
rect 42356 307498 42358 307507
rect 42410 307498 42412 307507
rect 42356 307433 42412 307442
rect 42358 306793 42410 306799
rect 42356 306758 42358 306767
rect 42410 306758 42412 306767
rect 42356 306693 42412 306702
rect 42358 305535 42410 305541
rect 42358 305477 42410 305483
rect 42370 305435 42398 305477
rect 42356 305426 42412 305435
rect 42356 305361 42412 305370
rect 43234 304103 43262 347541
rect 43318 328549 43370 328555
rect 43318 328491 43370 328497
rect 43330 320933 43358 328491
rect 43318 320927 43370 320933
rect 43318 320869 43370 320875
rect 43220 304094 43276 304103
rect 43220 304029 43276 304038
rect 43220 303946 43276 303955
rect 43220 303881 43276 303890
rect 41876 300394 41932 300403
rect 41876 300329 41932 300338
rect 37364 296694 37420 296703
rect 37364 296629 37420 296638
rect 37268 294030 37324 294039
rect 37268 293965 37324 293974
rect 37282 286819 37310 293965
rect 37378 292411 37406 296629
rect 40052 294770 40108 294779
rect 40052 294705 40108 294714
rect 37364 292402 37420 292411
rect 37364 292337 37420 292346
rect 37270 286813 37322 286819
rect 37270 286755 37322 286761
rect 40066 285339 40094 294705
rect 40148 294030 40204 294039
rect 40148 293965 40204 293974
rect 40054 285333 40106 285339
rect 40054 285275 40106 285281
rect 40162 285265 40190 293965
rect 40244 291662 40300 291671
rect 40244 291597 40300 291606
rect 40150 285259 40202 285265
rect 40150 285201 40202 285207
rect 40258 285191 40286 291597
rect 41782 289847 41834 289853
rect 41782 289789 41834 289795
rect 40534 286813 40586 286819
rect 40534 286755 40586 286761
rect 40246 285185 40298 285191
rect 40246 285127 40298 285133
rect 40546 284123 40574 286755
rect 40532 284114 40588 284123
rect 40532 284049 40588 284058
rect 41794 283859 41822 289789
rect 41890 285432 41918 300329
rect 42260 297286 42316 297295
rect 42260 297221 42316 297230
rect 42274 289853 42302 297221
rect 42452 292402 42508 292411
rect 42452 292337 42508 292346
rect 42262 289847 42314 289853
rect 42262 289789 42314 289795
rect 42260 288850 42316 288859
rect 42260 288785 42316 288794
rect 42274 288077 42302 288785
rect 42262 288071 42314 288077
rect 42262 288013 42314 288019
rect 41890 285404 42398 285432
rect 42262 285333 42314 285339
rect 42262 285275 42314 285281
rect 41782 283853 41834 283859
rect 41782 283795 41834 283801
rect 41782 283557 41834 283563
rect 41782 283499 41834 283505
rect 41794 283050 41822 283499
rect 42274 283383 42302 285275
rect 42260 283374 42316 283383
rect 42260 283309 42316 283318
rect 42370 281787 42398 285404
rect 42466 282495 42494 292337
rect 42932 291366 42988 291375
rect 42932 291301 42988 291310
rect 42452 282486 42508 282495
rect 42452 282421 42508 282430
rect 42166 281781 42218 281787
rect 42166 281723 42218 281729
rect 42358 281781 42410 281787
rect 42358 281723 42410 281729
rect 42178 281200 42206 281723
rect 42082 280159 42110 280534
rect 42070 280153 42122 280159
rect 42070 280095 42122 280101
rect 42358 280153 42410 280159
rect 42358 280095 42410 280101
rect 41780 279822 41836 279831
rect 41780 279757 41836 279766
rect 41794 279350 41822 279757
rect 42166 278599 42218 278605
rect 42166 278541 42218 278547
rect 42178 278166 42206 278541
rect 42166 277859 42218 277865
rect 42166 277801 42218 277807
rect 42178 277500 42206 277801
rect 42070 277415 42122 277421
rect 42070 277357 42122 277363
rect 42082 276908 42110 277357
rect 41780 276566 41836 276575
rect 41780 276501 41836 276510
rect 41794 276316 41822 276501
rect 42370 276459 42398 280095
rect 42946 278605 42974 291301
rect 43126 285259 43178 285265
rect 43126 285201 43178 285207
rect 43030 285185 43082 285191
rect 43030 285127 43082 285133
rect 42934 278599 42986 278605
rect 42934 278541 42986 278547
rect 43042 277421 43070 285127
rect 43138 277865 43166 285201
rect 43126 277859 43178 277865
rect 43126 277801 43178 277807
rect 43030 277415 43082 277421
rect 43030 277357 43082 277363
rect 42358 276453 42410 276459
rect 42358 276395 42410 276401
rect 41972 275530 42028 275539
rect 41972 275465 42028 275474
rect 41986 275058 42014 275465
rect 41780 274938 41836 274947
rect 41780 274873 41836 274882
rect 41794 274392 41822 274873
rect 42164 274198 42220 274207
rect 42164 274133 42220 274142
rect 42178 273845 42206 274133
rect 42260 273754 42316 273763
rect 42260 273689 42316 273698
rect 42274 273222 42302 273689
rect 42192 273194 42302 273222
rect 41780 273014 41836 273023
rect 41780 272949 41836 272958
rect 41794 272542 41822 272949
rect 41780 272274 41836 272283
rect 41780 272209 41836 272218
rect 41794 272024 41822 272209
rect 41780 270646 41836 270655
rect 41780 270581 41836 270590
rect 41794 270174 41822 270581
rect 42548 270498 42604 270507
rect 42548 270433 42604 270442
rect 41780 270054 41836 270063
rect 41780 269989 41836 269998
rect 41794 269508 41822 269989
rect 41780 269166 41836 269175
rect 41780 269101 41836 269110
rect 41794 268877 41822 269101
rect 42562 267820 42590 270433
rect 42562 267792 42782 267820
rect 42262 264317 42314 264323
rect 42260 264282 42262 264291
rect 42314 264282 42316 264291
rect 42260 264217 42316 264226
rect 42646 263281 42698 263287
rect 42644 263246 42646 263255
rect 42698 263246 42700 263255
rect 42644 263181 42700 263190
rect 42644 262506 42700 262515
rect 42644 262441 42700 262450
rect 42658 262325 42686 262441
rect 42646 262319 42698 262325
rect 42646 262261 42698 262267
rect 41300 259546 41356 259555
rect 41300 259481 41356 259490
rect 40244 251554 40300 251563
rect 40244 251489 40300 251498
rect 37364 250814 37420 250823
rect 37364 250749 37420 250758
rect 40052 250814 40108 250823
rect 40052 250749 40108 250758
rect 37378 241975 37406 250749
rect 40066 242123 40094 250749
rect 40148 248446 40204 248455
rect 40148 248381 40204 248390
rect 40054 242117 40106 242123
rect 40054 242059 40106 242065
rect 40162 242049 40190 248381
rect 40258 242091 40286 251489
rect 41314 246119 41342 259481
rect 42068 257178 42124 257187
rect 42068 257113 42124 257122
rect 41780 254366 41836 254375
rect 41780 254301 41836 254310
rect 41302 246113 41354 246119
rect 41302 246055 41354 246061
rect 40244 242082 40300 242091
rect 40150 242043 40202 242049
rect 40244 242017 40300 242026
rect 40150 241985 40202 241991
rect 37366 241969 37418 241975
rect 37366 241911 37418 241917
rect 41794 240643 41822 254301
rect 42082 244417 42110 257113
rect 42754 249912 42782 267792
rect 43234 260887 43262 303881
rect 43508 261618 43564 261627
rect 43508 261553 43564 261562
rect 43220 260878 43276 260887
rect 43220 260813 43276 260822
rect 43412 259398 43468 259407
rect 43412 259333 43468 259342
rect 42658 249893 42782 249912
rect 42166 249887 42218 249893
rect 42166 249829 42218 249835
rect 42646 249887 42782 249893
rect 42698 249884 42782 249887
rect 42646 249829 42698 249835
rect 42178 247123 42206 249829
rect 42548 249186 42604 249195
rect 42548 249121 42604 249130
rect 42164 247114 42220 247123
rect 42164 247049 42220 247058
rect 42356 246818 42412 246827
rect 42356 246753 42412 246762
rect 42370 245643 42398 246753
rect 42562 245916 42590 249121
rect 43028 247558 43084 247567
rect 43028 247493 43084 247502
rect 42562 245888 42686 245916
rect 42356 245634 42412 245643
rect 42356 245569 42412 245578
rect 42370 245009 42398 245569
rect 42358 245003 42410 245009
rect 42358 244945 42410 244951
rect 42070 244411 42122 244417
rect 42070 244353 42122 244359
rect 42550 244411 42602 244417
rect 42550 244353 42602 244359
rect 42358 242117 42410 242123
rect 42358 242059 42410 242065
rect 41782 240637 41834 240643
rect 41782 240579 41834 240585
rect 41782 240415 41834 240421
rect 41782 240357 41834 240363
rect 41794 239834 41822 240357
rect 42370 239427 42398 242059
rect 42356 239418 42412 239427
rect 42562 239385 42590 244353
rect 42356 239353 42412 239362
rect 42550 239379 42602 239385
rect 42550 239321 42602 239327
rect 42358 239305 42410 239311
rect 42658 239256 42686 245888
rect 42934 241969 42986 241975
rect 42934 241911 42986 241917
rect 42358 239247 42410 239253
rect 42370 238571 42398 239247
rect 42562 239237 42686 239256
rect 42550 239231 42686 239237
rect 42602 239228 42686 239231
rect 42550 239173 42602 239179
rect 42452 238974 42508 238983
rect 42452 238909 42508 238918
rect 42166 238565 42218 238571
rect 42166 238507 42218 238513
rect 42358 238565 42410 238571
rect 42358 238507 42410 238513
rect 42178 237984 42206 238507
rect 42466 238368 42494 238909
rect 42370 238340 42494 238368
rect 42166 237899 42218 237905
rect 42166 237841 42218 237847
rect 42178 237361 42206 237841
rect 42166 236715 42218 236721
rect 42166 236657 42218 236663
rect 42178 236165 42206 236657
rect 42166 235457 42218 235463
rect 42166 235399 42218 235405
rect 42178 234950 42206 235399
rect 42370 234871 42398 238340
rect 42946 236721 42974 241911
rect 42934 236715 42986 236721
rect 42934 236657 42986 236663
rect 43042 235463 43070 247493
rect 43318 246113 43370 246119
rect 43318 246055 43370 246061
rect 43126 242043 43178 242049
rect 43126 241985 43178 241991
rect 43030 235457 43082 235463
rect 43030 235399 43082 235405
rect 42166 234865 42218 234871
rect 42166 234807 42218 234813
rect 42358 234865 42410 234871
rect 42358 234807 42410 234813
rect 42178 234325 42206 234807
rect 43138 234205 43166 241985
rect 43222 239231 43274 239237
rect 43222 239173 43274 239179
rect 42070 234199 42122 234205
rect 42070 234141 42122 234147
rect 43126 234199 43178 234205
rect 43126 234141 43178 234147
rect 42082 233692 42110 234141
rect 41780 233350 41836 233359
rect 41780 233285 41836 233294
rect 41794 233129 41822 233285
rect 43234 232577 43262 239173
rect 42262 232571 42314 232577
rect 42262 232513 42314 232519
rect 43222 232571 43274 232577
rect 43222 232513 43274 232519
rect 41986 231731 42014 231842
rect 41972 231722 42028 231731
rect 41972 231657 42028 231666
rect 41986 230991 42014 231176
rect 41972 230982 42028 230991
rect 41972 230917 42028 230926
rect 42274 230672 42302 232513
rect 42192 230644 42302 230672
rect 41780 230390 41836 230399
rect 41780 230325 41836 230334
rect 41794 229992 41822 230325
rect 41780 229798 41836 229807
rect 41780 229733 41836 229742
rect 41794 229357 41822 229733
rect 41780 229058 41836 229067
rect 41780 228993 41836 229002
rect 41794 228808 41822 228993
rect 43222 227613 43274 227619
rect 43222 227555 43274 227561
rect 41780 227282 41836 227291
rect 41780 227217 41836 227226
rect 41794 226958 41822 227217
rect 41780 226690 41836 226699
rect 41780 226625 41836 226634
rect 41794 226321 41822 226625
rect 42068 226246 42124 226255
rect 42068 226181 42124 226190
rect 42082 225700 42110 226181
rect 42358 221101 42410 221107
rect 42356 221066 42358 221075
rect 42410 221066 42412 221075
rect 42356 221001 42412 221010
rect 42358 220361 42410 220367
rect 42356 220326 42358 220335
rect 42410 220326 42412 220335
rect 42356 220261 42412 220270
rect 42358 219473 42410 219479
rect 42356 219438 42358 219447
rect 42410 219438 42412 219447
rect 42356 219373 42412 219382
rect 43234 217671 43262 227555
rect 43220 217662 43276 217671
rect 43220 217597 43276 217606
rect 43330 216931 43358 246055
rect 43426 246045 43454 259333
rect 43414 246039 43466 246045
rect 43414 245981 43466 245987
rect 43316 216922 43372 216931
rect 43316 216857 43372 216866
rect 43426 216191 43454 245981
rect 43522 227619 43550 261553
rect 44578 255147 44606 544793
rect 44566 255141 44618 255147
rect 44566 255083 44618 255089
rect 44674 246415 44702 930925
rect 44770 627959 44798 988201
rect 44854 988185 44906 988191
rect 44854 988127 44906 988133
rect 44866 673765 44894 988127
rect 44950 988111 45002 988117
rect 44950 988053 45002 988059
rect 44962 714317 44990 988053
rect 45046 988037 45098 988043
rect 45046 987979 45098 987985
rect 45058 757533 45086 987979
rect 45142 987963 45194 987969
rect 45142 987905 45194 987911
rect 45154 800675 45182 987905
rect 47446 986557 47498 986563
rect 47446 986499 47498 986505
rect 46102 959103 46154 959109
rect 46102 959045 46154 959051
rect 46114 947935 46142 959045
rect 46102 947929 46154 947935
rect 46102 947871 46154 947877
rect 47458 946275 47486 986499
rect 47444 946266 47500 946275
rect 47444 946201 47500 946210
rect 47542 872671 47594 872677
rect 47542 872613 47594 872619
rect 47446 858315 47498 858321
rect 47446 858257 47498 858263
rect 45142 800669 45194 800675
rect 45142 800611 45194 800617
rect 45046 757527 45098 757533
rect 45046 757469 45098 757475
rect 44950 714311 45002 714317
rect 44950 714253 45002 714259
rect 44854 673759 44906 673765
rect 44854 673701 44906 673707
rect 44758 627953 44810 627959
rect 44758 627895 44810 627901
rect 44758 486761 44810 486767
rect 44758 486703 44810 486709
rect 44770 392343 44798 486703
rect 44854 472405 44906 472411
rect 44854 472347 44906 472353
rect 44866 393971 44894 472347
rect 45046 414759 45098 414765
rect 45046 414701 45098 414707
rect 44854 393965 44906 393971
rect 44854 393907 44906 393913
rect 44758 392337 44810 392343
rect 44758 392279 44810 392285
rect 44950 385973 45002 385979
rect 44950 385915 45002 385921
rect 44758 375243 44810 375249
rect 44758 375185 44810 375191
rect 44662 246409 44714 246415
rect 44662 246351 44714 246357
rect 44770 246341 44798 375185
rect 44854 313971 44906 313977
rect 44854 313913 44906 313919
rect 44758 246335 44810 246341
rect 44758 246277 44810 246283
rect 44566 241969 44618 241975
rect 44566 241911 44618 241917
rect 43510 227613 43562 227619
rect 43510 227555 43562 227561
rect 43412 216182 43468 216191
rect 43412 216117 43468 216126
rect 41972 213962 42028 213971
rect 41972 213897 42028 213906
rect 40244 210854 40300 210863
rect 40244 210789 40300 210798
rect 40052 207154 40108 207163
rect 40052 207089 40108 207098
rect 37364 206118 37420 206127
rect 37364 206053 37420 206062
rect 37378 198833 37406 206053
rect 40066 201497 40094 207089
rect 40148 205230 40204 205239
rect 40148 205165 40204 205174
rect 40054 201491 40106 201497
rect 40054 201433 40106 201439
rect 37366 198827 37418 198833
rect 37366 198769 37418 198775
rect 40162 198759 40190 205165
rect 40258 201571 40286 210789
rect 40246 201565 40298 201571
rect 40246 201507 40298 201513
rect 41782 201565 41834 201571
rect 41782 201507 41834 201513
rect 40150 198753 40202 198759
rect 40918 198753 40970 198759
rect 40150 198695 40202 198701
rect 40916 198718 40918 198727
rect 40970 198718 40972 198727
rect 40916 198653 40972 198662
rect 41794 197427 41822 201507
rect 41986 201127 42014 213897
rect 42068 209226 42124 209235
rect 42068 209161 42124 209170
rect 41974 201121 42026 201127
rect 41974 201063 42026 201069
rect 42082 197501 42110 209161
rect 42836 208930 42892 208939
rect 42836 208865 42892 208874
rect 42356 207894 42412 207903
rect 42356 207829 42412 207838
rect 42370 204531 42398 207829
rect 42358 204525 42410 204531
rect 42358 204467 42410 204473
rect 42358 204377 42410 204383
rect 42356 204342 42358 204351
rect 42410 204342 42412 204351
rect 42356 204277 42412 204286
rect 42370 202871 42398 204277
rect 42356 202862 42412 202871
rect 42356 202797 42412 202806
rect 42166 201491 42218 201497
rect 42166 201433 42218 201439
rect 42178 197543 42206 201433
rect 42358 201121 42410 201127
rect 42358 201063 42410 201069
rect 42164 197534 42220 197543
rect 42070 197495 42122 197501
rect 42164 197469 42220 197478
rect 42070 197437 42122 197443
rect 41782 197421 41834 197427
rect 41782 197363 41834 197369
rect 41782 197199 41834 197205
rect 41782 197141 41834 197147
rect 41794 196618 41822 197141
rect 42370 195355 42398 201063
rect 42850 195799 42878 208865
rect 43124 204934 43180 204943
rect 43124 204869 43180 204878
rect 43030 204525 43082 204531
rect 43030 204467 43082 204473
rect 42934 197495 42986 197501
rect 42934 197437 42986 197443
rect 42550 195793 42602 195799
rect 42838 195793 42890 195799
rect 42602 195753 42686 195781
rect 42550 195735 42602 195741
rect 42166 195349 42218 195355
rect 42166 195291 42218 195297
rect 42358 195349 42410 195355
rect 42358 195291 42410 195297
rect 42178 194805 42206 195291
rect 42356 195166 42412 195175
rect 42356 195101 42412 195110
rect 42070 194535 42122 194541
rect 42070 194477 42122 194483
rect 42082 194176 42110 194477
rect 42070 193499 42122 193505
rect 42070 193441 42122 193447
rect 42082 192992 42110 193441
rect 42166 192241 42218 192247
rect 42166 192183 42218 192189
rect 42178 191769 42206 192183
rect 42370 191507 42398 195101
rect 42070 191501 42122 191507
rect 42070 191443 42122 191449
rect 42358 191501 42410 191507
rect 42358 191443 42410 191449
rect 42082 191142 42110 191443
rect 41780 191022 41836 191031
rect 41780 190957 41836 190966
rect 41794 190476 41822 190957
rect 41780 190134 41836 190143
rect 41780 190069 41836 190078
rect 41794 189929 41822 190069
rect 41972 189098 42028 189107
rect 41972 189033 42028 189042
rect 41986 188626 42014 189033
rect 41780 188358 41836 188367
rect 41780 188293 41836 188302
rect 41794 188011 41822 188293
rect 41794 187997 42302 188011
rect 41808 187983 42302 187997
rect 42166 187727 42218 187733
rect 42166 187669 42218 187675
rect 42178 187442 42206 187669
rect 42274 187308 42302 187983
rect 42274 187280 42398 187308
rect 42262 187209 42314 187215
rect 42262 187151 42314 187157
rect 42166 187135 42218 187141
rect 42166 187077 42218 187083
rect 42178 186776 42206 187077
rect 42178 186124 42206 186184
rect 42274 186124 42302 187151
rect 42178 186096 42302 186124
rect 41780 185990 41836 185999
rect 41780 185925 41836 185934
rect 41794 185592 41822 185925
rect 42370 184792 42398 187280
rect 42550 187135 42602 187141
rect 42658 187123 42686 195753
rect 42838 195735 42890 195741
rect 42838 195645 42890 195651
rect 42838 195587 42890 195593
rect 42850 187733 42878 195587
rect 42838 187727 42890 187733
rect 42838 187669 42890 187675
rect 42946 187289 42974 197437
rect 43042 193505 43070 204467
rect 43030 193499 43082 193505
rect 43030 193441 43082 193447
rect 43138 192247 43166 204869
rect 44578 204383 44606 241911
rect 44866 219479 44894 313913
rect 44962 307539 44990 385915
rect 45058 350015 45086 414701
rect 47458 367405 47486 858257
rect 47554 823171 47582 872613
rect 47542 823165 47594 823171
rect 47542 823107 47594 823113
rect 47542 786313 47594 786319
rect 47542 786255 47594 786261
rect 47554 735703 47582 786255
rect 47542 735697 47594 735703
rect 47542 735639 47594 735645
rect 47542 728667 47594 728673
rect 47542 728609 47594 728615
rect 47554 692783 47582 728609
rect 47542 692777 47594 692783
rect 47542 692719 47594 692725
rect 47542 685525 47594 685531
rect 47542 685467 47594 685473
rect 47446 367399 47498 367405
rect 47446 367341 47498 367347
rect 45046 350009 45098 350015
rect 45046 349951 45098 349957
rect 45046 332027 45098 332033
rect 45046 331969 45098 331975
rect 44950 307533 45002 307539
rect 44950 307475 45002 307481
rect 44950 299615 45002 299621
rect 44950 299557 45002 299563
rect 44962 221107 44990 299557
rect 45058 252039 45086 331969
rect 45142 285185 45194 285191
rect 45142 285127 45194 285133
rect 45046 252033 45098 252039
rect 45046 251975 45098 251981
rect 44950 221101 45002 221107
rect 44950 221043 45002 221049
rect 45154 220367 45182 285127
rect 47554 237905 47582 685467
rect 47650 584743 47678 988275
rect 47926 986705 47978 986711
rect 47926 986647 47978 986653
rect 47734 986631 47786 986637
rect 47734 986573 47786 986579
rect 47746 946127 47774 986573
rect 47732 946118 47788 946127
rect 47732 946053 47788 946062
rect 47938 944795 47966 986647
rect 59444 975422 59500 975431
rect 59444 975357 59500 975366
rect 59458 973539 59486 975357
rect 50518 973533 50570 973539
rect 50518 973475 50570 973481
rect 59446 973533 59498 973539
rect 59446 973475 59498 973481
rect 47924 944786 47980 944795
rect 47924 944721 47980 944730
rect 50326 901531 50378 901537
rect 50326 901473 50378 901479
rect 47734 829529 47786 829535
rect 47734 829471 47786 829477
rect 47746 780473 47774 829471
rect 50338 822283 50366 901473
rect 50326 822277 50378 822283
rect 50326 822219 50378 822225
rect 50422 815099 50474 815105
rect 50422 815041 50474 815047
rect 50326 800669 50378 800675
rect 50326 800611 50378 800617
rect 47734 780467 47786 780473
rect 47734 780409 47786 780415
rect 47638 584737 47690 584743
rect 47638 584679 47690 584685
rect 48886 563499 48938 563505
rect 48886 563441 48938 563447
rect 48898 544709 48926 563441
rect 48886 544703 48938 544709
rect 48886 544645 48938 544651
rect 47638 501191 47690 501197
rect 47638 501133 47690 501139
rect 47650 436299 47678 501133
rect 47638 436293 47690 436299
rect 47638 436235 47690 436241
rect 47638 429189 47690 429195
rect 47638 429131 47690 429137
rect 47650 350755 47678 429131
rect 47734 371617 47786 371623
rect 47734 371559 47786 371565
rect 47638 350749 47690 350755
rect 47638 350691 47690 350697
rect 47746 306799 47774 371559
rect 50338 324189 50366 800611
rect 50434 779733 50462 815041
rect 50422 779727 50474 779733
rect 50422 779669 50474 779675
rect 50422 714311 50474 714317
rect 50422 714253 50474 714259
rect 50434 694041 50462 714253
rect 50422 694035 50474 694041
rect 50422 693977 50474 693983
rect 50422 671095 50474 671101
rect 50422 671037 50474 671043
rect 50434 649567 50462 671037
rect 50422 649561 50474 649567
rect 50422 649503 50474 649509
rect 50422 627879 50474 627885
rect 50422 627821 50474 627827
rect 50326 324183 50378 324189
rect 50326 324125 50378 324131
rect 47734 306793 47786 306799
rect 47734 306735 47786 306741
rect 47542 237899 47594 237905
rect 47542 237841 47594 237847
rect 45142 220361 45194 220367
rect 45142 220303 45194 220309
rect 44854 219473 44906 219479
rect 44854 219415 44906 219421
rect 44566 204377 44618 204383
rect 44566 204319 44618 204325
rect 43222 198827 43274 198833
rect 43222 198769 43274 198775
rect 43234 195651 43262 198769
rect 43222 195645 43274 195651
rect 43222 195587 43274 195593
rect 50434 194541 50462 627821
rect 50530 541527 50558 973475
rect 61858 962111 61886 993825
rect 62036 992146 62092 992155
rect 62036 992081 62092 992090
rect 62050 962259 62078 992081
rect 69154 987988 69182 995083
rect 77314 993667 77342 995508
rect 77698 993815 77726 995522
rect 77686 993809 77738 993815
rect 77686 993751 77738 993757
rect 78370 993741 78398 995522
rect 80194 993783 80222 995522
rect 80770 995263 80798 995522
rect 82032 995517 82334 995536
rect 82032 995511 82346 995517
rect 82032 995508 82294 995511
rect 82294 995453 82346 995459
rect 80756 995254 80812 995263
rect 82594 995221 82622 995522
rect 83232 995508 83486 995536
rect 80756 995189 80812 995198
rect 82582 995215 82634 995221
rect 82582 995157 82634 995163
rect 82594 993889 82622 995157
rect 82582 993883 82634 993889
rect 82582 993825 82634 993831
rect 80180 993774 80236 993783
rect 78358 993735 78410 993741
rect 80180 993709 80236 993718
rect 78358 993677 78410 993683
rect 77302 993661 77354 993667
rect 83458 993635 83486 995508
rect 84514 993931 84542 995522
rect 85104 995508 85406 995536
rect 86352 995508 86516 995536
rect 85378 995411 85406 995508
rect 92770 995517 92798 999449
rect 92854 999433 92906 999439
rect 92854 999375 92906 999381
rect 86516 995485 86572 995494
rect 92758 995511 92810 995517
rect 92758 995453 92810 995459
rect 85364 995402 85420 995411
rect 85364 995337 85420 995346
rect 84500 993922 84556 993931
rect 84500 993857 84556 993866
rect 92866 993635 92894 999375
rect 77302 993603 77354 993609
rect 83444 993626 83500 993635
rect 83444 993561 83500 993570
rect 92852 993626 92908 993635
rect 92852 993561 92908 993570
rect 89590 990553 89642 990559
rect 89590 990495 89642 990501
rect 73462 989295 73514 989301
rect 73462 989237 73514 989243
rect 69058 987960 69182 987988
rect 63286 986483 63338 986489
rect 63286 986425 63338 986431
rect 62036 962250 62092 962259
rect 62036 962185 62092 962194
rect 61844 962102 61900 962111
rect 61844 962037 61900 962046
rect 59540 960918 59596 960927
rect 59540 960853 59596 960862
rect 59554 959109 59582 960853
rect 59542 959103 59594 959109
rect 59542 959045 59594 959051
rect 53206 948447 53258 948453
rect 53206 948389 53258 948395
rect 53218 933135 53246 948389
rect 57814 947485 57866 947491
rect 57814 947427 57866 947433
rect 57826 946719 57854 947427
rect 57812 946710 57868 946719
rect 57812 946645 57868 946654
rect 53206 933129 53258 933135
rect 53206 933071 53258 933077
rect 59542 933129 59594 933135
rect 59542 933071 59594 933077
rect 59554 932363 59582 933071
rect 59540 932354 59596 932363
rect 59540 932289 59596 932298
rect 59540 917850 59596 917859
rect 59540 917785 59596 917794
rect 59554 915893 59582 917785
rect 53398 915887 53450 915893
rect 53398 915829 53450 915835
rect 59542 915887 59594 915893
rect 59542 915829 59594 915835
rect 53206 887175 53258 887181
rect 53206 887117 53258 887123
rect 53218 823911 53246 887117
rect 53302 843885 53354 843891
rect 53302 843827 53354 843833
rect 53206 823905 53258 823911
rect 53206 823847 53258 823853
rect 53206 805479 53258 805485
rect 53206 805421 53258 805427
rect 51862 649783 51914 649789
rect 51862 649725 51914 649731
rect 51874 644535 51902 649725
rect 51862 644529 51914 644535
rect 51862 644471 51914 644477
rect 51862 607751 51914 607757
rect 51862 607693 51914 607699
rect 51874 601911 51902 607693
rect 51862 601905 51914 601911
rect 51862 601847 51914 601853
rect 51862 564535 51914 564541
rect 51862 564477 51914 564483
rect 51874 561581 51902 564477
rect 51862 561575 51914 561581
rect 51862 561517 51914 561523
rect 50518 541521 50570 541527
rect 50518 541463 50570 541469
rect 50518 457975 50570 457981
rect 50518 457917 50570 457923
rect 50530 392935 50558 457917
rect 50518 392929 50570 392935
rect 50518 392871 50570 392877
rect 50518 342831 50570 342837
rect 50518 342773 50570 342779
rect 50530 264323 50558 342773
rect 50518 264317 50570 264323
rect 50518 264259 50570 264265
rect 53218 246489 53246 805421
rect 53314 778919 53342 843827
rect 53302 778913 53354 778919
rect 53302 778855 53354 778861
rect 53302 761967 53354 761973
rect 53302 761909 53354 761915
rect 53314 246563 53342 761909
rect 53410 406107 53438 915829
rect 59540 903494 59596 903503
rect 59540 903429 59596 903438
rect 59554 901537 59582 903429
rect 59542 901531 59594 901537
rect 59542 901473 59594 901479
rect 59540 889138 59596 889147
rect 59540 889073 59596 889082
rect 59554 887181 59582 889073
rect 59542 887175 59594 887181
rect 59542 887117 59594 887123
rect 59540 874782 59596 874791
rect 59540 874717 59596 874726
rect 59554 872677 59582 874717
rect 59542 872671 59594 872677
rect 59542 872613 59594 872619
rect 58580 860426 58636 860435
rect 58580 860361 58636 860370
rect 58594 858321 58622 860361
rect 58582 858315 58634 858321
rect 58582 858257 58634 858263
rect 59540 846070 59596 846079
rect 59540 846005 59596 846014
rect 59554 843891 59582 846005
rect 59542 843885 59594 843891
rect 59542 843827 59594 843833
rect 59540 831714 59596 831723
rect 59540 831649 59596 831658
rect 59554 829535 59582 831649
rect 59542 829529 59594 829535
rect 59542 829471 59594 829477
rect 59540 817358 59596 817367
rect 59540 817293 59596 817302
rect 59554 815105 59582 817293
rect 59542 815099 59594 815105
rect 59542 815041 59594 815047
rect 59540 802854 59596 802863
rect 59540 802789 59596 802798
rect 59554 800675 59582 802789
rect 59542 800669 59594 800675
rect 59542 800611 59594 800617
rect 59540 788646 59596 788655
rect 59540 788581 59596 788590
rect 59554 786319 59582 788581
rect 59542 786313 59594 786319
rect 59542 786255 59594 786261
rect 59540 774142 59596 774151
rect 59540 774077 59596 774086
rect 59554 771889 59582 774077
rect 53494 771883 53546 771889
rect 53494 771825 53546 771831
rect 59542 771883 59594 771889
rect 59542 771825 59594 771831
rect 53506 737257 53534 771825
rect 59540 759786 59596 759795
rect 59540 759721 59596 759730
rect 59554 757533 59582 759721
rect 53686 757527 53738 757533
rect 53686 757469 53738 757475
rect 59542 757527 59594 757533
rect 59542 757469 59594 757475
rect 53590 743097 53642 743103
rect 53590 743039 53642 743045
rect 53494 737251 53546 737257
rect 53494 737193 53546 737199
rect 53494 718751 53546 718757
rect 53494 718693 53546 718699
rect 53398 406101 53450 406107
rect 53398 406043 53450 406049
rect 53398 328401 53450 328407
rect 53398 328343 53450 328349
rect 53410 263287 53438 328343
rect 53398 263281 53450 263287
rect 53398 263223 53450 263229
rect 53506 246785 53534 718693
rect 53602 276459 53630 743039
rect 53698 736739 53726 757469
rect 59540 745578 59596 745587
rect 59540 745513 59596 745522
rect 59554 743103 59582 745513
rect 59542 743097 59594 743103
rect 59542 743039 59594 743045
rect 53686 736733 53738 736739
rect 53686 736675 53738 736681
rect 59540 731074 59596 731083
rect 59540 731009 59596 731018
rect 59554 728673 59582 731009
rect 59542 728667 59594 728673
rect 59542 728609 59594 728615
rect 59540 716718 59596 716727
rect 59540 716653 59596 716662
rect 59554 714317 59582 716653
rect 59542 714311 59594 714317
rect 59542 714253 59594 714259
rect 59540 702362 59596 702371
rect 59540 702297 59596 702306
rect 59554 699887 59582 702297
rect 59542 699881 59594 699887
rect 59542 699823 59594 699829
rect 59540 688006 59596 688015
rect 59540 687941 59596 687950
rect 59554 685531 59582 687941
rect 59542 685525 59594 685531
rect 59542 685467 59594 685473
rect 53686 675831 53738 675837
rect 53686 675773 53738 675779
rect 53590 276453 53642 276459
rect 53590 276395 53642 276401
rect 53494 246779 53546 246785
rect 53494 246721 53546 246727
rect 53698 246637 53726 675773
rect 59540 673650 59596 673659
rect 59540 673585 59596 673594
rect 59554 671101 59582 673585
rect 59542 671095 59594 671101
rect 59542 671037 59594 671043
rect 59540 659294 59596 659303
rect 59540 659229 59596 659238
rect 59554 656745 59582 659229
rect 59542 656739 59594 656745
rect 59542 656681 59594 656687
rect 59252 644938 59308 644947
rect 59252 644873 59308 644882
rect 59266 644535 59294 644873
rect 59254 644529 59306 644535
rect 59254 644471 59306 644477
rect 56086 630765 56138 630771
rect 56086 630707 56138 630713
rect 53878 606863 53930 606869
rect 53878 606805 53930 606811
rect 53780 589438 53836 589447
rect 53780 589373 53836 589382
rect 53794 252113 53822 589373
rect 53890 587481 53918 606805
rect 53878 587475 53930 587481
rect 53878 587417 53930 587423
rect 53878 515547 53930 515553
rect 53878 515489 53930 515495
rect 53890 437187 53918 515489
rect 53974 443619 54026 443625
rect 53974 443561 54026 443567
rect 53878 437181 53930 437187
rect 53878 437123 53930 437129
rect 53878 418459 53930 418465
rect 53878 418401 53930 418407
rect 53890 269281 53918 418401
rect 53986 349127 54014 443561
rect 53974 349121 54026 349127
rect 53974 349063 54026 349069
rect 53878 269275 53930 269281
rect 53878 269217 53930 269223
rect 53782 252107 53834 252113
rect 53782 252049 53834 252055
rect 56098 246859 56126 630707
rect 59540 630582 59596 630591
rect 59540 630517 59596 630526
rect 59554 627885 59582 630517
rect 59542 627879 59594 627885
rect 59542 627821 59594 627827
rect 59540 616226 59596 616235
rect 59540 616161 59596 616170
rect 59554 613529 59582 616161
rect 59542 613523 59594 613529
rect 59542 613465 59594 613471
rect 59542 601905 59594 601911
rect 59540 601870 59542 601879
rect 59594 601870 59596 601879
rect 59540 601805 59596 601814
rect 58196 587514 58252 587523
rect 58196 587449 58198 587458
rect 58250 587449 58252 587458
rect 58198 587417 58250 587423
rect 59540 573010 59596 573019
rect 59540 572945 59596 572954
rect 59554 570313 59582 572945
rect 59542 570307 59594 570313
rect 59542 570249 59594 570255
rect 59446 561575 59498 561581
rect 59446 561517 59498 561523
rect 59458 558959 59486 561517
rect 59444 558950 59500 558959
rect 59444 558885 59500 558894
rect 59542 544703 59594 544709
rect 59542 544645 59594 544651
rect 59554 544455 59582 544645
rect 59540 544446 59596 544455
rect 59540 544381 59596 544390
rect 59540 530090 59596 530099
rect 59540 530025 59596 530034
rect 59554 529983 59582 530025
rect 59542 529977 59594 529983
rect 59542 529919 59594 529925
rect 59540 515734 59596 515743
rect 59540 515669 59596 515678
rect 59554 515553 59582 515669
rect 59542 515547 59594 515553
rect 59542 515489 59594 515495
rect 59540 501230 59596 501239
rect 59540 501165 59542 501174
rect 59594 501165 59596 501174
rect 59542 501133 59594 501139
rect 58580 486874 58636 486883
rect 58580 486809 58636 486818
rect 58594 486767 58622 486809
rect 58582 486761 58634 486767
rect 58582 486703 58634 486709
rect 59540 472518 59596 472527
rect 59540 472453 59596 472462
rect 59554 472411 59582 472453
rect 59542 472405 59594 472411
rect 59542 472347 59594 472353
rect 59540 458162 59596 458171
rect 59540 458097 59596 458106
rect 59554 457981 59582 458097
rect 59542 457975 59594 457981
rect 59542 457917 59594 457923
rect 59540 443806 59596 443815
rect 59540 443741 59596 443750
rect 59554 443625 59582 443741
rect 59542 443619 59594 443625
rect 59542 443561 59594 443567
rect 59540 429450 59596 429459
rect 59540 429385 59596 429394
rect 59554 429195 59582 429385
rect 59542 429189 59594 429195
rect 59542 429131 59594 429137
rect 58388 415094 58444 415103
rect 58388 415029 58444 415038
rect 58402 414765 58430 415029
rect 58390 414759 58442 414765
rect 58390 414701 58442 414707
rect 57620 400738 57676 400747
rect 57620 400673 57676 400682
rect 57634 400409 57662 400673
rect 56278 400403 56330 400409
rect 56278 400345 56330 400351
rect 57622 400403 57674 400409
rect 57622 400345 57674 400351
rect 56182 357409 56234 357415
rect 56182 357351 56234 357357
rect 56194 262325 56222 357351
rect 56290 305541 56318 400345
rect 59252 386382 59308 386391
rect 59252 386317 59308 386326
rect 59266 385979 59294 386317
rect 59254 385973 59306 385979
rect 59254 385915 59306 385921
rect 59540 371878 59596 371887
rect 59540 371813 59596 371822
rect 59554 371623 59582 371813
rect 59542 371617 59594 371623
rect 59542 371559 59594 371565
rect 60212 357670 60268 357679
rect 60212 357605 60268 357614
rect 60226 357415 60254 357605
rect 60214 357409 60266 357415
rect 60214 357351 60266 357357
rect 58388 343166 58444 343175
rect 58388 343101 58444 343110
rect 58402 342837 58430 343101
rect 58390 342831 58442 342837
rect 58390 342773 58442 342779
rect 57812 328810 57868 328819
rect 57812 328745 57868 328754
rect 57826 328407 57854 328745
rect 57814 328401 57866 328407
rect 57814 328343 57866 328349
rect 58004 314602 58060 314611
rect 58004 314537 58060 314546
rect 58018 313977 58046 314537
rect 58006 313971 58058 313977
rect 58006 313913 58058 313919
rect 56278 305535 56330 305541
rect 56278 305477 56330 305483
rect 59444 300098 59500 300107
rect 59444 300033 59500 300042
rect 59458 299621 59486 300033
rect 59446 299615 59498 299621
rect 59446 299557 59498 299563
rect 56278 288071 56330 288077
rect 56278 288013 56330 288019
rect 56182 262319 56234 262325
rect 56182 262261 56234 262267
rect 56086 246853 56138 246859
rect 56086 246795 56138 246801
rect 56290 246711 56318 288013
rect 58100 285890 58156 285899
rect 58100 285825 58156 285834
rect 58114 285191 58142 285825
rect 58102 285185 58154 285191
rect 58102 285127 58154 285133
rect 60406 255141 60458 255147
rect 60406 255083 60458 255089
rect 56278 246705 56330 246711
rect 56278 246647 56330 246653
rect 53686 246631 53738 246637
rect 53686 246573 53738 246579
rect 53302 246557 53354 246563
rect 53302 246499 53354 246505
rect 53206 246483 53258 246489
rect 53206 246425 53258 246431
rect 60418 246267 60446 255083
rect 63298 246933 63326 986425
rect 65206 986409 65258 986415
rect 65206 986351 65258 986357
rect 65110 985003 65162 985009
rect 65110 984945 65162 984951
rect 64822 984189 64874 984195
rect 64822 984131 64874 984137
rect 64834 277939 64862 984131
rect 64918 983597 64970 983603
rect 64918 983539 64970 983545
rect 64930 278605 64958 983539
rect 65014 983523 65066 983529
rect 65014 983465 65066 983471
rect 64918 278599 64970 278605
rect 64918 278541 64970 278547
rect 64822 277933 64874 277939
rect 64822 277875 64874 277881
rect 65026 267875 65054 983465
rect 65014 267869 65066 267875
rect 65014 267811 65066 267817
rect 63286 246927 63338 246933
rect 63286 246869 63338 246875
rect 65122 246531 65150 984945
rect 65108 246522 65164 246531
rect 65108 246457 65164 246466
rect 60406 246261 60458 246267
rect 60406 246203 60458 246209
rect 65218 245939 65246 986351
rect 69058 984195 69086 987960
rect 69046 984189 69098 984195
rect 69046 984131 69098 984137
rect 73474 983534 73502 989237
rect 89602 983534 89630 990495
rect 92962 989301 92990 1005221
rect 93730 990559 93758 1005517
rect 93922 995887 93950 1010919
rect 97090 1005507 97118 1010919
rect 440662 1005723 440714 1005729
rect 440662 1005665 440714 1005671
rect 446614 1005723 446666 1005729
rect 446614 1005665 446666 1005671
rect 115702 1005649 115754 1005655
rect 115700 1005614 115702 1005623
rect 115754 1005614 115756 1005623
rect 115700 1005549 115756 1005558
rect 439222 1005575 439274 1005581
rect 439222 1005517 439274 1005523
rect 97078 1005501 97130 1005507
rect 118198 1005501 118250 1005507
rect 97078 1005443 97130 1005449
rect 102164 1005466 102220 1005475
rect 118198 1005443 118250 1005449
rect 298486 1005501 298538 1005507
rect 312790 1005501 312842 1005507
rect 298486 1005443 298538 1005449
rect 312788 1005466 312790 1005475
rect 365110 1005501 365162 1005507
rect 312842 1005466 312844 1005475
rect 102164 1005401 102166 1005410
rect 102218 1005401 102220 1005410
rect 102166 1005369 102218 1005375
rect 101494 1005353 101546 1005359
rect 101492 1005318 101494 1005327
rect 101546 1005318 101548 1005327
rect 101492 1005253 101548 1005262
rect 114164 1005318 114220 1005327
rect 114164 1005253 114166 1005262
rect 114218 1005253 114220 1005262
rect 114166 1005221 114218 1005227
rect 105430 1005205 105482 1005211
rect 105428 1005170 105430 1005179
rect 105482 1005170 105484 1005179
rect 105428 1005105 105484 1005114
rect 108886 1003725 108938 1003731
rect 108884 1003690 108886 1003699
rect 108938 1003690 108940 1003699
rect 108884 1003625 108940 1003634
rect 102836 1002506 102892 1002515
rect 97846 1002467 97898 1002473
rect 102836 1002441 102838 1002450
rect 97846 1002409 97898 1002415
rect 102890 1002441 102892 1002450
rect 102838 1002409 102890 1002415
rect 97750 1002319 97802 1002325
rect 97750 1002261 97802 1002267
rect 97762 999513 97790 1002261
rect 97750 999507 97802 999513
rect 97750 999449 97802 999455
rect 97858 995887 97886 1002409
rect 99766 1002393 99818 1002399
rect 103798 1002393 103850 1002399
rect 99766 1002335 99818 1002341
rect 100532 1002358 100588 1002367
rect 93910 995881 93962 995887
rect 93910 995823 93962 995829
rect 97846 995881 97898 995887
rect 97846 995823 97898 995829
rect 94964 995698 95020 995707
rect 94964 995633 95020 995642
rect 93718 990553 93770 990559
rect 93718 990495 93770 990501
rect 92950 989295 93002 989301
rect 92950 989237 93002 989243
rect 94978 985009 95006 995633
rect 99778 995263 99806 1002335
rect 103796 1002358 103798 1002367
rect 103850 1002358 103852 1002367
rect 100532 1002293 100534 1002302
rect 100586 1002293 100588 1002302
rect 100726 1002319 100778 1002325
rect 100534 1002261 100586 1002267
rect 103796 1002293 103852 1002302
rect 104468 1002358 104524 1002367
rect 104468 1002293 104470 1002302
rect 100726 1002261 100778 1002267
rect 104522 1002293 104524 1002302
rect 104470 1002261 104522 1002267
rect 99764 995254 99820 995263
rect 99764 995189 99820 995198
rect 100738 993815 100766 1002261
rect 115318 996103 115370 996109
rect 115318 996045 115370 996051
rect 106964 995994 107020 996003
rect 106498 995952 106964 995980
rect 106102 995807 106154 995813
rect 106102 995749 106154 995755
rect 100726 993809 100778 993815
rect 100726 993751 100778 993757
rect 94966 985003 95018 985009
rect 94966 984945 95018 984951
rect 106114 983548 106142 995749
rect 106498 993783 106526 995952
rect 106964 995929 107020 995938
rect 113300 995994 113356 996003
rect 113300 995929 113356 995938
rect 113314 995813 113342 995929
rect 115222 995881 115274 995887
rect 113396 995846 113452 995855
rect 113302 995807 113354 995813
rect 115222 995823 115274 995829
rect 113396 995781 113398 995790
rect 113302 995749 113354 995755
rect 113450 995781 113452 995790
rect 113398 995749 113450 995755
rect 115234 995559 115262 995823
rect 115220 995550 115276 995559
rect 115220 995485 115276 995494
rect 108212 995402 108268 995411
rect 108212 995337 108268 995346
rect 106484 993774 106540 993783
rect 106484 993709 106540 993718
rect 108226 993667 108254 995337
rect 109844 995254 109900 995263
rect 109844 995189 109900 995198
rect 109858 993741 109886 995189
rect 109846 993735 109898 993741
rect 109846 993677 109898 993683
rect 108214 993661 108266 993667
rect 108214 993603 108266 993609
rect 115234 986637 115262 995485
rect 115330 995411 115358 996045
rect 118102 995807 118154 995813
rect 118102 995749 118154 995755
rect 115316 995402 115372 995411
rect 115316 995337 115372 995346
rect 115330 986711 115358 995337
rect 115318 986705 115370 986711
rect 115318 986647 115370 986653
rect 115222 986631 115274 986637
rect 115222 986573 115274 986579
rect 118114 986563 118142 995749
rect 118210 995073 118238 1005443
rect 298390 1005427 298442 1005433
rect 298390 1005369 298442 1005375
rect 195478 1005205 195530 1005211
rect 209014 1005205 209066 1005211
rect 195478 1005147 195530 1005153
rect 209012 1005170 209014 1005179
rect 209066 1005170 209068 1005179
rect 143734 1002541 143786 1002547
rect 157942 1002541 157994 1002547
rect 143734 1002483 143786 1002489
rect 151220 1002506 151276 1002515
rect 143746 999532 143774 1002483
rect 144022 1002467 144074 1002473
rect 151220 1002441 151222 1002450
rect 144022 1002409 144074 1002415
rect 151274 1002441 151276 1002450
rect 157940 1002506 157942 1002515
rect 157994 1002506 157996 1002515
rect 157940 1002441 157996 1002450
rect 151222 1002409 151274 1002415
rect 143926 1002393 143978 1002399
rect 143926 1002335 143978 1002341
rect 143830 1000839 143882 1000845
rect 143830 1000781 143882 1000787
rect 143650 999504 143774 999532
rect 126646 999433 126698 999439
rect 126646 999375 126698 999381
rect 118198 995067 118250 995073
rect 118198 995009 118250 995015
rect 126658 993593 126686 999375
rect 127510 996103 127562 996109
rect 127510 996045 127562 996051
rect 127414 996029 127466 996035
rect 127414 995971 127466 995977
rect 127426 995887 127454 995971
rect 127522 995887 127550 996045
rect 127414 995881 127466 995887
rect 127414 995823 127466 995829
rect 127510 995881 127562 995887
rect 136724 995846 136780 995855
rect 127510 995823 127562 995829
rect 136464 995804 136724 995832
rect 137972 995846 138028 995855
rect 136724 995781 136780 995790
rect 137590 995807 137642 995813
rect 137760 995804 137972 995832
rect 142656 995813 143006 995832
rect 142656 995807 143018 995813
rect 142656 995804 142966 995807
rect 137972 995781 138028 995790
rect 137590 995749 137642 995755
rect 142966 995749 143018 995755
rect 133654 995733 133706 995739
rect 133440 995681 133654 995684
rect 137602 995707 137630 995749
rect 141046 995733 141098 995739
rect 133440 995675 133706 995681
rect 137588 995698 137644 995707
rect 133440 995656 133694 995675
rect 139220 995698 139276 995707
rect 138960 995656 139220 995684
rect 137588 995633 137644 995642
rect 140784 995681 141046 995684
rect 140784 995675 141098 995681
rect 140784 995656 141086 995675
rect 139220 995633 139276 995642
rect 132406 995585 132458 995591
rect 128482 993667 128510 995522
rect 129120 995508 129374 995536
rect 129346 993815 129374 995508
rect 129730 993931 129758 995522
rect 131616 995508 131870 995536
rect 132144 995533 132406 995536
rect 137396 995550 137452 995559
rect 132144 995527 132458 995533
rect 132144 995508 132446 995527
rect 132816 995508 133118 995536
rect 131842 994185 131870 995508
rect 133090 995443 133118 995508
rect 133078 995437 133130 995443
rect 133078 995379 133130 995385
rect 134002 995295 134030 995522
rect 133990 995289 134042 995295
rect 133990 995231 134042 995237
rect 131830 994179 131882 994185
rect 131830 994121 131882 994127
rect 129716 993922 129772 993931
rect 129716 993857 129772 993866
rect 129334 993809 129386 993815
rect 129334 993751 129386 993757
rect 128470 993661 128522 993667
rect 128470 993603 128522 993609
rect 134626 993593 134654 995522
rect 135936 995508 136286 995536
rect 137136 995508 137396 995536
rect 136258 995443 136286 995508
rect 140160 995508 140414 995536
rect 137396 995485 137452 995494
rect 136246 995437 136298 995443
rect 140386 995411 140414 995508
rect 143650 995443 143678 999504
rect 143734 999433 143786 999439
rect 143734 999375 143786 999381
rect 143746 995813 143774 999375
rect 143734 995807 143786 995813
rect 143734 995749 143786 995755
rect 143842 995739 143870 1000781
rect 143938 995855 143966 1002335
rect 144034 996003 144062 1002409
rect 150358 1002393 150410 1002399
rect 150356 1002358 150358 1002367
rect 150410 1002358 150412 1002367
rect 144118 1002319 144170 1002325
rect 150356 1002293 150412 1002302
rect 178486 1002319 178538 1002325
rect 144118 1002261 144170 1002267
rect 178486 1002261 178538 1002267
rect 144020 995994 144076 996003
rect 144020 995929 144076 995938
rect 144022 995881 144074 995887
rect 143924 995846 143980 995855
rect 144022 995823 144074 995829
rect 143924 995781 143980 995790
rect 143830 995733 143882 995739
rect 143830 995675 143882 995681
rect 144034 995591 144062 995823
rect 144022 995585 144074 995591
rect 144022 995527 144074 995533
rect 143638 995437 143690 995443
rect 141154 995411 141278 995425
rect 136246 995379 136298 995385
rect 140372 995402 140428 995411
rect 140372 995337 140428 995346
rect 141140 995402 141278 995411
rect 141196 995397 141278 995402
rect 141140 995337 141196 995346
rect 141250 995221 141278 995397
rect 144130 995388 144158 1002261
rect 160244 1000878 160300 1000887
rect 160244 1000813 160246 1000822
rect 160298 1000813 160300 1000822
rect 160246 1000781 160298 1000787
rect 156886 999433 156938 999439
rect 156884 999398 156886 999407
rect 156938 999398 156940 999407
rect 156884 999333 156940 999342
rect 163126 996177 163178 996183
rect 162260 996142 162316 996151
rect 162260 996077 162262 996086
rect 162314 996077 162316 996086
rect 163124 996142 163126 996151
rect 163178 996142 163180 996151
rect 163124 996077 163180 996086
rect 164084 996142 164140 996151
rect 164084 996077 164140 996086
rect 162262 996045 162314 996051
rect 164098 996035 164126 996077
rect 164086 996029 164138 996035
rect 145268 995994 145324 996003
rect 145268 995929 145324 995938
rect 149108 995994 149164 996003
rect 149492 995994 149548 996003
rect 149164 995952 149492 995980
rect 149108 995929 149164 995938
rect 149492 995929 149548 995938
rect 151988 995994 152044 996003
rect 151988 995929 151990 995938
rect 143638 995379 143690 995385
rect 143938 995360 144158 995388
rect 143938 995295 143966 995360
rect 143926 995289 143978 995295
rect 143926 995231 143978 995237
rect 141238 995215 141290 995221
rect 141238 995157 141290 995163
rect 126646 993587 126698 993593
rect 126646 993529 126698 993535
rect 134614 993587 134666 993593
rect 134614 993529 134666 993535
rect 138262 989295 138314 989301
rect 138262 989237 138314 989243
rect 122038 988333 122090 988339
rect 122038 988275 122090 988281
rect 118102 986557 118154 986563
rect 118102 986499 118154 986505
rect 105840 983520 106142 983548
rect 122050 983534 122078 988275
rect 138274 983534 138302 989237
rect 145282 986489 145310 995929
rect 152042 995929 152044 995938
rect 152852 995994 152908 996003
rect 152852 995929 152908 995938
rect 155348 995994 155404 996003
rect 164182 996029 164234 996035
rect 164086 995971 164138 995977
rect 164180 995994 164182 996003
rect 164234 995994 164236 996003
rect 155348 995929 155404 995938
rect 164180 995929 164236 995938
rect 151990 995897 152042 995903
rect 146806 995807 146858 995813
rect 146806 995749 146858 995755
rect 146818 995369 146846 995749
rect 151702 995733 151754 995739
rect 151702 995675 151754 995681
rect 146806 995363 146858 995369
rect 146806 995305 146858 995311
rect 151714 993815 151742 995675
rect 152866 995559 152894 995929
rect 155362 995887 155390 995929
rect 155350 995881 155402 995887
rect 154292 995846 154348 995855
rect 155350 995823 155402 995829
rect 156308 995846 156364 995855
rect 154292 995781 154294 995790
rect 154346 995781 154348 995790
rect 165620 995846 165676 995855
rect 156308 995781 156364 995790
rect 164086 995807 164138 995813
rect 154294 995749 154346 995755
rect 156322 995739 156350 995781
rect 165620 995781 165622 995790
rect 164086 995749 164138 995755
rect 165674 995781 165676 995790
rect 166196 995846 166252 995855
rect 166196 995781 166252 995790
rect 165622 995749 165674 995755
rect 156310 995733 156362 995739
rect 163990 995733 164042 995739
rect 156310 995675 156362 995681
rect 159572 995698 159628 995707
rect 163990 995675 164042 995681
rect 159572 995633 159628 995642
rect 152852 995550 152908 995559
rect 152852 995485 152908 995494
rect 158804 995550 158860 995559
rect 158804 995485 158860 995494
rect 158996 995550 159052 995559
rect 158996 995485 159052 995494
rect 158818 994185 158846 995485
rect 158806 994179 158858 994185
rect 158806 994121 158858 994127
rect 159010 993931 159038 995485
rect 158996 993922 159052 993931
rect 158996 993857 159052 993866
rect 151702 993809 151754 993815
rect 151702 993751 151754 993757
rect 159586 993667 159614 995633
rect 161204 995254 161260 995263
rect 161204 995189 161206 995198
rect 161258 995189 161260 995198
rect 161206 995157 161258 995163
rect 159574 993661 159626 993667
rect 159574 993603 159626 993609
rect 164002 989375 164030 995675
rect 154486 989369 154538 989375
rect 154486 989311 154538 989317
rect 163990 989369 164042 989375
rect 163990 989311 164042 989317
rect 145270 986483 145322 986489
rect 145270 986425 145322 986431
rect 154498 983534 154526 989311
rect 164098 989301 164126 995749
rect 166210 995739 166238 995781
rect 166198 995733 166250 995739
rect 178498 995707 178526 1002261
rect 195286 1001061 195338 1001067
rect 195286 1001003 195338 1001009
rect 195190 996547 195242 996553
rect 195190 996489 195242 996495
rect 195202 995855 195230 996489
rect 185108 995846 185164 995855
rect 184848 995804 185108 995832
rect 188756 995846 188812 995855
rect 187344 995813 187742 995832
rect 187344 995807 187754 995813
rect 187344 995804 187702 995807
rect 185108 995781 185164 995790
rect 188544 995804 188756 995832
rect 195188 995846 195244 995855
rect 190368 995813 190622 995832
rect 190368 995807 190634 995813
rect 190368 995804 190582 995807
rect 188756 995781 188812 995790
rect 187702 995749 187754 995755
rect 195188 995781 195244 995790
rect 190582 995749 190634 995755
rect 188086 995733 188138 995739
rect 166198 995675 166250 995681
rect 170324 995698 170380 995707
rect 170324 995633 170380 995642
rect 178484 995698 178540 995707
rect 178484 995633 178540 995642
rect 185204 995698 185260 995707
rect 185260 995670 185424 995684
rect 187872 995681 188086 995684
rect 195092 995698 195148 995707
rect 187872 995675 188138 995681
rect 185260 995656 185438 995670
rect 187872 995656 188126 995675
rect 194064 995665 194462 995684
rect 194064 995659 194474 995665
rect 194064 995656 194422 995659
rect 185204 995633 185260 995642
rect 166964 995254 167020 995263
rect 167020 995212 167198 995240
rect 166964 995189 167020 995198
rect 167170 995115 167198 995212
rect 167156 995106 167212 995115
rect 167156 995041 167212 995050
rect 164086 989295 164138 989301
rect 164086 989237 164138 989243
rect 170338 983548 170366 995633
rect 184340 995550 184396 995559
rect 179842 993667 179870 995522
rect 180514 993815 180542 995522
rect 181152 995508 181406 995536
rect 180502 993809 180554 993815
rect 180502 993751 180554 993757
rect 181378 993741 181406 995508
rect 181462 995215 181514 995221
rect 181462 995157 181514 995163
rect 181474 995115 181502 995157
rect 181460 995106 181516 995115
rect 181460 995041 181516 995050
rect 183010 994227 183038 995522
rect 183552 995508 183806 995536
rect 184176 995508 184340 995536
rect 183778 995263 183806 995508
rect 184340 995485 184396 995494
rect 183764 995254 183820 995263
rect 183764 995189 183820 995198
rect 182996 994218 183052 994227
rect 182996 994153 183052 994162
rect 185410 994079 185438 995656
rect 195298 995665 195326 1001003
rect 195382 1000839 195434 1000845
rect 195382 1000781 195434 1000787
rect 195092 995633 195148 995642
rect 195286 995659 195338 995665
rect 194422 995601 194474 995607
rect 192502 995585 192554 995591
rect 189428 995550 189484 995559
rect 186048 995508 186206 995536
rect 189168 995508 189428 995536
rect 185396 994070 185452 994079
rect 185396 994005 185452 994014
rect 181366 993735 181418 993741
rect 181366 993677 181418 993683
rect 179830 993661 179882 993667
rect 179830 993603 179882 993609
rect 186178 993593 186206 995508
rect 192192 995533 192502 995536
rect 192192 995527 192554 995533
rect 189428 995485 189484 995494
rect 191554 993931 191582 995522
rect 192192 995508 192542 995527
rect 191540 993922 191596 993931
rect 191540 993857 191596 993866
rect 186166 993587 186218 993593
rect 186166 993529 186218 993535
rect 186934 988259 186986 988265
rect 186934 988201 186986 988207
rect 170338 983520 170736 983548
rect 186946 983534 186974 988201
rect 195106 986415 195134 995633
rect 195286 995601 195338 995607
rect 195394 995591 195422 1000781
rect 195490 995887 195518 1005147
rect 209012 1005105 209068 1005114
rect 208342 1001061 208394 1001067
rect 208340 1001026 208342 1001035
rect 208394 1001026 208396 1001035
rect 208340 1000961 208396 1000970
rect 211700 1000878 211756 1000887
rect 211700 1000813 211702 1000822
rect 211754 1000813 211756 1000822
rect 211702 1000781 211754 1000787
rect 298102 1000025 298154 1000031
rect 298102 999967 298154 999973
rect 256436 999546 256492 999555
rect 246934 999507 246986 999513
rect 298114 999532 298142 999967
rect 298294 999729 298346 999735
rect 298294 999671 298346 999677
rect 256436 999481 256438 999490
rect 246934 999449 246986 999455
rect 256490 999481 256492 999490
rect 298018 999504 298142 999532
rect 298198 999507 298250 999513
rect 256438 999449 256490 999455
rect 195766 999433 195818 999439
rect 195766 999375 195818 999381
rect 224662 999433 224714 999439
rect 224662 999375 224714 999381
rect 246550 999433 246602 999439
rect 246550 999375 246602 999381
rect 195478 995881 195530 995887
rect 195478 995823 195530 995829
rect 195382 995585 195434 995591
rect 195382 995527 195434 995533
rect 195778 993593 195806 999375
rect 204212 996586 204268 996595
rect 204212 996521 204214 996530
rect 204266 996521 204268 996530
rect 204214 996489 204266 996495
rect 214102 996177 214154 996183
rect 213332 996142 213388 996151
rect 213332 996077 213334 996086
rect 213386 996077 213388 996086
rect 214100 996142 214102 996151
rect 214154 996142 214156 996151
rect 214100 996077 214156 996086
rect 215636 996142 215692 996151
rect 215636 996077 215638 996086
rect 213334 996045 213386 996051
rect 215690 996077 215692 996086
rect 215638 996045 215690 996051
rect 198644 995994 198700 996003
rect 198644 995929 198646 995938
rect 198698 995929 198700 995938
rect 203444 995994 203500 996003
rect 203444 995929 203446 995938
rect 198646 995897 198698 995903
rect 203498 995929 203500 995938
rect 205652 995994 205708 996003
rect 205652 995929 205708 995938
rect 206516 995994 206572 996003
rect 206516 995929 206572 995938
rect 213046 995955 213098 995961
rect 203446 995897 203498 995903
rect 201716 995846 201772 995855
rect 201716 995781 201772 995790
rect 202868 995846 202924 995855
rect 202868 995781 202924 995790
rect 204980 995846 205036 995855
rect 204980 995781 204982 995790
rect 201622 995659 201674 995665
rect 201622 995601 201674 995607
rect 201526 995215 201578 995221
rect 201526 995157 201578 995163
rect 201538 995115 201566 995157
rect 201524 995106 201580 995115
rect 201524 995041 201580 995050
rect 201634 993815 201662 995601
rect 201730 995559 201758 995781
rect 202882 995739 202910 995781
rect 205034 995781 205036 995790
rect 204982 995749 205034 995755
rect 202870 995733 202922 995739
rect 202870 995675 202922 995681
rect 201716 995550 201772 995559
rect 201716 995485 201772 995494
rect 205666 995411 205694 995929
rect 205652 995402 205708 995411
rect 205652 995337 205708 995346
rect 206530 995295 206558 995929
rect 213046 995897 213098 995903
rect 206996 995698 207052 995707
rect 206996 995633 206998 995642
rect 207050 995633 207052 995642
rect 206998 995601 207050 995607
rect 210260 995402 210316 995411
rect 210260 995337 210316 995346
rect 211028 995402 211084 995411
rect 211028 995337 211084 995346
rect 212660 995402 212716 995411
rect 212660 995337 212716 995346
rect 201718 995289 201770 995295
rect 201716 995254 201718 995263
rect 206518 995289 206570 995295
rect 201770 995254 201772 995263
rect 206518 995231 206570 995237
rect 201716 995189 201772 995198
rect 210274 994227 210302 995337
rect 210260 994218 210316 994227
rect 210260 994153 210316 994162
rect 201622 993809 201674 993815
rect 201622 993751 201674 993757
rect 211042 993667 211070 995337
rect 212674 993741 212702 995337
rect 212662 993735 212714 993741
rect 212662 993677 212714 993683
rect 211030 993661 211082 993667
rect 211030 993603 211082 993609
rect 195766 993587 195818 993593
rect 195766 993529 195818 993535
rect 213058 988857 213086 995897
rect 213346 995887 213374 996045
rect 215446 996029 215498 996035
rect 215444 995994 215446 996003
rect 215498 995994 215500 996003
rect 215444 995929 215500 995938
rect 217076 995994 217132 996003
rect 217076 995929 217078 995938
rect 217130 995929 217132 995938
rect 221780 995994 221836 996003
rect 221780 995929 221836 995938
rect 217078 995897 217130 995903
rect 213334 995881 213386 995887
rect 213334 995823 213386 995829
rect 221794 990559 221822 995929
rect 224674 995813 224702 999375
rect 241844 995846 241900 995855
rect 236256 995813 236510 995832
rect 224662 995807 224714 995813
rect 236256 995807 236522 995813
rect 236256 995804 236470 995807
rect 224662 995749 224714 995755
rect 241776 995804 241844 995832
rect 243860 995846 243916 995855
rect 243600 995804 243860 995832
rect 241844 995781 241900 995790
rect 243860 995781 243916 995790
rect 236470 995749 236522 995755
rect 246562 995739 246590 999375
rect 246946 996003 246974 999449
rect 259510 999433 259562 999439
rect 259508 999398 259510 999407
rect 259562 999398 259564 999407
rect 259508 999333 259564 999342
rect 263060 996586 263116 996595
rect 251254 996547 251306 996553
rect 263060 996521 263062 996530
rect 251254 996489 251306 996495
rect 263114 996521 263116 996530
rect 263062 996489 263114 996495
rect 246932 995994 246988 996003
rect 246932 995929 246988 995938
rect 247508 995994 247564 996003
rect 247508 995929 247564 995938
rect 250486 995955 250538 995961
rect 245686 995733 245738 995739
rect 222932 995698 222988 995707
rect 240788 995698 240844 995707
rect 222932 995633 222988 995642
rect 237238 995659 237290 995665
rect 219478 990553 219530 990559
rect 219478 990495 219530 990501
rect 221782 990553 221834 990559
rect 221782 990495 221834 990501
rect 203158 988851 203210 988857
rect 203158 988793 203210 988799
rect 213046 988851 213098 988857
rect 213046 988793 213098 988799
rect 195094 986409 195146 986415
rect 195094 986351 195146 986357
rect 203170 983534 203198 988793
rect 219490 983534 219518 990495
rect 222946 989375 222974 995633
rect 240576 995656 240788 995684
rect 245424 995681 245686 995684
rect 245424 995675 245738 995681
rect 246550 995733 246602 995739
rect 246550 995675 246602 995681
rect 245424 995656 245726 995675
rect 240788 995633 240844 995642
rect 237238 995601 237290 995607
rect 237250 995536 237278 995601
rect 239540 995550 239596 995559
rect 231264 995508 231518 995536
rect 231936 995508 232190 995536
rect 227348 995106 227404 995115
rect 227540 995106 227596 995115
rect 227404 995064 227540 995092
rect 227348 995041 227404 995050
rect 227540 995041 227596 995050
rect 231490 993815 231518 995508
rect 232162 994375 232190 995508
rect 232148 994366 232204 994375
rect 232148 994301 232204 994310
rect 231478 993809 231530 993815
rect 231478 993751 231530 993757
rect 232546 993741 232574 995522
rect 234370 994227 234398 995522
rect 234356 994218 234412 994227
rect 234356 994153 234412 994162
rect 234946 993963 234974 995522
rect 235584 995508 235838 995536
rect 237250 995522 237456 995536
rect 235810 994523 235838 995508
rect 235796 994514 235852 994523
rect 235796 994449 235852 994458
rect 236770 994079 236798 995522
rect 237250 995508 237470 995522
rect 236756 994070 236812 994079
rect 236756 994005 236812 994014
rect 234934 993957 234986 993963
rect 234934 993899 234986 993905
rect 232534 993735 232586 993741
rect 232534 993677 232586 993683
rect 237442 993667 237470 995508
rect 238690 993889 238718 995522
rect 239280 995508 239540 995536
rect 239952 995508 240254 995536
rect 242976 995508 243230 995536
rect 239540 995485 239596 995494
rect 240226 995411 240254 995508
rect 240212 995402 240268 995411
rect 240212 995337 240268 995346
rect 242324 994662 242380 994671
rect 242324 994597 242380 994606
rect 242338 994375 242366 994597
rect 242324 994366 242380 994375
rect 242324 994301 242380 994310
rect 242516 994366 242572 994375
rect 242516 994301 242572 994310
rect 242530 994079 242558 994301
rect 243202 994079 243230 995508
rect 247412 995106 247468 995115
rect 247412 995041 247468 995050
rect 247426 994999 247454 995041
rect 247414 994993 247466 994999
rect 247414 994935 247466 994941
rect 244820 994366 244876 994375
rect 244820 994301 244876 994310
rect 244834 994111 244862 994301
rect 244822 994105 244874 994111
rect 242516 994070 242572 994079
rect 242516 994005 242572 994014
rect 243188 994070 243244 994079
rect 244822 994047 244874 994053
rect 243188 994005 243244 994014
rect 238678 993883 238730 993889
rect 238678 993825 238730 993831
rect 237430 993661 237482 993667
rect 237430 993603 237482 993609
rect 222934 989369 222986 989375
rect 222934 989311 222986 989317
rect 235606 989369 235658 989375
rect 235606 989311 235658 989317
rect 235618 983534 235646 989311
rect 247522 987821 247550 995929
rect 250486 995897 250538 995903
rect 250102 995881 250154 995887
rect 250102 995823 250154 995829
rect 247606 995733 247658 995739
rect 247606 995675 247658 995681
rect 247618 994523 247646 995675
rect 250114 995411 250142 995823
rect 250100 995402 250156 995411
rect 250100 995337 250156 995346
rect 250498 994671 250526 995897
rect 251266 995855 251294 996489
rect 265942 996177 265994 996183
rect 265940 996142 265942 996151
rect 270742 996177 270794 996183
rect 265994 996142 265996 996151
rect 265940 996077 265996 996086
rect 266996 996142 267052 996151
rect 270742 996119 270794 996125
rect 266996 996077 266998 996086
rect 267050 996077 267052 996086
rect 266998 996045 267050 996051
rect 264694 996029 264746 996035
rect 258836 995994 258892 996003
rect 258836 995929 258838 995938
rect 258890 995929 258892 995938
rect 264692 995994 264694 996003
rect 267766 996029 267818 996035
rect 264746 995994 264748 996003
rect 267862 996029 267914 996035
rect 267818 995977 267862 995980
rect 267766 995971 267914 995977
rect 267778 995952 267902 995971
rect 264692 995929 264748 995938
rect 258838 995897 258890 995903
rect 255574 995881 255626 995887
rect 251252 995846 251308 995855
rect 251252 995781 251308 995790
rect 254804 995846 254860 995855
rect 254804 995781 254806 995790
rect 254858 995781 254860 995790
rect 255572 995846 255574 995855
rect 255626 995846 255628 995855
rect 255572 995781 255628 995790
rect 257492 995846 257548 995855
rect 257492 995781 257548 995790
rect 258260 995846 258316 995855
rect 258260 995781 258316 995790
rect 260756 995846 260812 995855
rect 260756 995781 260812 995790
rect 268244 995846 268300 995855
rect 268244 995781 268246 995790
rect 254806 995749 254858 995755
rect 257506 995739 257534 995781
rect 257494 995733 257546 995739
rect 257494 995675 257546 995681
rect 258274 995665 258302 995781
rect 253078 995659 253130 995665
rect 253078 995601 253130 995607
rect 258262 995659 258314 995665
rect 258262 995601 258314 995607
rect 250484 994662 250540 994671
rect 250484 994597 250540 994606
rect 247604 994514 247660 994523
rect 247604 994449 247660 994458
rect 253090 993963 253118 995601
rect 254708 995402 254764 995411
rect 254708 995337 254764 995346
rect 254722 994227 254750 995337
rect 259124 995106 259180 995115
rect 259124 995041 259180 995050
rect 259138 994999 259166 995041
rect 259126 994993 259178 994999
rect 259126 994935 259178 994941
rect 254708 994218 254764 994227
rect 254708 994153 254764 994162
rect 253078 993957 253130 993963
rect 253078 993899 253130 993905
rect 260770 993889 260798 995781
rect 268298 995781 268300 995790
rect 268436 995846 268492 995855
rect 268436 995781 268492 995790
rect 268246 995749 268298 995755
rect 262388 995698 262444 995707
rect 262388 995633 262444 995642
rect 262196 995106 262252 995115
rect 262196 995041 262252 995050
rect 262210 994819 262238 995041
rect 262196 994810 262252 994819
rect 262196 994745 262252 994754
rect 260758 993883 260810 993889
rect 260758 993825 260810 993831
rect 262402 993815 262430 995633
rect 264020 995402 264076 995411
rect 264020 995337 264076 995346
rect 262390 993809 262442 993815
rect 262390 993751 262442 993757
rect 264034 993741 264062 995337
rect 264022 993735 264074 993741
rect 264022 993677 264074 993683
rect 251830 988185 251882 988191
rect 251830 988127 251882 988133
rect 244726 987815 244778 987821
rect 244726 987757 244778 987763
rect 247510 987815 247562 987821
rect 247510 987757 247562 987763
rect 244738 983603 244766 987757
rect 244726 983597 244778 983603
rect 244726 983539 244778 983545
rect 251842 983534 251870 988127
rect 268450 983548 268478 995781
rect 270754 995707 270782 996119
rect 273620 995846 273676 995855
rect 283124 995846 283180 995855
rect 273620 995781 273676 995790
rect 273718 995807 273770 995813
rect 270740 995698 270796 995707
rect 270740 995633 270796 995642
rect 273634 989375 273662 995781
rect 282864 995804 283124 995832
rect 294836 995846 294892 995855
rect 283536 995813 283838 995832
rect 290880 995813 291230 995832
rect 283536 995807 283850 995813
rect 283536 995804 283798 995807
rect 283124 995781 283180 995790
rect 273718 995749 273770 995755
rect 283798 995749 283850 995755
rect 289462 995807 289514 995813
rect 290880 995807 291242 995813
rect 290880 995804 291190 995807
rect 289462 995749 289514 995755
rect 294576 995804 294836 995832
rect 294836 995781 294892 995790
rect 291190 995749 291242 995755
rect 273622 989369 273674 989375
rect 273622 989311 273674 989317
rect 273730 989301 273758 995749
rect 286292 995698 286348 995707
rect 286032 995656 286292 995684
rect 286292 995633 286348 995642
rect 284160 995517 284414 995536
rect 284160 995511 284426 995517
rect 284160 995508 284374 995511
rect 286560 995508 286814 995536
rect 284374 995453 284426 995459
rect 286786 995443 286814 995508
rect 286774 995437 286826 995443
rect 286774 995379 286826 995385
rect 287170 995221 287198 995522
rect 287158 995215 287210 995221
rect 287158 995157 287210 995163
rect 287842 994999 287870 995522
rect 288130 995508 288384 995536
rect 289056 995508 289310 995536
rect 287830 994993 287882 994999
rect 287830 994935 287882 994941
rect 279286 994105 279338 994111
rect 279286 994047 279338 994053
rect 279298 993593 279326 994047
rect 288130 993593 288158 995508
rect 289282 994555 289310 995508
rect 289474 995221 289502 995749
rect 291766 995733 291818 995739
rect 291504 995681 291766 995684
rect 291504 995675 291818 995681
rect 291504 995656 291806 995675
rect 297072 995665 297374 995684
rect 297072 995659 297386 995665
rect 297072 995656 297334 995659
rect 297334 995601 297386 995607
rect 295414 995585 295466 995591
rect 292532 995550 292588 995559
rect 289462 995215 289514 995221
rect 289462 995157 289514 995163
rect 290338 994851 290366 995522
rect 292176 995508 292532 995536
rect 293376 995517 293726 995536
rect 295200 995533 295414 995536
rect 295200 995527 295466 995533
rect 293376 995511 293738 995517
rect 293376 995508 293686 995511
rect 292532 995485 292588 995494
rect 295200 995508 295454 995527
rect 298018 995517 298046 999504
rect 298198 999449 298250 999455
rect 298102 999433 298154 999439
rect 298102 999375 298154 999381
rect 298114 995665 298142 999375
rect 298102 995659 298154 995665
rect 298102 995601 298154 995607
rect 298210 995591 298238 999449
rect 298306 995855 298334 999671
rect 298402 996003 298430 1005369
rect 298388 995994 298444 996003
rect 298388 995929 298444 995938
rect 298292 995846 298348 995855
rect 298292 995781 298348 995790
rect 298498 995707 298526 1005443
rect 312788 1005401 312844 1005410
rect 313844 1005466 313900 1005475
rect 313844 1005401 313846 1005410
rect 313898 1005401 313900 1005410
rect 321044 1005466 321100 1005475
rect 321428 1005466 321484 1005475
rect 321100 1005424 321428 1005452
rect 321044 1005401 321100 1005410
rect 321428 1005401 321484 1005410
rect 325460 1005466 325516 1005475
rect 325460 1005401 325516 1005410
rect 365108 1005466 365110 1005475
rect 383638 1005501 383690 1005507
rect 365162 1005466 365164 1005475
rect 433174 1005501 433226 1005507
rect 383638 1005443 383690 1005449
rect 430868 1005466 430924 1005475
rect 365108 1005401 365164 1005410
rect 313846 1005369 313898 1005375
rect 298678 1005353 298730 1005359
rect 309622 1005353 309674 1005359
rect 298678 1005295 298730 1005301
rect 308756 1005318 308812 1005327
rect 298582 999581 298634 999587
rect 298582 999523 298634 999529
rect 298484 995698 298540 995707
rect 298484 995633 298540 995642
rect 298198 995585 298250 995591
rect 298198 995527 298250 995533
rect 298006 995511 298058 995517
rect 293686 995453 293738 995459
rect 298006 995453 298058 995459
rect 298594 995443 298622 999523
rect 298582 995437 298634 995443
rect 298582 995379 298634 995385
rect 298690 995221 298718 1005295
rect 298774 1005279 298826 1005285
rect 308756 1005253 308758 1005262
rect 298774 1005221 298826 1005227
rect 308810 1005253 308812 1005262
rect 309620 1005318 309622 1005327
rect 309674 1005318 309676 1005327
rect 309620 1005253 309676 1005262
rect 318644 1005318 318700 1005327
rect 318644 1005253 318646 1005262
rect 308758 1005221 308810 1005227
rect 318698 1005253 318700 1005262
rect 318646 1005221 318698 1005227
rect 298786 995887 298814 1005221
rect 325474 1005211 325502 1005401
rect 358678 1005353 358730 1005359
rect 358676 1005318 358678 1005327
rect 366262 1005353 366314 1005359
rect 358730 1005318 358732 1005327
rect 328726 1005279 328778 1005285
rect 358676 1005253 358732 1005262
rect 359924 1005318 359980 1005327
rect 366262 1005295 366314 1005301
rect 359924 1005253 359926 1005262
rect 328726 1005221 328778 1005227
rect 359978 1005253 359980 1005262
rect 359926 1005221 359978 1005227
rect 299542 1005205 299594 1005211
rect 310294 1005205 310346 1005211
rect 299542 1005147 299594 1005153
rect 310292 1005170 310294 1005179
rect 325462 1005205 325514 1005211
rect 310346 1005170 310348 1005179
rect 299554 996572 299582 1005147
rect 325462 1005147 325514 1005153
rect 310292 1005105 310348 1005114
rect 308084 1002654 308140 1002663
rect 308084 1002589 308140 1002598
rect 308098 1000031 308126 1002589
rect 308086 1000025 308138 1000031
rect 308086 999967 308138 999973
rect 315478 999581 315530 999587
rect 314708 999546 314764 999555
rect 314708 999481 314710 999490
rect 314762 999481 314764 999490
rect 315476 999546 315478 999555
rect 315530 999546 315532 999555
rect 315476 999481 315532 999490
rect 314710 999449 314762 999455
rect 311446 999433 311498 999439
rect 311444 999398 311446 999407
rect 311498 999398 311500 999407
rect 311444 999333 311500 999342
rect 320950 997953 321002 997959
rect 320950 997895 321002 997901
rect 302422 997805 302474 997811
rect 302422 997747 302474 997753
rect 299458 996544 299582 996572
rect 299458 995961 299486 996544
rect 299446 995955 299498 995961
rect 299446 995897 299498 995903
rect 298774 995881 298826 995887
rect 298774 995823 298826 995829
rect 299156 995698 299212 995707
rect 299156 995633 299212 995642
rect 298678 995215 298730 995221
rect 298678 995157 298730 995163
rect 290326 994845 290378 994851
rect 290326 994787 290378 994793
rect 289270 994549 289322 994555
rect 289270 994491 289322 994497
rect 296662 994549 296714 994555
rect 296662 994491 296714 994497
rect 289282 993667 289310 994491
rect 296674 994227 296702 994491
rect 296660 994218 296716 994227
rect 296660 994153 296716 994162
rect 289270 993661 289322 993667
rect 289270 993603 289322 993609
rect 279286 993587 279338 993593
rect 279286 993529 279338 993535
rect 288118 993587 288170 993593
rect 288118 993529 288170 993535
rect 284278 989369 284330 989375
rect 284278 989311 284330 989317
rect 273718 989295 273770 989301
rect 273718 989237 273770 989243
rect 277942 985151 277994 985157
rect 277942 985093 277994 985099
rect 268176 983520 268478 983548
rect 277954 983529 277982 985093
rect 284290 983534 284318 989311
rect 299170 988709 299198 995633
rect 302434 995147 302462 997747
rect 319798 996473 319850 996479
rect 319798 996415 319850 996421
rect 318646 996177 318698 996183
rect 317108 996142 317164 996151
rect 317108 996077 317110 996086
rect 317162 996077 317164 996086
rect 318644 996142 318646 996151
rect 318698 996142 318700 996151
rect 318644 996077 318700 996086
rect 317110 996045 317162 996051
rect 316342 996029 316394 996035
rect 305588 995994 305644 996003
rect 305588 995929 305644 995938
rect 316340 995994 316342 996003
rect 319702 996029 319754 996035
rect 316394 995994 316396 996003
rect 319810 995980 319838 996415
rect 320962 996109 320990 997895
rect 328738 997737 328766 1005221
rect 331222 1005205 331274 1005211
rect 357046 1005205 357098 1005211
rect 331222 1005147 331274 1005153
rect 357044 1005170 357046 1005179
rect 357098 1005170 357100 1005179
rect 328726 997731 328778 997737
rect 328726 997673 328778 997679
rect 320950 996103 321002 996109
rect 320950 996045 321002 996051
rect 319754 995977 319838 995980
rect 319702 995971 319838 995977
rect 319714 995952 319838 995971
rect 328244 995994 328300 996003
rect 316340 995929 316396 995938
rect 328244 995929 328300 995938
rect 305602 995813 305630 995929
rect 306452 995846 306508 995855
rect 305590 995807 305642 995813
rect 306452 995781 306508 995790
rect 307412 995846 307468 995855
rect 307412 995781 307468 995790
rect 311924 995846 311980 995855
rect 311924 995781 311980 995790
rect 305590 995749 305642 995755
rect 302422 995141 302474 995147
rect 302422 995083 302474 995089
rect 306466 994999 306494 995781
rect 307426 995739 307454 995781
rect 307414 995733 307466 995739
rect 307414 995675 307466 995681
rect 306454 994993 306506 994999
rect 306454 994935 306506 994941
rect 311938 994851 311966 995781
rect 325268 995698 325324 995707
rect 325268 995633 325324 995642
rect 316724 995254 316780 995263
rect 316724 995189 316780 995198
rect 316738 995115 316766 995189
rect 316724 995106 316780 995115
rect 316724 995041 316780 995050
rect 311926 994845 311978 994851
rect 311926 994787 311978 994793
rect 325282 989301 325310 995633
rect 328258 989375 328286 995929
rect 331234 992631 331262 1005147
rect 357044 1005105 357100 1005114
rect 364244 1005170 364300 1005179
rect 364244 1005105 364246 1005114
rect 364298 1005105 364300 1005114
rect 364246 1005073 364298 1005079
rect 357622 1003873 357674 1003879
rect 357620 1003838 357622 1003847
rect 357674 1003838 357676 1003847
rect 357620 1003773 357676 1003782
rect 359060 1003838 359116 1003847
rect 359060 1003773 359062 1003782
rect 359114 1003773 359116 1003782
rect 359062 1003741 359114 1003747
rect 355990 1003725 356042 1003731
rect 355988 1003690 355990 1003699
rect 356042 1003690 356044 1003699
rect 355988 1003625 356044 1003634
rect 361558 1000913 361610 1000919
rect 360692 1000878 360748 1000887
rect 360692 1000813 360694 1000822
rect 360746 1000813 360748 1000822
rect 361556 1000878 361558 1000887
rect 361610 1000878 361612 1000887
rect 361556 1000813 361612 1000822
rect 360694 1000781 360746 1000787
rect 331798 999433 331850 999439
rect 331798 999375 331850 999381
rect 331810 997885 331838 999375
rect 366274 999291 366302 1005295
rect 381718 1005279 381770 1005285
rect 381718 1005221 381770 1005227
rect 368566 1005205 368618 1005211
rect 368566 1005147 368618 1005153
rect 368578 999365 368606 1005147
rect 380086 1003873 380138 1003879
rect 380086 1003815 380138 1003821
rect 378262 1003799 378314 1003805
rect 378262 1003741 378314 1003747
rect 378274 1001955 378302 1003741
rect 379318 1003725 379370 1003731
rect 379318 1003667 379370 1003673
rect 378262 1001949 378314 1001955
rect 378262 1001891 378314 1001897
rect 368566 999359 368618 999365
rect 368566 999301 368618 999307
rect 366262 999285 366314 999291
rect 366262 999227 366314 999233
rect 367894 997953 367946 997959
rect 367892 997918 367894 997927
rect 367946 997918 367948 997927
rect 331798 997879 331850 997885
rect 367892 997853 367948 997862
rect 331798 997821 331850 997827
rect 348694 997805 348746 997811
rect 348694 997747 348746 997753
rect 369044 997770 369100 997779
rect 348706 995855 348734 997747
rect 369044 997705 369046 997714
rect 369098 997705 369100 997714
rect 369046 997673 369098 997679
rect 367126 996473 367178 996479
rect 367126 996415 367178 996421
rect 367138 996035 367166 996415
rect 368662 996177 368714 996183
rect 368662 996119 368714 996125
rect 367126 996029 367178 996035
rect 362324 995994 362380 996003
rect 362324 995929 362380 995938
rect 367124 995994 367126 996003
rect 367178 995994 367180 996003
rect 367124 995929 367180 995938
rect 348692 995846 348748 995855
rect 348692 995781 348748 995790
rect 339764 995254 339820 995263
rect 339764 995189 339820 995198
rect 339778 994967 339806 995189
rect 339764 994958 339820 994967
rect 339764 994893 339820 994902
rect 362338 993667 362366 995929
rect 365876 995846 365932 995855
rect 365876 995781 365932 995790
rect 366644 995846 366700 995855
rect 366644 995781 366646 995790
rect 365890 995739 365918 995781
rect 366698 995781 366700 995790
rect 366646 995749 366698 995755
rect 365878 995733 365930 995739
rect 368674 995707 368702 996119
rect 379330 996003 379358 1003667
rect 380098 999384 380126 1003815
rect 380470 1001949 380522 1001955
rect 380470 1001891 380522 1001897
rect 380098 999356 380318 999384
rect 380182 997953 380234 997959
rect 380182 997895 380234 997901
rect 380194 996109 380222 997895
rect 380182 996103 380234 996109
rect 380182 996045 380234 996051
rect 377300 995994 377356 996003
rect 377300 995929 377356 995938
rect 379316 995994 379372 996003
rect 379316 995929 379372 995938
rect 371828 995846 371884 995855
rect 371828 995781 371830 995790
rect 371882 995781 371884 995790
rect 371830 995749 371882 995755
rect 365878 995675 365930 995681
rect 368660 995698 368716 995707
rect 368660 995633 368716 995642
rect 374420 995698 374476 995707
rect 374420 995633 374476 995642
rect 362804 995254 362860 995263
rect 362804 995189 362860 995198
rect 368468 995254 368524 995263
rect 368468 995189 368524 995198
rect 362818 995115 362846 995189
rect 362804 995106 362860 995115
rect 362804 995041 362860 995050
rect 368482 994819 368510 995189
rect 368468 994810 368524 994819
rect 368468 994745 368524 994754
rect 362326 993661 362378 993667
rect 362326 993603 362378 993609
rect 331222 992625 331274 992631
rect 331222 992567 331274 992573
rect 332566 992625 332618 992631
rect 332566 992567 332618 992573
rect 328246 989369 328298 989375
rect 328246 989311 328298 989317
rect 300502 989295 300554 989301
rect 300502 989237 300554 989243
rect 325270 989295 325322 989301
rect 325270 989237 325322 989243
rect 288022 988703 288074 988709
rect 288022 988645 288074 988651
rect 299158 988703 299210 988709
rect 299158 988645 299210 988651
rect 288034 985157 288062 988645
rect 288022 985151 288074 985157
rect 288022 985093 288074 985099
rect 300514 983534 300542 989237
rect 316726 988111 316778 988117
rect 316726 988053 316778 988059
rect 316738 983534 316766 988053
rect 332578 983548 332606 992567
rect 374434 989449 374462 995633
rect 374516 995550 374572 995559
rect 374516 995485 374572 995494
rect 374422 989443 374474 989449
rect 374422 989385 374474 989391
rect 349174 989369 349226 989375
rect 349174 989311 349226 989317
rect 277942 983523 277994 983529
rect 332578 983520 332976 983548
rect 349186 983534 349214 989311
rect 374530 989301 374558 995485
rect 377314 989375 377342 995929
rect 377398 995733 377450 995739
rect 377398 995675 377450 995681
rect 377410 995411 377438 995675
rect 380290 995559 380318 999356
rect 380276 995550 380332 995559
rect 380482 995517 380510 1001891
rect 381730 995707 381758 1005221
rect 382966 1005131 383018 1005137
rect 382966 1005073 383018 1005079
rect 382978 995887 383006 1005073
rect 383650 1001012 383678 1005443
rect 430868 1005401 430870 1005410
rect 430922 1005401 430924 1005410
rect 433172 1005466 433174 1005475
rect 433226 1005466 433228 1005475
rect 433172 1005401 433228 1005410
rect 430870 1005369 430922 1005375
rect 431542 1005353 431594 1005359
rect 425300 1005318 425356 1005327
rect 425300 1005253 425302 1005262
rect 425354 1005253 425356 1005262
rect 431540 1005318 431542 1005327
rect 431594 1005318 431596 1005327
rect 431540 1005253 431596 1005262
rect 425302 1005221 425354 1005227
rect 427606 1005205 427658 1005211
rect 427604 1005170 427606 1005179
rect 427658 1005170 427660 1005179
rect 427604 1005105 427660 1005114
rect 435572 1005170 435628 1005179
rect 435572 1005105 435574 1005114
rect 435626 1005105 435628 1005114
rect 435574 1005073 435626 1005079
rect 428084 1003986 428140 1003995
rect 428084 1003921 428086 1003930
rect 428138 1003921 428140 1003930
rect 428086 1003889 428138 1003895
rect 426454 1003873 426506 1003879
rect 423380 1003838 423436 1003847
rect 423380 1003773 423382 1003782
rect 423434 1003773 423436 1003782
rect 426452 1003838 426454 1003847
rect 426506 1003838 426508 1003847
rect 426452 1003773 426508 1003782
rect 423382 1003741 423434 1003747
rect 425782 1003725 425834 1003731
rect 425780 1003690 425782 1003699
rect 425834 1003690 425836 1003699
rect 425780 1003625 425836 1003634
rect 434036 1001174 434092 1001183
rect 434036 1001109 434038 1001118
rect 434090 1001109 434092 1001118
rect 434038 1001077 434090 1001083
rect 432500 1001026 432556 1001035
rect 383650 1000984 383774 1001012
rect 383638 1000913 383690 1000919
rect 383638 1000855 383690 1000861
rect 383542 1000839 383594 1000845
rect 383542 1000781 383594 1000787
rect 383062 999359 383114 999365
rect 383062 999301 383114 999307
rect 382966 995881 383018 995887
rect 382966 995823 383018 995829
rect 381716 995698 381772 995707
rect 381716 995633 381772 995642
rect 383074 995591 383102 999301
rect 383254 999285 383306 999291
rect 383254 999227 383306 999233
rect 383158 997879 383210 997885
rect 383158 997821 383210 997827
rect 383062 995585 383114 995591
rect 383062 995527 383114 995533
rect 380276 995485 380332 995494
rect 380470 995511 380522 995517
rect 380470 995453 380522 995459
rect 377396 995402 377452 995411
rect 377396 995337 377452 995346
rect 383170 995147 383198 997821
rect 383158 995141 383210 995147
rect 383266 995115 383294 999227
rect 383554 995739 383582 1000781
rect 383650 995813 383678 1000855
rect 383638 995807 383690 995813
rect 383638 995749 383690 995755
rect 383542 995733 383594 995739
rect 383542 995675 383594 995681
rect 383746 995665 383774 1000984
rect 432500 1000961 432502 1000970
rect 432554 1000961 432556 1000970
rect 432502 1000929 432554 1000935
rect 428950 1000913 429002 1000919
rect 424148 1000878 424204 1000887
rect 424148 1000813 424150 1000822
rect 424202 1000813 424204 1000822
rect 428948 1000878 428950 1000887
rect 429002 1000878 429004 1000887
rect 428948 1000813 429004 1000822
rect 424150 1000781 424202 1000787
rect 399958 999433 400010 999439
rect 399958 999375 400010 999381
rect 399860 996142 399916 996151
rect 399860 996077 399916 996086
rect 385844 995846 385900 995855
rect 384994 995813 385296 995832
rect 384982 995807 385296 995813
rect 385034 995804 385296 995807
rect 389108 995846 389164 995855
rect 385900 995804 385968 995832
rect 387490 995813 387792 995832
rect 387478 995807 387792 995813
rect 385844 995781 385900 995790
rect 384982 995749 385034 995755
rect 387530 995804 387792 995807
rect 388992 995804 389108 995832
rect 389108 995781 389164 995790
rect 393716 995846 393772 995855
rect 393772 995804 393984 995832
rect 396336 995813 396638 995832
rect 396336 995807 396650 995813
rect 396336 995804 396598 995807
rect 393716 995781 393772 995790
rect 387478 995749 387530 995755
rect 396598 995749 396650 995755
rect 388054 995733 388106 995739
rect 384418 995665 384672 995684
rect 389396 995698 389452 995707
rect 388106 995681 388368 995684
rect 388054 995675 388368 995681
rect 383734 995659 383786 995665
rect 383734 995601 383786 995607
rect 384406 995659 384672 995665
rect 384458 995656 384672 995659
rect 388066 995656 388368 995675
rect 389452 995656 389664 995684
rect 389396 995633 389452 995642
rect 384406 995601 384458 995607
rect 392374 995585 392426 995591
rect 386324 995550 386380 995559
rect 391796 995550 391852 995559
rect 386324 995485 386380 995494
rect 386338 995263 386366 995485
rect 386324 995254 386380 995263
rect 386324 995189 386380 995198
rect 383158 995083 383210 995089
rect 383252 995106 383308 995115
rect 383252 995041 383308 995050
rect 390178 993593 390206 995522
rect 390850 994227 390878 995522
rect 391852 995508 392112 995536
rect 392426 995533 392688 995536
rect 392374 995527 392688 995533
rect 392386 995508 392688 995527
rect 393058 995508 393312 995536
rect 394882 995517 395184 995536
rect 394870 995511 395184 995517
rect 391796 995485 391852 995494
rect 393058 995115 393086 995508
rect 394922 995508 395184 995511
rect 396706 995508 397008 995536
rect 394870 995453 394922 995459
rect 396706 995411 396734 995508
rect 396692 995402 396748 995411
rect 396692 995337 396748 995346
rect 393044 995106 393100 995115
rect 393044 995041 393100 995050
rect 390836 994218 390892 994227
rect 390836 994153 390892 994162
rect 398818 993667 398846 995522
rect 399874 994819 399902 996077
rect 399970 995813 399998 999375
rect 422518 999359 422570 999365
rect 422518 999301 422570 999307
rect 429142 999359 429194 999365
rect 429142 999301 429194 999307
rect 422530 995855 422558 999301
rect 422516 995846 422572 995855
rect 399958 995807 400010 995813
rect 422516 995781 422572 995790
rect 399958 995749 400010 995755
rect 399860 994810 399916 994819
rect 399860 994745 399916 994754
rect 398806 993661 398858 993667
rect 398806 993603 398858 993609
rect 390166 993587 390218 993593
rect 390166 993529 390218 993535
rect 397846 989443 397898 989449
rect 397846 989385 397898 989391
rect 377302 989369 377354 989375
rect 377302 989311 377354 989317
rect 365398 989295 365450 989301
rect 365398 989237 365450 989243
rect 374518 989295 374570 989301
rect 374518 989237 374570 989243
rect 365410 983534 365438 989237
rect 381622 988037 381674 988043
rect 381622 987979 381674 987985
rect 381634 983534 381662 987979
rect 397858 983534 397886 989385
rect 414070 989369 414122 989375
rect 414070 989311 414122 989317
rect 414082 983534 414110 989311
rect 429154 983529 429182 999301
rect 436340 996290 436396 996299
rect 436340 996225 436396 996234
rect 436354 996183 436382 996225
rect 436342 996177 436394 996183
rect 436438 996177 436490 996183
rect 436342 996119 436394 996125
rect 436436 996142 436438 996151
rect 436490 996142 436492 996151
rect 436436 996077 436492 996086
rect 439234 996035 439262 1005517
rect 440674 1005137 440702 1005665
rect 446422 1005575 446474 1005581
rect 446422 1005517 446474 1005523
rect 446038 1005427 446090 1005433
rect 446038 1005369 446090 1005375
rect 440662 1005131 440714 1005137
rect 440662 1005073 440714 1005079
rect 440674 996109 440702 1005073
rect 446050 1002325 446078 1005369
rect 446434 1005359 446462 1005517
rect 446626 1005433 446654 1005665
rect 460822 1005501 460874 1005507
rect 558742 1005501 558794 1005507
rect 460822 1005443 460874 1005449
rect 554516 1005466 554572 1005475
rect 446614 1005427 446666 1005433
rect 446614 1005369 446666 1005375
rect 446326 1005353 446378 1005359
rect 446326 1005295 446378 1005301
rect 446422 1005353 446474 1005359
rect 446422 1005295 446474 1005301
rect 446338 1002344 446366 1005295
rect 457846 1003947 457898 1003953
rect 457846 1003889 457898 1003895
rect 456310 1003873 456362 1003879
rect 456310 1003815 456362 1003821
rect 446038 1002319 446090 1002325
rect 446338 1002316 446462 1002344
rect 446038 1002261 446090 1002267
rect 446434 1001067 446462 1002316
rect 446518 1002319 446570 1002325
rect 446518 1002261 446570 1002267
rect 446530 1001215 446558 1002261
rect 446518 1001209 446570 1001215
rect 446518 1001151 446570 1001157
rect 446422 1001061 446474 1001067
rect 446422 1001003 446474 1001009
rect 456322 1000327 456350 1003815
rect 457858 1002196 457886 1003889
rect 457858 1002168 457982 1002196
rect 456310 1000321 456362 1000327
rect 456310 1000263 456362 1000269
rect 457954 997737 457982 1002168
rect 458806 1000321 458858 1000327
rect 458806 1000263 458858 1000269
rect 457942 997731 457994 997737
rect 457942 997673 457994 997679
rect 458818 996849 458846 1000263
rect 460834 999143 460862 1005443
rect 469846 1005427 469898 1005433
rect 558742 1005443 558794 1005449
rect 572854 1005501 572906 1005507
rect 572854 1005443 572906 1005449
rect 554516 1005401 554518 1005410
rect 469846 1005369 469898 1005375
rect 554570 1005401 554572 1005410
rect 554518 1005369 554570 1005375
rect 463606 1005279 463658 1005285
rect 463606 1005221 463658 1005227
rect 463618 1005008 463646 1005221
rect 466582 1005205 466634 1005211
rect 466582 1005147 466634 1005153
rect 463618 1004980 463742 1005008
rect 463714 1000771 463742 1004980
rect 466486 1003799 466538 1003805
rect 466486 1003741 466538 1003747
rect 463702 1000765 463754 1000771
rect 463702 1000707 463754 1000713
rect 466498 999236 466526 1003741
rect 466594 999513 466622 1005147
rect 467062 1001209 467114 1001215
rect 467062 1001151 467114 1001157
rect 466582 999507 466634 999513
rect 466582 999449 466634 999455
rect 466498 999208 466622 999236
rect 460822 999137 460874 999143
rect 460822 999079 460874 999085
rect 458806 996843 458858 996849
rect 458806 996785 458858 996791
rect 440662 996103 440714 996109
rect 440662 996045 440714 996051
rect 434134 996029 434186 996035
rect 429716 995994 429772 996003
rect 429716 995929 429772 995938
rect 434132 995994 434134 996003
rect 439222 996029 439274 996035
rect 434186 995994 434188 996003
rect 439222 995971 439274 995977
rect 446228 995994 446284 996003
rect 434132 995929 434188 995938
rect 446228 995929 446284 995938
rect 429730 993667 429758 995929
rect 438740 995846 438796 995855
rect 438740 995781 438742 995790
rect 438794 995781 438796 995790
rect 444502 995807 444554 995813
rect 438742 995749 438794 995755
rect 444502 995749 444554 995755
rect 440756 995698 440812 995707
rect 440756 995633 440812 995642
rect 429718 993661 429770 993667
rect 429718 993603 429770 993609
rect 440770 989301 440798 995633
rect 443542 995289 443594 995295
rect 443540 995254 443542 995263
rect 443594 995254 443596 995263
rect 443540 995189 443596 995198
rect 444514 990559 444542 995749
rect 444502 990553 444554 990559
rect 444502 990495 444554 990501
rect 446242 989375 446270 995929
rect 466594 995517 466622 999208
rect 467074 995707 467102 1001151
rect 469858 996035 469886 1005369
rect 470038 1005353 470090 1005359
rect 556918 1005353 556970 1005359
rect 470038 1005295 470090 1005301
rect 500660 1005318 500716 1005327
rect 470050 996109 470078 1005295
rect 556916 1005318 556918 1005327
rect 556970 1005318 556972 1005327
rect 500660 1005253 500662 1005262
rect 500714 1005253 500716 1005262
rect 512566 1005279 512618 1005285
rect 500662 1005221 500714 1005227
rect 556916 1005253 556972 1005262
rect 512566 1005221 512618 1005227
rect 501142 1005205 501194 1005211
rect 498164 1005170 498220 1005179
rect 498164 1005105 498220 1005114
rect 501140 1005170 501142 1005179
rect 512470 1005205 512522 1005211
rect 501194 1005170 501196 1005179
rect 512470 1005147 512522 1005153
rect 501140 1005105 501196 1005114
rect 498178 1003805 498206 1005105
rect 498166 1003799 498218 1003805
rect 498166 1003741 498218 1003747
rect 471766 1003725 471818 1003731
rect 471766 1003667 471818 1003673
rect 471670 999433 471722 999439
rect 471670 999375 471722 999381
rect 470038 996103 470090 996109
rect 470038 996045 470090 996051
rect 469846 996029 469898 996035
rect 469846 995971 469898 995977
rect 467060 995698 467116 995707
rect 467060 995633 467116 995642
rect 466582 995511 466634 995517
rect 466582 995453 466634 995459
rect 463604 995402 463660 995411
rect 463604 995337 463660 995346
rect 463618 995295 463646 995337
rect 463606 995289 463658 995295
rect 463606 995231 463658 995237
rect 471682 995221 471710 999375
rect 471778 995411 471806 1003667
rect 501046 1002615 501098 1002621
rect 501046 1002557 501098 1002563
rect 472642 1001141 472766 1001160
rect 472630 1001135 472766 1001141
rect 472682 1001132 472766 1001135
rect 472630 1001077 472682 1001083
rect 472342 1001061 472394 1001067
rect 472342 1001003 472394 1001009
rect 471958 1000839 472010 1000845
rect 471958 1000781 472010 1000787
rect 471862 999137 471914 999143
rect 471862 999079 471914 999085
rect 471874 996003 471902 999079
rect 471860 995994 471916 996003
rect 471860 995929 471916 995938
rect 471970 995443 471998 1000781
rect 472150 1000765 472202 1000771
rect 472150 1000707 472202 1000713
rect 472054 996843 472106 996849
rect 472054 996785 472106 996791
rect 472066 995961 472094 996785
rect 472054 995955 472106 995961
rect 472054 995897 472106 995903
rect 472162 995559 472190 1000707
rect 472246 997731 472298 997737
rect 472246 997673 472298 997679
rect 472258 995855 472286 997673
rect 472244 995846 472300 995855
rect 472244 995781 472300 995790
rect 472354 995591 472382 1001003
rect 472630 1000987 472682 1000993
rect 472630 1000929 472682 1000935
rect 472534 1000913 472586 1000919
rect 472534 1000855 472586 1000861
rect 472438 999507 472490 999513
rect 472438 999449 472490 999455
rect 472450 995887 472478 999449
rect 472438 995881 472490 995887
rect 472438 995823 472490 995829
rect 472546 995739 472574 1000855
rect 472642 995813 472670 1000929
rect 472630 995807 472682 995813
rect 472630 995749 472682 995755
rect 472534 995733 472586 995739
rect 472534 995675 472586 995681
rect 472738 995665 472766 1001132
rect 488950 999433 489002 999439
rect 488852 999398 488908 999407
rect 488950 999375 489002 999381
rect 497588 999398 497644 999407
rect 488852 999333 488908 999342
rect 477044 995846 477100 995855
rect 473314 995813 473664 995832
rect 473302 995807 473664 995813
rect 473354 995804 473664 995807
rect 485780 995846 485836 995855
rect 477100 995804 477360 995832
rect 477730 995813 477984 995832
rect 483874 995813 484176 995832
rect 477718 995807 477984 995813
rect 477044 995781 477100 995790
rect 473302 995749 473354 995755
rect 477770 995804 477984 995807
rect 483862 995807 484176 995813
rect 477718 995749 477770 995755
rect 483914 995804 484176 995807
rect 485376 995813 485726 995832
rect 485376 995807 485738 995813
rect 485376 995804 485686 995807
rect 483862 995749 483914 995755
rect 485836 995804 486000 995832
rect 485780 995781 485836 995790
rect 485686 995749 485738 995755
rect 474070 995733 474122 995739
rect 480980 995698 481036 995707
rect 474122 995681 474336 995684
rect 474070 995675 474336 995681
rect 472726 995659 472778 995665
rect 474082 995656 474336 995675
rect 474658 995665 474960 995684
rect 474646 995659 474960 995665
rect 472726 995601 472778 995607
rect 474698 995656 474960 995659
rect 481036 995656 481104 995684
rect 480980 995633 481036 995642
rect 474646 995601 474698 995607
rect 472342 995585 472394 995591
rect 472148 995550 472204 995559
rect 472342 995527 472394 995533
rect 476374 995585 476426 995591
rect 488866 995559 488894 999333
rect 488962 995813 488990 999375
rect 497588 999333 497590 999342
rect 497642 999333 497644 999342
rect 497590 999301 497642 999307
rect 488950 995807 489002 995813
rect 488950 995749 489002 995755
rect 478388 995550 478444 995559
rect 476426 995533 476784 995536
rect 476374 995527 476784 995533
rect 476386 995508 476784 995527
rect 472148 995485 472204 995494
rect 479924 995550 479980 995559
rect 478444 995508 478656 995536
rect 479856 995522 479924 995536
rect 478388 995485 478444 995494
rect 471958 995437 472010 995443
rect 471764 995402 471820 995411
rect 471958 995379 472010 995385
rect 471764 995337 471820 995346
rect 471670 995215 471722 995221
rect 471670 995157 471722 995163
rect 479170 993593 479198 995522
rect 479842 995508 479924 995522
rect 479842 994227 479870 995508
rect 488852 995550 488908 995559
rect 479924 995485 479980 995494
rect 481378 995508 481680 995536
rect 482050 995508 482352 995536
rect 482722 995517 482976 995536
rect 482710 995511 482976 995517
rect 481378 995443 481406 995508
rect 481366 995437 481418 995443
rect 482050 995411 482078 995508
rect 482762 995508 482976 995511
rect 482710 995453 482762 995459
rect 481366 995379 481418 995385
rect 482036 995402 482092 995411
rect 482036 995337 482092 995346
rect 479828 994218 479884 994227
rect 479828 994153 479884 994162
rect 487810 993667 487838 995522
rect 488852 995485 488908 995494
rect 487798 993661 487850 993667
rect 487798 993603 487850 993609
rect 501058 993593 501086 1002557
rect 503446 1002541 503498 1002547
rect 503444 1002506 503446 1002515
rect 503498 1002506 503500 1002515
rect 503444 1002441 503500 1002450
rect 505076 1002358 505132 1002367
rect 505076 1002293 505078 1002302
rect 505130 1002293 505132 1002302
rect 505078 1002261 505130 1002267
rect 509396 1000730 509452 1000739
rect 509396 1000665 509398 1000674
rect 509450 1000665 509452 1000674
rect 509398 1000633 509450 1000639
rect 503060 999990 503116 999999
rect 503060 999925 503062 999934
rect 503114 999925 503116 999934
rect 503062 999893 503114 999899
rect 509876 999842 509932 999851
rect 509876 999777 509878 999786
rect 509930 999777 509932 999786
rect 509878 999745 509930 999751
rect 506230 999729 506282 999735
rect 506228 999694 506230 999703
rect 506282 999694 506284 999703
rect 506228 999629 506284 999638
rect 507764 999694 507820 999703
rect 507764 999629 507766 999638
rect 507818 999629 507820 999638
rect 507766 999597 507818 999603
rect 502390 999581 502442 999587
rect 502388 999546 502390 999555
rect 502442 999546 502444 999555
rect 502388 999481 502444 999490
rect 508628 999546 508684 999555
rect 508628 999481 508630 999490
rect 508682 999481 508684 999490
rect 508630 999449 508682 999455
rect 512482 999291 512510 1005147
rect 512578 999384 512606 1005221
rect 558754 1005211 558782 1005443
rect 570454 1005427 570506 1005433
rect 570454 1005369 570506 1005375
rect 553750 1005205 553802 1005211
rect 553748 1005170 553750 1005179
rect 558742 1005205 558794 1005211
rect 553802 1005170 553804 1005179
rect 562486 1005205 562538 1005211
rect 558742 1005147 558794 1005153
rect 562484 1005170 562486 1005179
rect 562538 1005170 562540 1005179
rect 553748 1005105 553804 1005114
rect 562484 1005105 562540 1005114
rect 554902 1003873 554954 1003879
rect 554900 1003838 554902 1003847
rect 567190 1003873 567242 1003879
rect 554954 1003838 554956 1003847
rect 515734 1003799 515786 1003805
rect 567190 1003815 567242 1003821
rect 554900 1003773 554956 1003782
rect 515734 1003741 515786 1003747
rect 512578 999356 512702 999384
rect 512470 999285 512522 999291
rect 512470 999227 512522 999233
rect 512674 996553 512702 999356
rect 512662 996547 512714 996553
rect 512662 996489 512714 996495
rect 511894 996251 511946 996257
rect 511894 996193 511946 996199
rect 511124 996142 511180 996151
rect 511124 996077 511126 996086
rect 511178 996077 511180 996086
rect 511126 996045 511178 996051
rect 511906 996035 511934 996193
rect 513430 996177 513482 996183
rect 513428 996142 513430 996151
rect 513482 996142 513484 996151
rect 513428 996077 513484 996086
rect 511894 996029 511946 996035
rect 511892 995994 511894 996003
rect 513334 996029 513386 996035
rect 511946 995994 511948 996003
rect 511892 995929 511948 995938
rect 513332 995994 513334 996003
rect 513386 995994 513388 996003
rect 513332 995929 513388 995938
rect 504692 995846 504748 995855
rect 504692 995781 504694 995790
rect 504746 995781 504748 995790
rect 504694 995749 504746 995755
rect 515746 995295 515774 1003741
rect 555670 1003725 555722 1003731
rect 555668 1003690 555670 1003699
rect 555722 1003690 555724 1003699
rect 555668 1003625 555724 1003634
rect 519286 1002615 519338 1002621
rect 519286 1002557 519338 1002563
rect 517174 1002393 517226 1002399
rect 517174 1002335 517226 1002341
rect 516694 1000691 516746 1000697
rect 516694 1000633 516746 1000639
rect 516706 1000295 516734 1000633
rect 516692 1000286 516748 1000295
rect 516692 1000221 516748 1000230
rect 516694 999951 516746 999957
rect 516694 999893 516746 999899
rect 516706 999407 516734 999893
rect 516884 999842 516940 999851
rect 516884 999777 516940 999786
rect 516790 999729 516842 999735
rect 516788 999694 516790 999703
rect 516842 999694 516844 999703
rect 516788 999629 516844 999638
rect 516790 999581 516842 999587
rect 516788 999546 516790 999555
rect 516842 999546 516844 999555
rect 516788 999481 516844 999490
rect 516692 999398 516748 999407
rect 516898 999365 516926 999777
rect 516692 999333 516748 999342
rect 516886 999359 516938 999365
rect 516886 999301 516938 999307
rect 517186 996151 517214 1002335
rect 517172 996142 517228 996151
rect 517172 996077 517228 996086
rect 518710 995807 518762 995813
rect 518710 995749 518762 995755
rect 518722 995707 518750 995749
rect 518516 995698 518572 995707
rect 518516 995633 518572 995642
rect 518708 995698 518764 995707
rect 518708 995633 518764 995642
rect 515734 995289 515786 995295
rect 506612 995254 506668 995263
rect 515734 995231 515786 995237
rect 506612 995189 506668 995198
rect 506626 993741 506654 995189
rect 509684 995106 509740 995115
rect 509740 995064 509918 995092
rect 509684 995041 509740 995050
rect 509890 994819 509918 995064
rect 509876 994810 509932 994819
rect 509876 994745 509932 994754
rect 506614 993735 506666 993741
rect 506614 993677 506666 993683
rect 479158 993587 479210 993593
rect 479158 993529 479210 993535
rect 501046 993587 501098 993593
rect 501046 993529 501098 993535
rect 462742 990553 462794 990559
rect 462742 990495 462794 990501
rect 446230 989369 446282 989375
rect 446230 989311 446282 989317
rect 430294 989295 430346 989301
rect 430294 989237 430346 989243
rect 440758 989295 440810 989301
rect 440758 989237 440810 989243
rect 430306 983534 430334 989237
rect 446518 987963 446570 987969
rect 446518 987905 446570 987911
rect 446530 983534 446558 987905
rect 462754 983534 462782 990495
rect 518530 989375 518558 995633
rect 518708 995550 518764 995559
rect 518708 995485 518764 995494
rect 478966 989369 479018 989375
rect 478966 989311 479018 989317
rect 518518 989369 518570 989375
rect 518518 989311 518570 989317
rect 478978 983534 479006 989311
rect 518722 989301 518750 995485
rect 519298 994967 519326 1002557
rect 559126 1002541 559178 1002547
rect 559124 1002506 559126 1002515
rect 566134 1002541 566186 1002547
rect 559178 1002506 559180 1002515
rect 559124 1002441 559180 1002450
rect 560564 1002506 560620 1002515
rect 566134 1002483 566186 1002489
rect 560564 1002441 560566 1002450
rect 560618 1002441 560620 1002450
rect 560566 1002409 560618 1002415
rect 560086 1002393 560138 1002399
rect 560084 1002358 560086 1002367
rect 564694 1002393 564746 1002399
rect 560138 1002358 560140 1002367
rect 523606 1002319 523658 1002325
rect 560084 1002293 560140 1002302
rect 561524 1002358 561580 1002367
rect 564790 1002393 564842 1002399
rect 564694 1002335 564746 1002341
rect 564788 1002358 564790 1002367
rect 564842 1002358 564844 1002367
rect 561524 1002293 561526 1002302
rect 523606 1002261 523658 1002267
rect 561578 1002293 561580 1002302
rect 561526 1002261 561578 1002267
rect 523508 999842 523564 999851
rect 521686 999803 521738 999809
rect 523508 999777 523564 999786
rect 521686 999745 521738 999751
rect 521590 999655 521642 999661
rect 521590 999597 521642 999603
rect 521302 999359 521354 999365
rect 521302 999301 521354 999307
rect 521314 995369 521342 999301
rect 521494 996547 521546 996553
rect 521494 996489 521546 996495
rect 521396 995994 521452 996003
rect 521396 995929 521452 995938
rect 521302 995363 521354 995369
rect 521302 995305 521354 995311
rect 519284 994958 519340 994967
rect 519284 994893 519340 994902
rect 521410 989523 521438 995929
rect 521506 995559 521534 996489
rect 521602 996003 521630 999597
rect 521588 995994 521644 996003
rect 521588 995929 521644 995938
rect 521492 995550 521548 995559
rect 521492 995485 521548 995494
rect 521698 995263 521726 999745
rect 521782 999285 521834 999291
rect 521782 999227 521834 999233
rect 521794 995517 521822 999227
rect 521782 995511 521834 995517
rect 521782 995453 521834 995459
rect 523522 995443 523550 999777
rect 523618 995665 523646 1002261
rect 564706 1001067 564734 1002335
rect 564788 1002293 564844 1002302
rect 565174 1002319 565226 1002325
rect 565174 1002261 565226 1002267
rect 564694 1001061 564746 1001067
rect 564694 1001003 564746 1001009
rect 565186 1000919 565214 1002261
rect 565174 1000913 565226 1000919
rect 565174 1000855 565226 1000861
rect 523796 1000286 523852 1000295
rect 523796 1000221 523852 1000230
rect 523700 999546 523756 999555
rect 523700 999481 523756 999490
rect 523714 995887 523742 999481
rect 523702 995881 523754 995887
rect 523702 995823 523754 995829
rect 523810 995739 523838 1000221
rect 523892 999694 523948 999703
rect 523892 999629 523948 999638
rect 540310 999655 540362 999661
rect 523906 995813 523934 999629
rect 540310 999597 540362 999603
rect 523990 999507 524042 999513
rect 523990 999449 524042 999455
rect 524002 995855 524030 999449
rect 524084 999398 524140 999407
rect 524084 999333 524140 999342
rect 524098 995961 524126 999333
rect 524086 995955 524138 995961
rect 524086 995897 524138 995903
rect 523988 995846 524044 995855
rect 523894 995807 523946 995813
rect 527924 995846 527980 995855
rect 525346 995813 525744 995832
rect 523988 995781 524044 995790
rect 525334 995807 525744 995813
rect 523894 995749 523946 995755
rect 525386 995804 525744 995807
rect 532244 995846 532300 995855
rect 527980 995804 528192 995832
rect 529858 995813 530064 995832
rect 529846 995807 530064 995813
rect 527924 995781 527980 995790
rect 525334 995749 525386 995755
rect 529898 995804 530064 995807
rect 535316 995846 535372 995855
rect 532300 995804 532512 995832
rect 533410 995813 533712 995832
rect 533398 995807 533712 995813
rect 532244 995781 532300 995790
rect 529846 995749 529898 995755
rect 533450 995804 533712 995807
rect 535372 995804 535584 995832
rect 536784 995813 537182 995832
rect 540322 995813 540350 999597
rect 552982 999433 553034 999439
rect 552980 999398 552982 999407
rect 555862 999433 555914 999439
rect 553034 999398 553036 999407
rect 555862 999375 555914 999381
rect 552980 999333 553036 999342
rect 555874 996553 555902 999375
rect 566146 999291 566174 1002483
rect 566422 1002467 566474 1002473
rect 566422 1002409 566474 1002415
rect 566134 999285 566186 999291
rect 566134 999227 566186 999233
rect 557300 997918 557356 997927
rect 557300 997853 557302 997862
rect 557354 997853 557356 997862
rect 557302 997821 557354 997827
rect 566434 997811 566462 1002409
rect 567202 999217 567230 1003815
rect 567286 1003725 567338 1003731
rect 567286 1003667 567338 1003673
rect 567298 999384 567326 1003667
rect 567670 1002393 567722 1002399
rect 567670 1002335 567722 1002341
rect 567298 999356 567422 999384
rect 567190 999211 567242 999217
rect 567190 999153 567242 999159
rect 567394 998625 567422 999356
rect 567382 998619 567434 998625
rect 567382 998561 567434 998567
rect 566422 997805 566474 997811
rect 566422 997747 566474 997753
rect 555862 996547 555914 996553
rect 555862 996489 555914 996495
rect 561430 996547 561482 996553
rect 561430 996489 561482 996495
rect 558164 995846 558220 995855
rect 536784 995807 537194 995813
rect 536784 995804 537142 995807
rect 535316 995781 535372 995790
rect 533398 995749 533450 995755
rect 537142 995749 537194 995755
rect 540310 995807 540362 995813
rect 558164 995781 558220 995790
rect 540310 995749 540362 995755
rect 523798 995733 523850 995739
rect 523798 995675 523850 995681
rect 524758 995733 524810 995739
rect 529076 995698 529132 995707
rect 524810 995681 525072 995684
rect 524758 995675 525072 995681
rect 523606 995659 523658 995665
rect 524770 995656 525072 995675
rect 528418 995665 528768 995684
rect 528406 995659 528768 995665
rect 523606 995601 523658 995607
rect 528458 995656 528768 995659
rect 534068 995698 534124 995707
rect 529132 995656 529392 995684
rect 529076 995633 529132 995642
rect 544244 995698 544300 995707
rect 534124 995656 534384 995684
rect 534068 995633 534124 995642
rect 544244 995633 544300 995642
rect 528406 995601 528458 995607
rect 526114 995508 526368 995536
rect 530592 995508 530750 995536
rect 523510 995437 523562 995443
rect 526114 995411 526142 995508
rect 530722 995411 530750 995508
rect 531106 995522 531216 995536
rect 531106 995508 531230 995522
rect 532834 995517 533088 995536
rect 531106 995443 531134 995508
rect 531094 995437 531146 995443
rect 523510 995379 523562 995385
rect 526100 995402 526156 995411
rect 526100 995337 526156 995346
rect 526484 995402 526540 995411
rect 526484 995337 526540 995346
rect 530708 995402 530764 995411
rect 531094 995379 531146 995385
rect 530708 995337 530764 995346
rect 521684 995254 521740 995263
rect 521684 995189 521740 995198
rect 526498 994967 526526 995337
rect 526484 994958 526540 994967
rect 526484 994893 526540 994902
rect 531202 993667 531230 995508
rect 532822 995511 533088 995517
rect 532874 995508 533088 995511
rect 537154 995508 537408 995536
rect 538978 995508 539232 995536
rect 532822 995453 532874 995459
rect 536852 995402 536908 995411
rect 536852 995337 536908 995346
rect 536866 994227 536894 995337
rect 537154 995263 537182 995508
rect 537140 995254 537196 995263
rect 537140 995189 537196 995198
rect 536852 994218 536908 994227
rect 536852 994153 536908 994162
rect 538978 993741 539006 995508
rect 538966 993735 539018 993741
rect 538966 993677 539018 993683
rect 531190 993661 531242 993667
rect 531190 993603 531242 993609
rect 521398 989517 521450 989523
rect 521398 989459 521450 989465
rect 527638 989369 527690 989375
rect 527638 989311 527690 989317
rect 543766 989369 543818 989375
rect 543766 989311 543818 989317
rect 495190 989295 495242 989301
rect 495190 989237 495242 989243
rect 518710 989295 518762 989301
rect 518710 989237 518762 989243
rect 495202 983534 495230 989237
rect 511414 987889 511466 987895
rect 511414 987831 511466 987837
rect 511426 983534 511454 987831
rect 527650 983534 527678 989311
rect 543778 983534 543806 989311
rect 544258 986415 544286 995633
rect 558178 993889 558206 995781
rect 561442 994375 561470 996489
rect 563734 996177 563786 996183
rect 563734 996119 563786 996125
rect 562870 996103 562922 996109
rect 562870 996045 562922 996051
rect 562882 996003 562910 996045
rect 562868 995994 562924 996003
rect 562868 995929 562924 995938
rect 562882 995887 562910 995929
rect 562870 995881 562922 995887
rect 563746 995855 563774 996119
rect 564790 996029 564842 996035
rect 564788 995994 564790 996003
rect 564842 995994 564844 996003
rect 564788 995929 564844 995938
rect 567092 995994 567148 996003
rect 567092 995929 567094 995938
rect 567146 995929 567148 995938
rect 567094 995897 567146 995903
rect 567382 995881 567434 995887
rect 562870 995823 562922 995829
rect 563732 995846 563788 995855
rect 563732 995781 563788 995790
rect 566324 995846 566380 995855
rect 567382 995823 567434 995829
rect 566324 995781 566326 995790
rect 563746 995739 563774 995781
rect 566378 995781 566380 995790
rect 566326 995749 566378 995755
rect 563734 995733 563786 995739
rect 563734 995675 563786 995681
rect 561718 995437 561770 995443
rect 561620 995402 561676 995411
rect 561718 995379 561770 995385
rect 561620 995337 561676 995346
rect 561634 995240 561662 995337
rect 561730 995240 561758 995379
rect 561634 995212 561758 995240
rect 561526 995067 561578 995073
rect 561526 995009 561578 995015
rect 561428 994366 561484 994375
rect 561428 994301 561484 994310
rect 558166 993883 558218 993889
rect 558166 993825 558218 993831
rect 560086 989295 560138 989301
rect 560086 989237 560138 989243
rect 544246 986409 544298 986415
rect 544246 986351 544298 986357
rect 560098 983534 560126 989237
rect 561538 988265 561566 995009
rect 561526 988259 561578 988265
rect 561526 988201 561578 988207
rect 567394 986563 567422 995823
rect 567478 995733 567530 995739
rect 567478 995675 567530 995681
rect 567382 986557 567434 986563
rect 567382 986499 567434 986505
rect 567490 986489 567518 995675
rect 567682 989301 567710 1002335
rect 570166 1001061 570218 1001067
rect 570166 1001003 570218 1001009
rect 568342 1000913 568394 1000919
rect 568342 1000855 568394 1000861
rect 568354 998329 568382 1000855
rect 568342 998323 568394 998329
rect 568342 998265 568394 998271
rect 570178 997756 570206 1001003
rect 570178 997728 570302 997756
rect 570274 997460 570302 997728
rect 570466 997589 570494 1005369
rect 570550 1005205 570602 1005211
rect 570550 1005147 570602 1005153
rect 570562 997663 570590 1005147
rect 572470 999433 572522 999439
rect 572470 999375 572522 999381
rect 572482 997959 572510 999375
rect 572470 997953 572522 997959
rect 572470 997895 572522 997901
rect 570550 997657 570602 997663
rect 570550 997599 570602 997605
rect 570454 997583 570506 997589
rect 570454 997525 570506 997531
rect 570274 997432 570494 997460
rect 570262 995955 570314 995961
rect 570262 995897 570314 995903
rect 570274 989523 570302 995897
rect 570358 995807 570410 995813
rect 570358 995749 570410 995755
rect 570262 989517 570314 989523
rect 570262 989459 570314 989465
rect 570370 989375 570398 995749
rect 570466 995115 570494 997432
rect 570452 995106 570508 995115
rect 570452 995041 570508 995050
rect 572866 994819 572894 1005443
rect 574486 1005353 574538 1005359
rect 574486 1005295 574538 1005301
rect 573046 999285 573098 999291
rect 573046 999227 573098 999233
rect 572950 998323 573002 998329
rect 572950 998265 573002 998271
rect 572852 994810 572908 994819
rect 572852 994745 572908 994754
rect 572962 994523 572990 998265
rect 573058 996447 573086 999227
rect 574498 997737 574526 1005295
rect 616054 999729 616106 999735
rect 616054 999671 616106 999677
rect 625750 999729 625802 999735
rect 625750 999671 625802 999677
rect 600406 999581 600458 999587
rect 600406 999523 600458 999529
rect 598774 999507 598826 999513
rect 598774 999449 598826 999455
rect 596086 999433 596138 999439
rect 596086 999375 596138 999381
rect 575350 999211 575402 999217
rect 575350 999153 575402 999159
rect 574486 997731 574538 997737
rect 574486 997673 574538 997679
rect 573044 996438 573100 996447
rect 573044 996373 573100 996382
rect 573140 995846 573196 995855
rect 573140 995781 573196 995790
rect 572948 994514 573004 994523
rect 572948 994449 573004 994458
rect 573154 989449 573182 995781
rect 575362 994671 575390 999153
rect 575446 998619 575498 998625
rect 575446 998561 575498 998567
rect 575458 994967 575486 998561
rect 596098 997885 596126 999375
rect 596086 997879 596138 997885
rect 596086 997821 596138 997827
rect 598786 997811 598814 999449
rect 598774 997805 598826 997811
rect 598774 997747 598826 997753
rect 600418 997663 600446 999523
rect 616066 999513 616094 999671
rect 616150 999655 616202 999661
rect 616150 999597 616202 999603
rect 616054 999507 616106 999513
rect 616054 999449 616106 999455
rect 616162 999439 616190 999597
rect 625654 999507 625706 999513
rect 625654 999449 625706 999455
rect 616150 999433 616202 999439
rect 616150 999375 616202 999381
rect 616246 999433 616298 999439
rect 616246 999375 616298 999381
rect 600406 997657 600458 997663
rect 600406 997599 600458 997605
rect 616258 997589 616286 999375
rect 617782 997953 617834 997959
rect 617782 997895 617834 997901
rect 616246 997583 616298 997589
rect 616246 997525 616298 997531
rect 604820 996438 604876 996447
rect 604820 996373 604822 996382
rect 604874 996373 604876 996382
rect 604822 996341 604874 996347
rect 617794 995591 617822 997895
rect 619126 997731 619178 997737
rect 619126 997673 619178 997679
rect 619138 995887 619166 997673
rect 624886 996399 624938 996405
rect 624886 996341 624938 996347
rect 624898 996003 624926 996341
rect 624884 995994 624940 996003
rect 624884 995929 624940 995938
rect 619126 995881 619178 995887
rect 619126 995823 619178 995829
rect 625666 995665 625694 999449
rect 625762 995813 625790 999671
rect 625846 999655 625898 999661
rect 625846 999597 625898 999603
rect 625858 999532 625886 999597
rect 625858 999504 625982 999532
rect 625846 999433 625898 999439
rect 625846 999375 625898 999381
rect 625858 995961 625886 999375
rect 625846 995955 625898 995961
rect 625846 995897 625898 995903
rect 625750 995807 625802 995813
rect 625750 995749 625802 995755
rect 625954 995739 625982 999504
rect 634100 995846 634156 995855
rect 626530 995813 626880 995832
rect 630178 995813 630576 995832
rect 626518 995807 626880 995813
rect 626570 995804 626880 995807
rect 630166 995807 630576 995813
rect 626518 995749 626570 995755
rect 630218 995804 630576 995807
rect 634156 995804 634320 995832
rect 635266 995813 635520 995832
rect 635254 995807 635520 995813
rect 634100 995781 634156 995790
rect 630166 995749 630218 995755
rect 635306 995804 635520 995807
rect 635254 995749 635306 995755
rect 625942 995733 625994 995739
rect 625942 995675 625994 995681
rect 627094 995733 627146 995739
rect 635828 995698 635884 995707
rect 627146 995681 627504 995684
rect 627094 995675 627504 995681
rect 625654 995659 625706 995665
rect 627106 995656 627504 995675
rect 627874 995665 628176 995684
rect 627862 995659 628176 995665
rect 625654 995601 625706 995607
rect 627914 995656 628176 995659
rect 635884 995656 636144 995684
rect 635828 995633 635884 995642
rect 627862 995601 627914 995607
rect 617782 995585 617834 995591
rect 617782 995527 617834 995533
rect 629206 995585 629258 995591
rect 629206 995527 629258 995533
rect 581686 995437 581738 995443
rect 581684 995402 581686 995411
rect 581738 995402 581740 995411
rect 581684 995337 581740 995346
rect 584756 995254 584812 995263
rect 584756 995189 584812 995198
rect 604724 995254 604780 995263
rect 604724 995189 604780 995198
rect 584770 995073 584798 995189
rect 604738 995073 604766 995189
rect 584758 995067 584810 995073
rect 584758 995009 584810 995015
rect 604726 995067 604778 995073
rect 604726 995009 604778 995015
rect 575444 994958 575500 994967
rect 575444 994893 575500 994902
rect 575348 994662 575404 994671
rect 575348 994597 575404 994606
rect 592438 989517 592490 989523
rect 592438 989459 592490 989465
rect 573142 989443 573194 989449
rect 573142 989385 573194 989391
rect 570358 989369 570410 989375
rect 570358 989311 570410 989317
rect 567670 989295 567722 989301
rect 567670 989237 567722 989243
rect 576310 988259 576362 988265
rect 576310 988201 576362 988207
rect 567478 986483 567530 986489
rect 567478 986425 567530 986431
rect 576322 983534 576350 988201
rect 592450 983534 592478 989459
rect 608758 989443 608810 989449
rect 608758 989385 608810 989391
rect 608770 983534 608798 989385
rect 624982 989369 625034 989375
rect 624982 989311 625034 989317
rect 624994 983534 625022 989311
rect 629218 986637 629246 995527
rect 629986 995115 630014 995522
rect 630946 995508 631200 995536
rect 629972 995106 630028 995115
rect 629972 995041 630028 995050
rect 630946 994967 630974 995508
rect 630932 994958 630988 994967
rect 630932 994893 630988 994902
rect 631810 994819 631838 995522
rect 631796 994810 631852 994819
rect 631796 994745 631852 994754
rect 632386 994227 632414 995522
rect 633024 995508 633086 995536
rect 632372 994218 632428 994227
rect 632372 994153 632428 994162
rect 629206 986631 629258 986637
rect 629206 986573 629258 986579
rect 632386 983677 632414 994153
rect 633058 993667 633086 995508
rect 634882 994375 634910 995522
rect 636502 995141 636554 995147
rect 636502 995083 636554 995089
rect 634868 994366 634924 994375
rect 634868 994301 634924 994310
rect 633046 993661 633098 993667
rect 633046 993603 633098 993609
rect 632374 983671 632426 983677
rect 632374 983613 632426 983619
rect 633058 983603 633086 993603
rect 636514 993593 636542 995083
rect 637378 994671 637406 995522
rect 638530 994671 638558 995522
rect 637364 994662 637420 994671
rect 637364 994597 637420 994606
rect 638516 994662 638572 994671
rect 638516 994597 638572 994606
rect 639202 994523 639230 995522
rect 640726 995363 640778 995369
rect 640726 995305 640778 995311
rect 639188 994514 639244 994523
rect 639188 994449 639244 994458
rect 640532 993922 640588 993931
rect 640532 993857 640588 993866
rect 636502 993587 636554 993593
rect 636502 993529 636554 993535
rect 640546 987821 640574 993857
rect 640738 990781 640766 995305
rect 640916 994070 640972 994079
rect 640916 994005 640972 994014
rect 640726 990775 640778 990781
rect 640726 990717 640778 990723
rect 640534 987815 640586 987821
rect 640534 987757 640586 987763
rect 640930 987599 640958 994005
rect 641026 993889 641054 995522
rect 642646 995289 642698 995295
rect 642646 995231 642698 995237
rect 641108 995106 641164 995115
rect 641108 995041 641164 995050
rect 641014 993883 641066 993889
rect 641014 993825 641066 993831
rect 640918 987593 640970 987599
rect 640918 987535 640970 987541
rect 633046 983597 633098 983603
rect 633046 983539 633098 983545
rect 641122 983534 641150 995041
rect 642658 993519 642686 995231
rect 643414 995215 643466 995221
rect 643414 995157 643466 995163
rect 642646 993513 642698 993519
rect 642646 993455 642698 993461
rect 643426 987673 643454 995157
rect 649844 994662 649900 994671
rect 649844 994597 649900 994606
rect 643606 993587 643658 993593
rect 643606 993529 643658 993535
rect 643618 987747 643646 993529
rect 649462 993513 649514 993519
rect 649462 993455 649514 993461
rect 645142 990701 645194 990707
rect 645142 990643 645194 990649
rect 643606 987741 643658 987747
rect 643606 987683 643658 987689
rect 643414 987667 643466 987673
rect 643414 987609 643466 987615
rect 645154 984935 645182 990643
rect 645142 984929 645194 984935
rect 645142 984871 645194 984877
rect 429142 983523 429194 983529
rect 277942 983465 277994 983471
rect 429142 983465 429194 983471
rect 649366 983523 649418 983529
rect 649366 983465 649418 983471
rect 372884 278638 372940 278647
rect 67606 278599 67658 278605
rect 67606 278541 67658 278547
rect 299254 278599 299306 278605
rect 299254 278541 299306 278547
rect 299494 278599 299546 278605
rect 299494 278541 299546 278547
rect 339586 278596 339902 278624
rect 65890 273277 65918 277870
rect 67042 273499 67070 277870
rect 67030 273493 67082 273499
rect 67030 273435 67082 273441
rect 65878 273271 65930 273277
rect 65878 273213 65930 273219
rect 67618 270761 67646 278541
rect 226678 278525 226730 278531
rect 82868 278490 82924 278499
rect 82608 278448 82868 278476
rect 219312 278457 219614 278476
rect 226416 278473 226678 278476
rect 226416 278467 226730 278473
rect 219312 278451 219626 278457
rect 219312 278448 219574 278451
rect 82868 278425 82924 278434
rect 226416 278448 226718 278467
rect 219574 278393 219626 278399
rect 292054 278377 292106 278383
rect 292054 278319 292106 278325
rect 291670 278007 291722 278013
rect 291670 277949 291722 277955
rect 191446 277933 191498 277939
rect 68194 272907 68222 277870
rect 68182 272901 68234 272907
rect 68182 272843 68234 272849
rect 69046 272901 69098 272907
rect 69046 272843 69098 272849
rect 67606 270755 67658 270761
rect 67606 270697 67658 270703
rect 65204 245930 65260 245939
rect 65204 245865 65260 245874
rect 69058 243381 69086 272843
rect 69442 272283 69470 277870
rect 70594 272431 70622 277870
rect 71746 272875 71774 277870
rect 71732 272866 71788 272875
rect 71732 272801 71788 272810
rect 70580 272422 70636 272431
rect 70580 272357 70636 272366
rect 69428 272274 69484 272283
rect 69428 272209 69484 272218
rect 72994 266955 73022 277870
rect 74146 272135 74174 277870
rect 75394 272907 75422 277870
rect 75382 272901 75434 272907
rect 75382 272843 75434 272849
rect 76546 272579 76574 277870
rect 77686 272901 77738 272907
rect 77686 272843 77738 272849
rect 76532 272570 76588 272579
rect 76532 272505 76588 272514
rect 74132 272126 74188 272135
rect 74132 272061 74188 272070
rect 72980 266946 73036 266955
rect 72980 266881 73036 266890
rect 77698 243455 77726 272843
rect 77794 269619 77822 277870
rect 78946 272727 78974 277870
rect 80208 277856 80606 277884
rect 78932 272718 78988 272727
rect 78932 272653 78988 272662
rect 77780 269610 77836 269619
rect 77780 269545 77836 269554
rect 77782 267795 77834 267801
rect 77782 267737 77834 267743
rect 77794 263657 77822 267737
rect 77782 263651 77834 263657
rect 77782 263593 77834 263599
rect 80578 243529 80606 277856
rect 81346 273023 81374 277870
rect 83650 273319 83678 277870
rect 83636 273310 83692 273319
rect 83636 273245 83692 273254
rect 81332 273014 81388 273023
rect 81332 272949 81388 272958
rect 84898 272167 84926 277870
rect 86050 273171 86078 277870
rect 86036 273162 86092 273171
rect 86036 273097 86092 273106
rect 84886 272161 84938 272167
rect 84886 272103 84938 272109
rect 86326 272161 86378 272167
rect 86326 272103 86378 272109
rect 81814 270681 81866 270687
rect 81814 270623 81866 270629
rect 81826 264989 81854 270623
rect 85268 269610 85324 269619
rect 85268 269545 85270 269554
rect 85322 269545 85324 269554
rect 85270 269513 85322 269519
rect 81814 264983 81866 264989
rect 81814 264925 81866 264931
rect 86338 243603 86366 272103
rect 87202 271395 87230 277870
rect 88450 273467 88478 277870
rect 88436 273458 88492 273467
rect 88436 273393 88492 273402
rect 89602 272093 89630 277870
rect 89590 272087 89642 272093
rect 89590 272029 89642 272035
rect 90850 271691 90878 277870
rect 90836 271682 90892 271691
rect 90836 271617 90892 271626
rect 92002 271543 92030 277870
rect 92086 272087 92138 272093
rect 92086 272029 92138 272035
rect 91988 271534 92044 271543
rect 91988 271469 92044 271478
rect 87188 271386 87244 271395
rect 87188 271321 87244 271330
rect 86518 269571 86570 269577
rect 86518 269513 86570 269519
rect 86530 269471 86558 269513
rect 86516 269462 86572 269471
rect 86516 269397 86572 269406
rect 90646 264983 90698 264989
rect 90646 264925 90698 264931
rect 87766 263651 87818 263657
rect 87766 263593 87818 263599
rect 87778 260771 87806 263593
rect 87766 260765 87818 260771
rect 87766 260707 87818 260713
rect 90658 260697 90686 264925
rect 90646 260691 90698 260697
rect 90646 260633 90698 260639
rect 90742 247001 90794 247007
rect 90742 246943 90794 246949
rect 90644 246670 90700 246679
rect 90754 246637 90782 246943
rect 90644 246605 90700 246614
rect 90742 246631 90794 246637
rect 90658 246563 90686 246605
rect 90742 246573 90794 246579
rect 90646 246557 90698 246563
rect 90646 246499 90698 246505
rect 92098 243677 92126 272029
rect 93250 271987 93278 277870
rect 94416 277856 95006 277884
rect 93236 271978 93292 271987
rect 93236 271913 93292 271922
rect 93334 260765 93386 260771
rect 93334 260707 93386 260713
rect 93346 256331 93374 260707
rect 93334 256325 93386 256331
rect 93334 256267 93386 256273
rect 94978 243751 95006 277856
rect 95650 271247 95678 277870
rect 96802 271839 96830 277870
rect 98050 272907 98078 277870
rect 98038 272901 98090 272907
rect 98038 272843 98090 272849
rect 99202 272241 99230 277870
rect 99190 272235 99242 272241
rect 99190 272177 99242 272183
rect 100354 272167 100382 277870
rect 101506 272907 101534 277870
rect 102658 273573 102686 277870
rect 102646 273567 102698 273573
rect 102646 273509 102698 273515
rect 100726 272901 100778 272907
rect 100726 272843 100778 272849
rect 101494 272901 101546 272907
rect 101494 272843 101546 272849
rect 103606 272901 103658 272907
rect 103606 272843 103658 272849
rect 100342 272161 100394 272167
rect 100342 272103 100394 272109
rect 96788 271830 96844 271839
rect 96788 271765 96844 271774
rect 95636 271238 95692 271247
rect 95636 271173 95692 271182
rect 97846 256325 97898 256331
rect 97846 256267 97898 256273
rect 97858 250504 97886 256267
rect 100738 253001 100766 272843
rect 102550 260691 102602 260697
rect 102550 260633 102602 260639
rect 100150 252995 100202 253001
rect 100150 252937 100202 252943
rect 100726 252995 100778 253001
rect 100726 252937 100778 252943
rect 97858 250476 97982 250504
rect 97954 244861 97982 250476
rect 97942 244855 97994 244861
rect 97942 244797 97994 244803
rect 100162 243825 100190 252937
rect 100246 247001 100298 247007
rect 100246 246943 100298 246949
rect 100258 246637 100286 246943
rect 100532 246670 100588 246679
rect 100246 246631 100298 246637
rect 100532 246605 100588 246614
rect 100246 246573 100298 246579
rect 100546 246563 100574 246605
rect 100534 246557 100586 246563
rect 100534 246499 100586 246505
rect 100246 246409 100298 246415
rect 100630 246409 100682 246415
rect 100298 246357 100630 246360
rect 100246 246351 100682 246357
rect 100258 246332 100670 246351
rect 102562 244713 102590 260633
rect 102550 244707 102602 244713
rect 102550 244649 102602 244655
rect 103618 243899 103646 272843
rect 103906 272463 103934 277870
rect 105058 272685 105086 277870
rect 105046 272679 105098 272685
rect 105046 272621 105098 272627
rect 103894 272457 103946 272463
rect 103894 272399 103946 272405
rect 106306 271871 106334 277870
rect 106486 272679 106538 272685
rect 106486 272621 106538 272627
rect 106294 271865 106346 271871
rect 106294 271807 106346 271813
rect 106498 243973 106526 272621
rect 107458 272315 107486 277870
rect 108720 277856 109406 277884
rect 107446 272309 107498 272315
rect 107446 272251 107498 272257
rect 109378 244047 109406 277856
rect 109858 271797 109886 277870
rect 111106 272537 111134 277870
rect 111094 272531 111146 272537
rect 111094 272473 111146 272479
rect 109846 271791 109898 271797
rect 109846 271733 109898 271739
rect 112258 244121 112286 277870
rect 113506 276723 113534 277870
rect 113492 276714 113548 276723
rect 113492 276649 113548 276658
rect 114658 272685 114686 277870
rect 115810 272907 115838 277870
rect 116564 273606 116620 273615
rect 116564 273541 116620 273550
rect 115798 272901 115850 272907
rect 115798 272843 115850 272849
rect 114646 272679 114698 272685
rect 114646 272621 114698 272627
rect 116578 271691 116606 273541
rect 116564 271682 116620 271691
rect 116564 271617 116620 271626
rect 116962 267843 116990 277870
rect 118006 272901 118058 272907
rect 118006 272843 118058 272849
rect 116948 267834 117004 267843
rect 116948 267769 117004 267778
rect 118018 244195 118046 272843
rect 118114 272611 118142 277870
rect 119362 272907 119390 277870
rect 120514 276871 120542 277870
rect 120500 276862 120556 276871
rect 120500 276797 120556 276806
rect 119350 272901 119402 272907
rect 119350 272843 119402 272849
rect 120886 272901 120938 272907
rect 120886 272843 120938 272849
rect 118102 272605 118154 272611
rect 118102 272547 118154 272553
rect 118100 269906 118156 269915
rect 118100 269841 118156 269850
rect 118114 269471 118142 269841
rect 118100 269462 118156 269471
rect 118100 269397 118156 269406
rect 120898 244269 120926 272843
rect 121762 271691 121790 277870
rect 122914 272907 122942 277870
rect 122902 272901 122954 272907
rect 122902 272843 122954 272849
rect 123766 272901 123818 272907
rect 123766 272843 123818 272849
rect 121748 271682 121804 271691
rect 121748 271617 121804 271626
rect 123778 244343 123806 272843
rect 124162 271501 124190 277870
rect 125314 272685 125342 277870
rect 126576 277856 126686 277884
rect 125302 272679 125354 272685
rect 125302 272621 125354 272627
rect 124150 271495 124202 271501
rect 124150 271437 124202 271443
rect 126658 244417 126686 277856
rect 127714 271427 127742 277870
rect 128962 272759 128990 277870
rect 130114 272907 130142 277870
rect 130102 272901 130154 272907
rect 130102 272843 130154 272849
rect 128950 272753 129002 272759
rect 128950 272695 129002 272701
rect 127702 271421 127754 271427
rect 127702 271363 127754 271369
rect 131266 271353 131294 277870
rect 132406 272901 132458 272907
rect 132406 272843 132458 272849
rect 131254 271347 131306 271353
rect 131254 271289 131306 271295
rect 132418 244491 132446 272843
rect 132514 266807 132542 277870
rect 133570 272907 133598 277870
rect 133558 272901 133610 272907
rect 133558 272843 133610 272849
rect 134818 271057 134846 277870
rect 135286 272901 135338 272907
rect 135286 272843 135338 272849
rect 134806 271051 134858 271057
rect 134806 270993 134858 270999
rect 132500 266798 132556 266807
rect 132500 266733 132556 266742
rect 135298 244565 135326 272843
rect 135970 272833 135998 277870
rect 137218 272907 137246 277870
rect 138370 272907 138398 277870
rect 139618 273055 139646 277870
rect 140784 277856 141086 277884
rect 139606 273049 139658 273055
rect 139606 272991 139658 272997
rect 137206 272901 137258 272907
rect 137206 272843 137258 272849
rect 138166 272901 138218 272907
rect 138166 272843 138218 272849
rect 138358 272901 138410 272907
rect 138358 272843 138410 272849
rect 140950 272901 141002 272907
rect 140950 272843 141002 272849
rect 135958 272827 136010 272833
rect 135958 272769 136010 272775
rect 138178 244639 138206 272843
rect 140962 247567 140990 272843
rect 140948 247558 141004 247567
rect 140948 247493 141004 247502
rect 138166 244633 138218 244639
rect 138166 244575 138218 244581
rect 135286 244559 135338 244565
rect 135286 244501 135338 244507
rect 132406 244485 132458 244491
rect 132406 244427 132458 244433
rect 126646 244411 126698 244417
rect 126646 244353 126698 244359
rect 123766 244337 123818 244343
rect 123766 244279 123818 244285
rect 120886 244263 120938 244269
rect 120886 244205 120938 244211
rect 118006 244189 118058 244195
rect 118006 244131 118058 244137
rect 112246 244115 112298 244121
rect 112246 244057 112298 244063
rect 109366 244041 109418 244047
rect 109366 243983 109418 243989
rect 106486 243967 106538 243973
rect 106486 243909 106538 243915
rect 103606 243893 103658 243899
rect 103606 243835 103658 243841
rect 100150 243819 100202 243825
rect 100150 243761 100202 243767
rect 94966 243745 95018 243751
rect 94966 243687 95018 243693
rect 92086 243671 92138 243677
rect 92086 243613 92138 243619
rect 86326 243597 86378 243603
rect 86326 243539 86378 243545
rect 80566 243523 80618 243529
rect 80566 243465 80618 243471
rect 77686 243449 77738 243455
rect 77686 243391 77738 243397
rect 69046 243375 69098 243381
rect 69046 243317 69098 243323
rect 141058 224659 141086 277856
rect 142018 272907 142046 277870
rect 143170 273647 143198 277870
rect 143158 273641 143210 273647
rect 143158 273583 143210 273589
rect 144418 273351 144446 277870
rect 144406 273345 144458 273351
rect 144406 273287 144458 273293
rect 142006 272901 142058 272907
rect 142006 272843 142058 272849
rect 143926 272901 143978 272907
rect 143926 272843 143978 272849
rect 141142 271569 141194 271575
rect 141142 271511 141194 271517
rect 141154 271427 141182 271511
rect 141142 271421 141194 271427
rect 141142 271363 141194 271369
rect 141140 269758 141196 269767
rect 141140 269693 141196 269702
rect 141154 269619 141182 269693
rect 141140 269610 141196 269619
rect 141140 269545 141196 269554
rect 143938 247715 143966 272843
rect 145570 272093 145598 277870
rect 146722 272981 146750 277870
rect 146900 273606 146956 273615
rect 146956 273564 147134 273592
rect 146900 273541 146956 273550
rect 146806 273345 146858 273351
rect 146806 273287 146858 273293
rect 146710 272975 146762 272981
rect 146710 272917 146762 272923
rect 145558 272087 145610 272093
rect 145558 272029 145610 272035
rect 146710 272087 146762 272093
rect 146710 272029 146762 272035
rect 143924 247706 143980 247715
rect 143924 247641 143980 247650
rect 146722 247419 146750 272029
rect 146708 247410 146764 247419
rect 146708 247345 146764 247354
rect 146818 246212 146846 273287
rect 147106 271691 147134 273564
rect 147970 273129 147998 277870
rect 149136 277856 149630 277884
rect 147958 273123 148010 273129
rect 147958 273065 148010 273071
rect 146900 271682 146956 271691
rect 146900 271617 146956 271626
rect 147092 271682 147148 271691
rect 147092 271617 147148 271626
rect 146914 270803 146942 271617
rect 147190 271569 147242 271575
rect 147190 271511 147242 271517
rect 147202 271279 147230 271511
rect 147190 271273 147242 271279
rect 147190 271215 147242 271221
rect 146900 270794 146956 270803
rect 146900 270729 146956 270738
rect 149602 247123 149630 277856
rect 149686 273123 149738 273129
rect 149686 273065 149738 273071
rect 149588 247114 149644 247123
rect 149588 247049 149644 247058
rect 146626 246184 146846 246212
rect 144598 244781 144650 244787
rect 144598 244723 144650 244729
rect 142966 244707 143018 244713
rect 142966 244649 143018 244655
rect 141142 242265 141194 242271
rect 141142 242207 141194 242213
rect 141154 241975 141182 242207
rect 141142 241969 141194 241975
rect 141142 241911 141194 241917
rect 142978 239015 143006 244649
rect 144610 240495 144638 244723
rect 146324 240602 146380 240611
rect 146324 240537 146380 240546
rect 144598 240489 144650 240495
rect 144598 240431 144650 240437
rect 142966 239009 143018 239015
rect 142966 238951 143018 238957
rect 145556 236902 145612 236911
rect 145556 236837 145612 236846
rect 145570 236203 145598 236837
rect 145558 236197 145610 236203
rect 145558 236139 145610 236145
rect 146134 235235 146186 235241
rect 146134 235177 146186 235183
rect 144404 232166 144460 232175
rect 144404 232101 144460 232110
rect 144418 230505 144446 232101
rect 144406 230499 144458 230505
rect 144406 230441 144458 230447
rect 144020 226690 144076 226699
rect 144020 226625 144076 226634
rect 144034 226435 144062 226625
rect 144022 226429 144074 226435
rect 144022 226371 144074 226377
rect 144020 225062 144076 225071
rect 144020 224997 144076 225006
rect 144034 224733 144062 224997
rect 144022 224727 144074 224733
rect 144022 224669 144074 224675
rect 141046 224653 141098 224659
rect 141046 224595 141098 224601
rect 144116 223730 144172 223739
rect 144116 223665 144172 223674
rect 144020 222990 144076 222999
rect 144020 222925 144076 222934
rect 144034 221921 144062 222925
rect 144022 221915 144074 221921
rect 144022 221857 144074 221863
rect 144130 221847 144158 223665
rect 144118 221841 144170 221847
rect 144118 221783 144170 221789
rect 146146 221773 146174 235177
rect 146338 227545 146366 240537
rect 146422 236197 146474 236203
rect 146422 236139 146474 236145
rect 146434 235241 146462 236139
rect 146422 235235 146474 235241
rect 146422 235177 146474 235183
rect 146420 235126 146476 235135
rect 146420 235061 146476 235070
rect 146326 227539 146378 227545
rect 146326 227481 146378 227487
rect 146134 221767 146186 221773
rect 146134 221709 146186 221715
rect 146230 221767 146282 221773
rect 146230 221709 146282 221715
rect 144020 220178 144076 220187
rect 144020 220113 144076 220122
rect 144034 218961 144062 220113
rect 145364 218994 145420 219003
rect 144022 218955 144074 218961
rect 145364 218929 145420 218938
rect 144022 218897 144074 218903
rect 144020 218254 144076 218263
rect 144020 218189 144076 218198
rect 144034 216075 144062 218189
rect 144022 216069 144074 216075
rect 144022 216011 144074 216017
rect 144116 215294 144172 215303
rect 144116 215229 144172 215238
rect 144020 214554 144076 214563
rect 144020 214489 144076 214498
rect 144034 213189 144062 214489
rect 144130 213263 144158 215229
rect 144118 213257 144170 213263
rect 144118 213199 144170 213205
rect 144022 213183 144074 213189
rect 144022 213125 144074 213131
rect 144116 209818 144172 209827
rect 144116 209753 144172 209762
rect 144022 207485 144074 207491
rect 144020 207450 144022 207459
rect 144074 207450 144076 207459
rect 144130 207417 144158 209753
rect 144020 207385 144076 207394
rect 144118 207411 144170 207417
rect 144118 207353 144170 207359
rect 144020 205674 144076 205683
rect 144020 205609 144076 205618
rect 144034 204531 144062 205609
rect 144022 204525 144074 204531
rect 144022 204467 144074 204473
rect 144020 203454 144076 203463
rect 144020 203389 144076 203398
rect 144034 201645 144062 203389
rect 144596 202122 144652 202131
rect 144596 202057 144652 202066
rect 144022 201639 144074 201645
rect 144022 201581 144074 201587
rect 144116 201382 144172 201391
rect 144116 201317 144172 201326
rect 144020 199014 144076 199023
rect 144020 198949 144076 198958
rect 144034 198833 144062 198949
rect 144130 198907 144158 201317
rect 144118 198901 144170 198907
rect 144118 198843 144170 198849
rect 144022 198827 144074 198833
rect 144022 198769 144074 198775
rect 144020 197830 144076 197839
rect 144020 197765 144076 197774
rect 144034 195873 144062 197765
rect 144404 196646 144460 196655
rect 144404 196581 144460 196590
rect 144022 195867 144074 195873
rect 144022 195809 144074 195815
rect 144308 194870 144364 194879
rect 144308 194805 144364 194814
rect 50422 194535 50474 194541
rect 50422 194477 50474 194483
rect 144020 192946 144076 192955
rect 144020 192881 144076 192890
rect 43126 192241 43178 192247
rect 43126 192183 43178 192189
rect 144034 190175 144062 192881
rect 144022 190169 144074 190175
rect 144022 190111 144074 190117
rect 42934 187283 42986 187289
rect 42934 187225 42986 187231
rect 42602 187095 42686 187123
rect 42550 187077 42602 187083
rect 42370 184764 42494 184792
rect 41780 184214 41836 184223
rect 41780 184149 41836 184158
rect 41794 183742 41822 184149
rect 41780 183622 41836 183631
rect 41780 183557 41836 183566
rect 41794 183121 41822 183557
rect 41780 182882 41836 182891
rect 41780 182817 41836 182826
rect 41794 182484 41822 182817
rect 42466 125351 42494 184764
rect 144022 175665 144074 175671
rect 144022 175607 144074 175613
rect 144034 166717 144062 175607
rect 144022 166711 144074 166717
rect 144022 166653 144074 166659
rect 144020 166602 144076 166611
rect 144020 166537 144076 166546
rect 144034 164201 144062 166537
rect 144022 164195 144074 164201
rect 144022 164137 144074 164143
rect 144020 162902 144076 162911
rect 144020 162837 144076 162846
rect 144034 161315 144062 162837
rect 144022 161309 144074 161315
rect 144022 161251 144074 161257
rect 144116 159942 144172 159951
rect 144116 159877 144172 159886
rect 144020 159350 144076 159359
rect 144020 159285 144076 159294
rect 144034 158503 144062 159285
rect 144022 158497 144074 158503
rect 144022 158439 144074 158445
rect 144130 156524 144158 159877
rect 144212 158166 144268 158175
rect 144212 158101 144268 158110
rect 144034 156496 144158 156524
rect 144034 155932 144062 156496
rect 144116 156390 144172 156399
rect 144116 156325 144172 156334
rect 143938 155904 144062 155932
rect 143938 155636 143966 155904
rect 144020 155798 144076 155807
rect 144020 155733 144022 155742
rect 144074 155733 144076 155742
rect 144022 155701 144074 155707
rect 144130 155691 144158 156325
rect 144118 155685 144170 155691
rect 143938 155608 144062 155636
rect 144118 155627 144170 155633
rect 144226 155617 144254 158101
rect 144034 154600 144062 155608
rect 144214 155611 144266 155617
rect 144214 155553 144266 155559
rect 144034 154572 144254 154600
rect 144116 154466 144172 154475
rect 144116 154401 144172 154410
rect 144020 152986 144076 152995
rect 144020 152921 144076 152930
rect 144034 152805 144062 152921
rect 144022 152799 144074 152805
rect 144022 152741 144074 152747
rect 144130 152731 144158 154401
rect 144118 152725 144170 152731
rect 144118 152667 144170 152673
rect 144116 151654 144172 151663
rect 144116 151589 144172 151598
rect 144020 150914 144076 150923
rect 144020 150849 144076 150858
rect 144034 149845 144062 150849
rect 144130 149919 144158 151589
rect 144118 149913 144170 149919
rect 144118 149855 144170 149861
rect 144022 149839 144074 149845
rect 144022 149781 144074 149787
rect 144022 149691 144074 149697
rect 144022 149633 144074 149639
rect 144034 147181 144062 149633
rect 144226 147200 144254 154572
rect 144022 147175 144074 147181
rect 144022 147117 144074 147123
rect 144130 147172 144254 147200
rect 144130 147052 144158 147172
rect 144034 147024 144158 147052
rect 144212 147066 144268 147075
rect 143924 141294 143980 141303
rect 143924 141229 143980 141238
rect 143828 138334 143884 138343
rect 143828 138269 143830 138278
rect 143882 138269 143884 138278
rect 143830 138237 143882 138243
rect 143938 138227 143966 141229
rect 143926 138221 143978 138227
rect 143926 138163 143978 138169
rect 143926 130155 143978 130161
rect 143926 130097 143978 130103
rect 143938 126757 143966 130097
rect 143926 126751 143978 126757
rect 143926 126693 143978 126699
rect 39862 125345 39914 125351
rect 39860 125310 39862 125319
rect 42454 125345 42506 125351
rect 39914 125310 39916 125319
rect 42454 125287 42506 125293
rect 39860 125245 39916 125254
rect 143830 115207 143882 115213
rect 143830 115149 143882 115155
rect 143734 115133 143786 115139
rect 143734 115075 143786 115081
rect 143746 103373 143774 115075
rect 143842 106555 143870 115149
rect 143830 106549 143882 106555
rect 143830 106491 143882 106497
rect 144034 104927 144062 147024
rect 144212 147001 144268 147010
rect 144118 146953 144170 146959
rect 144118 146895 144170 146901
rect 144130 115139 144158 146895
rect 144226 146145 144254 147001
rect 144214 146139 144266 146145
rect 144214 146081 144266 146087
rect 144212 146030 144268 146039
rect 144212 145965 144268 145974
rect 144226 144369 144254 145965
rect 144214 144363 144266 144369
rect 144214 144305 144266 144311
rect 144212 144254 144268 144263
rect 144212 144189 144268 144198
rect 144226 144073 144254 144189
rect 144214 144067 144266 144073
rect 144214 144009 144266 144015
rect 144212 143218 144268 143227
rect 144212 143153 144268 143162
rect 144226 142593 144254 143153
rect 144214 142587 144266 142593
rect 144214 142529 144266 142535
rect 144212 142478 144268 142487
rect 144212 142413 144268 142422
rect 144226 141187 144254 142413
rect 144214 141181 144266 141187
rect 144214 141123 144266 141129
rect 144214 140885 144266 140891
rect 144214 140827 144266 140833
rect 144226 134897 144254 140827
rect 144214 134891 144266 134897
rect 144214 134833 144266 134839
rect 144212 134782 144268 134791
rect 144212 134717 144268 134726
rect 144226 134231 144254 134717
rect 144214 134225 144266 134231
rect 144214 134167 144266 134173
rect 144212 134042 144268 134051
rect 144212 133977 144268 133986
rect 144226 132751 144254 133977
rect 144214 132745 144266 132751
rect 144214 132687 144266 132693
rect 144214 132597 144266 132603
rect 144214 132539 144266 132545
rect 144226 130161 144254 132539
rect 144214 130155 144266 130161
rect 144214 130097 144266 130103
rect 144212 130046 144268 130055
rect 144212 129981 144268 129990
rect 144226 129643 144254 129981
rect 144214 129637 144266 129643
rect 144214 129579 144266 129585
rect 144214 126751 144266 126757
rect 144214 126693 144266 126699
rect 144118 115133 144170 115139
rect 144118 115075 144170 115081
rect 144118 114985 144170 114991
rect 144118 114927 144170 114933
rect 144022 104921 144074 104927
rect 144022 104863 144074 104869
rect 144130 104835 144158 114927
rect 144034 104807 144158 104835
rect 144034 104428 144062 104807
rect 144116 104738 144172 104747
rect 144116 104673 144172 104682
rect 143938 104400 144062 104428
rect 143938 103984 143966 104400
rect 143938 103956 144062 103984
rect 143734 103367 143786 103373
rect 143734 103309 143786 103315
rect 144034 101764 144062 103956
rect 144130 103743 144158 104673
rect 144118 103737 144170 103743
rect 144118 103679 144170 103685
rect 144116 102814 144172 102823
rect 144116 102749 144172 102758
rect 143938 101736 144062 101764
rect 143938 101468 143966 101736
rect 144020 101630 144076 101639
rect 144020 101565 144022 101574
rect 144074 101565 144076 101574
rect 144022 101533 144074 101539
rect 143938 101440 144062 101468
rect 144034 100709 144062 101440
rect 144130 100857 144158 102749
rect 144118 100851 144170 100857
rect 144118 100793 144170 100799
rect 144022 100703 144074 100709
rect 144022 100645 144074 100651
rect 143926 100037 143978 100043
rect 143926 99979 143978 99985
rect 143938 80729 143966 99979
rect 144116 99114 144172 99123
rect 144116 99049 144172 99058
rect 144022 98113 144074 98119
rect 144020 98078 144022 98087
rect 144074 98078 144076 98087
rect 144130 98045 144158 99049
rect 144020 98013 144076 98022
rect 144118 98039 144170 98045
rect 144118 97981 144170 97987
rect 144116 96302 144172 96311
rect 144116 96237 144172 96246
rect 144020 95562 144076 95571
rect 144020 95497 144076 95506
rect 144034 95159 144062 95497
rect 144022 95153 144074 95159
rect 144022 95095 144074 95101
rect 144130 95085 144158 96237
rect 144118 95079 144170 95085
rect 144118 95021 144170 95027
rect 144116 94378 144172 94387
rect 144116 94313 144172 94322
rect 144020 92750 144076 92759
rect 144020 92685 144076 92694
rect 144034 92199 144062 92685
rect 144130 92273 144158 94313
rect 144118 92267 144170 92273
rect 144118 92209 144170 92215
rect 144022 92193 144074 92199
rect 144022 92135 144074 92141
rect 144116 91418 144172 91427
rect 144116 91353 144172 91362
rect 144020 89642 144076 89651
rect 144020 89577 144076 89586
rect 144034 89461 144062 89577
rect 144022 89455 144074 89461
rect 144022 89397 144074 89403
rect 144130 89313 144158 91353
rect 144118 89307 144170 89313
rect 144118 89249 144170 89255
rect 144116 87866 144172 87875
rect 144116 87801 144172 87810
rect 143926 80723 143978 80729
rect 143926 80665 143978 80671
rect 144020 75138 144076 75147
rect 144020 75073 144076 75082
rect 144034 75031 144062 75073
rect 144022 75025 144074 75031
rect 144130 74999 144158 87801
rect 144022 74967 144074 74973
rect 144116 74990 144172 74999
rect 144116 74925 144172 74934
rect 144118 74137 144170 74143
rect 144118 74079 144170 74085
rect 144130 72779 144158 74079
rect 144116 72770 144172 72779
rect 144116 72705 144172 72714
rect 144020 70994 144076 71003
rect 144020 70929 144076 70938
rect 144034 70295 144062 70929
rect 144022 70289 144074 70295
rect 144022 70231 144074 70237
rect 144020 69810 144076 69819
rect 144020 69745 144076 69754
rect 144034 69185 144062 69745
rect 144022 69179 144074 69185
rect 144022 69121 144074 69127
rect 144116 67442 144172 67451
rect 144116 67377 144172 67386
rect 144130 67261 144158 67377
rect 144118 67255 144170 67261
rect 144118 67197 144170 67203
rect 144022 66219 144074 66225
rect 144022 66161 144074 66167
rect 144034 62969 144062 66161
rect 144118 65035 144170 65041
rect 144118 64977 144170 64983
rect 144022 62963 144074 62969
rect 144022 62905 144074 62911
rect 144020 62854 144076 62863
rect 144020 62789 144076 62798
rect 144034 62525 144062 62789
rect 144022 62519 144074 62525
rect 144022 62461 144074 62467
rect 144022 59633 144074 59639
rect 144020 59598 144022 59607
rect 144074 59598 144076 59607
rect 144020 59533 144076 59542
rect 144022 59041 144074 59047
rect 144022 58983 144074 58989
rect 144034 58719 144062 58983
rect 144020 58710 144076 58719
rect 144020 58645 144076 58654
rect 144022 57117 144074 57123
rect 144020 57082 144022 57091
rect 144074 57082 144076 57091
rect 144020 57017 144076 57026
rect 144022 56525 144074 56531
rect 144022 56467 144074 56473
rect 144034 56203 144062 56467
rect 144020 56194 144076 56203
rect 144020 56129 144076 56138
rect 144020 54714 144076 54723
rect 144020 54649 144022 54658
rect 144074 54649 144076 54658
rect 144022 54617 144074 54623
rect 144022 54157 144074 54163
rect 144022 54099 144074 54105
rect 144034 53835 144062 54099
rect 144020 53826 144076 53835
rect 144020 53761 144076 53770
rect 137494 52307 137546 52313
rect 137494 52249 137546 52255
rect 137506 51888 137534 52249
rect 137280 51860 137534 51888
rect 144130 50019 144158 64977
rect 144226 50241 144254 126693
rect 144322 115213 144350 194805
rect 144418 115213 144446 196581
rect 144500 185250 144556 185259
rect 144500 185185 144556 185194
rect 144514 184477 144542 185185
rect 144502 184471 144554 184477
rect 144502 184413 144554 184419
rect 144500 164826 144556 164835
rect 144500 164761 144556 164770
rect 144514 149697 144542 164761
rect 144502 149691 144554 149697
rect 144502 149633 144554 149639
rect 144500 147954 144556 147963
rect 144500 147889 144556 147898
rect 144514 146959 144542 147889
rect 144502 146953 144554 146959
rect 144502 146895 144554 146901
rect 144502 146287 144554 146293
rect 144502 146229 144554 146235
rect 144514 140891 144542 146229
rect 144502 140885 144554 140891
rect 144502 140827 144554 140833
rect 144500 139518 144556 139527
rect 144500 139453 144556 139462
rect 144514 138375 144542 139453
rect 144502 138369 144554 138375
rect 144502 138311 144554 138317
rect 144502 138221 144554 138227
rect 144502 138163 144554 138169
rect 144514 132973 144542 138163
rect 144502 132967 144554 132973
rect 144502 132909 144554 132915
rect 144500 132858 144556 132867
rect 144500 132793 144556 132802
rect 144514 132603 144542 132793
rect 144502 132597 144554 132603
rect 144502 132539 144554 132545
rect 144500 131082 144556 131091
rect 144500 131017 144556 131026
rect 144514 129717 144542 131017
rect 144502 129711 144554 129717
rect 144502 129653 144554 129659
rect 144502 129563 144554 129569
rect 144502 129505 144554 129511
rect 144514 115213 144542 129505
rect 144310 115207 144362 115213
rect 144310 115149 144362 115155
rect 144406 115207 144458 115213
rect 144406 115149 144458 115155
rect 144502 115207 144554 115213
rect 144502 115149 144554 115155
rect 144610 115107 144638 202057
rect 144692 180514 144748 180523
rect 144692 180449 144748 180458
rect 144706 163757 144734 180449
rect 145268 179774 145324 179783
rect 145268 179709 145324 179718
rect 145282 178705 145310 179709
rect 145270 178699 145322 178705
rect 145270 178641 145322 178647
rect 145268 176074 145324 176083
rect 145268 176009 145324 176018
rect 145172 174446 145228 174455
rect 145172 174381 145228 174390
rect 144884 172078 144940 172087
rect 144884 172013 144940 172022
rect 144694 163751 144746 163757
rect 144694 163693 144746 163699
rect 144692 163642 144748 163651
rect 144692 163577 144748 163586
rect 144706 147255 144734 163577
rect 144788 161422 144844 161431
rect 144788 161357 144844 161366
rect 144694 147249 144746 147255
rect 144694 147191 144746 147197
rect 144694 147101 144746 147107
rect 144694 147043 144746 147049
rect 144706 136969 144734 147043
rect 144694 136963 144746 136969
rect 144694 136905 144746 136911
rect 144802 136840 144830 161357
rect 144706 136812 144830 136840
rect 144308 115098 144364 115107
rect 144308 115033 144364 115042
rect 144596 115098 144652 115107
rect 144596 115033 144652 115042
rect 144322 106056 144350 115033
rect 144502 114985 144554 114991
rect 144502 114927 144554 114933
rect 144598 114985 144650 114991
rect 144598 114927 144650 114933
rect 144404 113174 144460 113183
rect 144404 113109 144460 113118
rect 144418 112475 144446 113109
rect 144406 112469 144458 112475
rect 144406 112411 144458 112417
rect 144404 111250 144460 111259
rect 144404 111185 144460 111194
rect 144418 109589 144446 111185
rect 144406 109583 144458 109589
rect 144406 109525 144458 109531
rect 144404 108290 144460 108299
rect 144404 108225 144460 108234
rect 144418 106703 144446 108225
rect 144406 106697 144458 106703
rect 144406 106639 144458 106645
rect 144322 106028 144446 106056
rect 144308 105922 144364 105931
rect 144308 105857 144364 105866
rect 144322 103817 144350 105857
rect 144310 103811 144362 103817
rect 144310 103753 144362 103759
rect 144308 103702 144364 103711
rect 144308 103637 144364 103646
rect 144322 100043 144350 103637
rect 144418 100635 144446 106028
rect 144406 100629 144458 100635
rect 144406 100571 144458 100577
rect 144310 100037 144362 100043
rect 144310 99979 144362 99985
rect 144308 99854 144364 99863
rect 144308 99789 144364 99798
rect 144322 97971 144350 99789
rect 144310 97965 144362 97971
rect 144310 97907 144362 97913
rect 144308 90826 144364 90835
rect 144308 90761 144364 90770
rect 144322 89387 144350 90761
rect 144310 89381 144362 89387
rect 144310 89323 144362 89329
rect 144514 86501 144542 114927
rect 144610 103521 144638 114927
rect 144706 106523 144734 136812
rect 144790 136741 144842 136747
rect 144790 136683 144842 136689
rect 144692 106514 144748 106523
rect 144692 106449 144748 106458
rect 144802 106352 144830 136683
rect 144706 106324 144830 106352
rect 144598 103515 144650 103521
rect 144598 103457 144650 103463
rect 144598 103367 144650 103373
rect 144598 103309 144650 103315
rect 144610 94937 144638 103309
rect 144598 94931 144650 94937
rect 144598 94873 144650 94879
rect 144706 86520 144734 106324
rect 144790 104255 144842 104261
rect 144790 104197 144842 104203
rect 144802 104007 144830 104197
rect 144788 103998 144844 104007
rect 144788 103933 144844 103942
rect 144502 86495 144554 86501
rect 144706 86492 144830 86520
rect 144502 86437 144554 86443
rect 144502 86347 144554 86353
rect 144502 86289 144554 86295
rect 144404 80762 144460 80771
rect 144404 80697 144460 80706
rect 144308 78690 144364 78699
rect 144308 78625 144364 78634
rect 144322 77917 144350 78625
rect 144310 77911 144362 77917
rect 144310 77853 144362 77859
rect 144308 77506 144364 77515
rect 144308 77441 144364 77450
rect 144322 74957 144350 77441
rect 144310 74951 144362 74957
rect 144310 74893 144362 74899
rect 144310 74211 144362 74217
rect 144310 74153 144362 74159
rect 144322 65041 144350 74153
rect 144310 65035 144362 65041
rect 144310 64977 144362 64983
rect 144310 64887 144362 64893
rect 144310 64829 144362 64835
rect 144322 64639 144350 64829
rect 144308 64630 144364 64639
rect 144308 64565 144364 64574
rect 144310 62963 144362 62969
rect 144310 62905 144362 62911
rect 144322 51351 144350 62905
rect 144418 52091 144446 80697
rect 144406 52085 144458 52091
rect 144406 52027 144458 52033
rect 144310 51345 144362 51351
rect 144310 51287 144362 51293
rect 144514 50389 144542 86289
rect 144596 83574 144652 83583
rect 144596 83509 144652 83518
rect 144610 52017 144638 83509
rect 144694 80723 144746 80729
rect 144694 80665 144746 80671
rect 144706 66225 144734 80665
rect 144802 66267 144830 86492
rect 144788 66258 144844 66267
rect 144694 66219 144746 66225
rect 144788 66193 144844 66202
rect 144694 66161 144746 66167
rect 144598 52011 144650 52017
rect 144598 51953 144650 51959
rect 144898 50759 144926 172013
rect 145076 170154 145132 170163
rect 145076 170089 145132 170098
rect 144980 168378 145036 168387
rect 144980 168313 145036 168322
rect 144994 65652 145022 168313
rect 145090 65781 145118 170089
rect 145078 65775 145130 65781
rect 145078 65717 145130 65723
rect 144994 65624 145118 65652
rect 144980 65518 145036 65527
rect 144980 65453 145036 65462
rect 144994 64819 145022 65453
rect 144982 64813 145034 64819
rect 144982 64755 145034 64761
rect 144980 64630 145036 64639
rect 144980 64565 145036 64574
rect 144886 50753 144938 50759
rect 144886 50695 144938 50701
rect 144502 50383 144554 50389
rect 144502 50325 144554 50331
rect 144214 50235 144266 50241
rect 144214 50177 144266 50183
rect 144994 50167 145022 64565
rect 145090 50685 145118 65624
rect 145078 50679 145130 50685
rect 145078 50621 145130 50627
rect 145186 50537 145214 174381
rect 145282 50611 145310 176009
rect 145378 51573 145406 218929
rect 145460 216478 145516 216487
rect 145460 216413 145516 216422
rect 145474 74217 145502 216413
rect 145556 211742 145612 211751
rect 145556 211677 145612 211686
rect 145462 74211 145514 74217
rect 145462 74153 145514 74159
rect 145462 74063 145514 74069
rect 145462 74005 145514 74011
rect 145474 65929 145502 74005
rect 145462 65923 145514 65929
rect 145462 65865 145514 65871
rect 145462 65775 145514 65781
rect 145462 65717 145514 65723
rect 145366 51567 145418 51573
rect 145366 51509 145418 51515
rect 145270 50605 145322 50611
rect 145270 50547 145322 50553
rect 145174 50531 145226 50537
rect 145174 50473 145226 50479
rect 145474 50463 145502 65717
rect 145570 51499 145598 211677
rect 146242 211635 146270 221709
rect 146434 213485 146462 235061
rect 146518 227539 146570 227545
rect 146518 227481 146570 227487
rect 146530 217777 146558 227481
rect 146626 224585 146654 246184
rect 146708 238678 146764 238687
rect 146708 238613 146764 238622
rect 146722 236203 146750 238613
rect 148342 237603 148394 237609
rect 148342 237545 148394 237551
rect 146804 236310 146860 236319
rect 146804 236245 146806 236254
rect 146858 236245 146860 236254
rect 146806 236213 146858 236219
rect 146710 236197 146762 236203
rect 146710 236139 146762 236145
rect 146804 233646 146860 233655
rect 146804 233581 146860 233590
rect 146818 233317 146846 233581
rect 146806 233311 146858 233317
rect 146806 233253 146858 233259
rect 146804 231426 146860 231435
rect 146804 231361 146860 231370
rect 146818 230579 146846 231361
rect 146806 230573 146858 230579
rect 146806 230515 146858 230521
rect 146708 230242 146764 230251
rect 146708 230177 146764 230186
rect 146722 227693 146750 230177
rect 146804 229058 146860 229067
rect 146804 228993 146860 229002
rect 146818 228803 146846 228993
rect 146806 228797 146858 228803
rect 146806 228739 146858 228745
rect 146804 227726 146860 227735
rect 146710 227687 146762 227693
rect 146804 227661 146860 227670
rect 146710 227629 146762 227635
rect 146818 227619 146846 227661
rect 146806 227613 146858 227619
rect 146806 227555 146858 227561
rect 146614 224579 146666 224585
rect 146614 224521 146666 224527
rect 146518 217771 146570 217777
rect 146518 217713 146570 217719
rect 146518 217623 146570 217629
rect 146518 217565 146570 217571
rect 146422 213479 146474 213485
rect 146422 213421 146474 213427
rect 146420 213370 146476 213379
rect 146420 213305 146422 213314
rect 146474 213305 146476 213314
rect 146422 213273 146474 213279
rect 146530 211728 146558 217565
rect 146710 213479 146762 213485
rect 146710 213421 146762 213427
rect 146434 211700 146558 211728
rect 146230 211629 146282 211635
rect 146230 211571 146282 211577
rect 145748 210558 145804 210567
rect 145748 210493 145804 210502
rect 145652 208042 145708 208051
rect 145652 207977 145708 207986
rect 145558 51493 145610 51499
rect 145558 51435 145610 51441
rect 145666 51277 145694 207977
rect 145654 51271 145706 51277
rect 145654 51213 145706 51219
rect 145762 51203 145790 210493
rect 145844 205082 145900 205091
rect 145844 205017 145900 205026
rect 145750 51197 145802 51203
rect 145750 51139 145802 51145
rect 145462 50457 145514 50463
rect 145462 50399 145514 50405
rect 144982 50161 145034 50167
rect 144982 50103 145034 50109
rect 145858 50093 145886 205017
rect 146228 199606 146284 199615
rect 146228 199541 146284 199550
rect 146242 198759 146270 199541
rect 146230 198753 146282 198759
rect 146230 198695 146282 198701
rect 146434 197224 146462 211700
rect 146518 211629 146570 211635
rect 146518 211571 146570 211577
rect 146338 197196 146462 197224
rect 145940 193686 145996 193695
rect 145940 193621 145996 193630
rect 145954 51425 145982 193621
rect 146036 191762 146092 191771
rect 146036 191697 146092 191706
rect 146050 74069 146078 191697
rect 146228 190134 146284 190143
rect 146228 190069 146284 190078
rect 146132 189394 146188 189403
rect 146132 189329 146188 189338
rect 146038 74063 146090 74069
rect 146038 74005 146090 74011
rect 146036 73954 146092 73963
rect 146036 73889 146092 73898
rect 146050 72071 146078 73889
rect 146038 72065 146090 72071
rect 146038 72007 146090 72013
rect 146038 69253 146090 69259
rect 146038 69195 146090 69201
rect 145942 51419 145994 51425
rect 145942 51361 145994 51367
rect 146050 50315 146078 69195
rect 146146 51129 146174 189329
rect 146134 51123 146186 51129
rect 146134 51065 146186 51071
rect 146242 51055 146270 190069
rect 146338 146293 146366 197196
rect 146420 188210 146476 188219
rect 146420 188145 146476 188154
rect 146434 187289 146462 188145
rect 146422 187283 146474 187289
rect 146422 187225 146474 187231
rect 146420 186434 146476 186443
rect 146420 186369 146476 186378
rect 146326 146287 146378 146293
rect 146326 146229 146378 146235
rect 146326 146139 146378 146145
rect 146326 146081 146378 146087
rect 146338 129569 146366 146081
rect 146326 129563 146378 129569
rect 146326 129505 146378 129511
rect 146324 127530 146380 127539
rect 146324 127465 146380 127474
rect 146338 126757 146366 127465
rect 146326 126751 146378 126757
rect 146326 126693 146378 126699
rect 146324 125162 146380 125171
rect 146324 125097 146380 125106
rect 146338 123945 146366 125097
rect 146326 123939 146378 123945
rect 146326 123881 146378 123887
rect 146326 123791 146378 123797
rect 146326 123733 146378 123739
rect 146338 119209 146366 123733
rect 146326 119203 146378 119209
rect 146326 119145 146378 119151
rect 146324 119094 146380 119103
rect 146324 119029 146380 119038
rect 146338 118173 146366 119029
rect 146326 118167 146378 118173
rect 146326 118109 146378 118115
rect 146326 118019 146378 118025
rect 146326 117961 146378 117967
rect 146338 115213 146366 117961
rect 146326 115207 146378 115213
rect 146326 115149 146378 115155
rect 146326 115059 146378 115065
rect 146326 115001 146378 115007
rect 146338 103595 146366 115001
rect 146326 103589 146378 103595
rect 146326 103531 146378 103537
rect 146324 84166 146380 84175
rect 146324 84101 146380 84110
rect 146338 69259 146366 84101
rect 146326 69253 146378 69259
rect 146326 69195 146378 69201
rect 146324 69070 146380 69079
rect 146324 69005 146380 69014
rect 146338 66447 146366 69005
rect 146326 66441 146378 66447
rect 146326 66383 146378 66389
rect 146326 65923 146378 65929
rect 146326 65865 146378 65871
rect 146230 51049 146282 51055
rect 146230 50991 146282 50997
rect 146038 50309 146090 50315
rect 146038 50251 146090 50257
rect 145846 50087 145898 50093
rect 145846 50029 145898 50035
rect 144118 50013 144170 50019
rect 144118 49955 144170 49961
rect 146338 49945 146366 65865
rect 146434 50981 146462 186369
rect 146530 175671 146558 211571
rect 146612 183326 146668 183335
rect 146612 183261 146668 183270
rect 146518 175665 146570 175671
rect 146518 175607 146570 175613
rect 146518 166711 146570 166717
rect 146518 166653 146570 166659
rect 146530 126799 146558 166653
rect 146516 126790 146572 126799
rect 146516 126725 146572 126734
rect 146516 115246 146572 115255
rect 146516 115181 146572 115190
rect 146530 104853 146558 115181
rect 146518 104847 146570 104853
rect 146518 104789 146570 104795
rect 146518 104699 146570 104705
rect 146518 104641 146570 104647
rect 146530 95011 146558 104641
rect 146518 95005 146570 95011
rect 146518 94947 146570 94953
rect 146516 87126 146572 87135
rect 146516 87061 146572 87070
rect 146530 77640 146558 87061
rect 146626 77769 146654 183261
rect 146722 134601 146750 213421
rect 148246 213183 148298 213189
rect 148246 213125 148298 213131
rect 146804 184510 146860 184519
rect 146804 184445 146860 184454
rect 146818 184403 146846 184445
rect 146806 184397 146858 184403
rect 146806 184339 146858 184345
rect 146804 181846 146860 181855
rect 146804 181781 146860 181790
rect 146818 181517 146846 181781
rect 146806 181511 146858 181517
rect 146806 181453 146858 181459
rect 146806 178625 146858 178631
rect 146804 178590 146806 178599
rect 146858 178590 146860 178599
rect 146804 178525 146860 178534
rect 146804 176814 146860 176823
rect 146804 176749 146860 176758
rect 146818 175745 146846 176749
rect 146806 175739 146858 175745
rect 146806 175681 146858 175687
rect 146804 173410 146860 173419
rect 146804 173345 146860 173354
rect 146818 172859 146846 173345
rect 146806 172853 146858 172859
rect 146806 172795 146858 172801
rect 146804 171338 146860 171347
rect 146804 171273 146806 171282
rect 146858 171273 146860 171282
rect 146806 171241 146858 171247
rect 146804 167638 146860 167647
rect 146804 167573 146860 167582
rect 146818 167309 146846 167573
rect 146806 167303 146858 167309
rect 146806 167245 146858 167251
rect 146806 163751 146858 163757
rect 146806 163693 146858 163699
rect 146818 155932 146846 163693
rect 146818 155904 146942 155932
rect 146914 155636 146942 155904
rect 146818 155608 146942 155636
rect 146710 134595 146762 134601
rect 146710 134537 146762 134543
rect 146818 134495 146846 155608
rect 146900 137594 146956 137603
rect 146900 137529 146956 137538
rect 146914 136303 146942 137529
rect 146902 136297 146954 136303
rect 146902 136239 146954 136245
rect 146900 136114 146956 136123
rect 146900 136049 146956 136058
rect 146914 136007 146942 136049
rect 146902 136001 146954 136007
rect 146902 135943 146954 135949
rect 146998 134891 147050 134897
rect 146998 134833 147050 134839
rect 146804 134486 146860 134495
rect 146804 134421 146860 134430
rect 146806 134373 146858 134379
rect 146858 134321 146942 134324
rect 146806 134315 146942 134321
rect 146818 134296 146942 134315
rect 146806 134225 146858 134231
rect 146806 134167 146858 134173
rect 146818 132677 146846 134167
rect 146806 132671 146858 132677
rect 146806 132613 146858 132619
rect 146804 132562 146860 132571
rect 146804 132497 146860 132506
rect 146708 129306 146764 129315
rect 146708 129241 146764 129250
rect 146722 126831 146750 129241
rect 146710 126825 146762 126831
rect 146710 126767 146762 126773
rect 146708 124422 146764 124431
rect 146708 124357 146764 124366
rect 146722 124093 146750 124357
rect 146710 124087 146762 124093
rect 146710 124029 146762 124035
rect 146708 122646 146764 122655
rect 146708 122581 146764 122590
rect 146722 121059 146750 122581
rect 146710 121053 146762 121059
rect 146710 120995 146762 121001
rect 146708 120870 146764 120879
rect 146708 120805 146764 120814
rect 146722 118617 146750 120805
rect 146710 118611 146762 118617
rect 146710 118553 146762 118559
rect 146708 118502 146764 118511
rect 146708 118437 146764 118446
rect 146722 118321 146750 118437
rect 146710 118315 146762 118321
rect 146710 118257 146762 118263
rect 146708 116726 146764 116735
rect 146708 116661 146764 116670
rect 146722 115287 146750 116661
rect 146710 115281 146762 115287
rect 146710 115223 146762 115229
rect 146708 114210 146764 114219
rect 146708 114145 146764 114154
rect 146722 112697 146750 114145
rect 146710 112691 146762 112697
rect 146710 112633 146762 112639
rect 146708 112434 146764 112443
rect 146708 112369 146710 112378
rect 146762 112369 146764 112378
rect 146710 112337 146762 112343
rect 146708 109770 146764 109779
rect 146708 109705 146764 109714
rect 146722 109515 146750 109705
rect 146710 109509 146762 109515
rect 146710 109451 146762 109457
rect 146708 107550 146764 107559
rect 146708 107485 146764 107494
rect 146722 106629 146750 107485
rect 146710 106623 146762 106629
rect 146710 106565 146762 106571
rect 146710 106475 146762 106481
rect 146710 106417 146762 106423
rect 146722 100783 146750 106417
rect 146710 100777 146762 100783
rect 146710 100719 146762 100725
rect 146708 85942 146764 85951
rect 146708 85877 146764 85886
rect 146722 85021 146750 85877
rect 146710 85015 146762 85021
rect 146710 84957 146762 84963
rect 146708 82390 146764 82399
rect 146708 82325 146764 82334
rect 146722 82135 146750 82325
rect 146710 82129 146762 82135
rect 146710 82071 146762 82077
rect 146708 79430 146764 79439
rect 146708 79365 146764 79374
rect 146722 77843 146750 79365
rect 146710 77837 146762 77843
rect 146710 77779 146762 77785
rect 146614 77763 146666 77769
rect 146614 77705 146666 77711
rect 146530 77612 146750 77640
rect 146614 77467 146666 77473
rect 146614 77409 146666 77415
rect 146516 75730 146572 75739
rect 146516 75665 146572 75674
rect 146530 75105 146558 75665
rect 146518 75099 146570 75105
rect 146518 75041 146570 75047
rect 146516 74990 146572 74999
rect 146516 74925 146572 74934
rect 146530 51943 146558 74925
rect 146518 51937 146570 51943
rect 146518 51879 146570 51885
rect 146422 50975 146474 50981
rect 146422 50917 146474 50923
rect 146626 50907 146654 77409
rect 146722 52165 146750 77612
rect 146818 66540 146846 132497
rect 146914 123797 146942 134296
rect 146902 123791 146954 123797
rect 146902 123733 146954 123739
rect 146900 121462 146956 121471
rect 146900 121397 146956 121406
rect 146914 121133 146942 121397
rect 146902 121127 146954 121133
rect 146902 121069 146954 121075
rect 146900 115986 146956 115995
rect 146900 115921 146956 115930
rect 146914 115583 146942 115921
rect 146902 115577 146954 115583
rect 146902 115519 146954 115525
rect 147010 115065 147038 134833
rect 147092 126938 147148 126947
rect 147092 126873 147094 126882
rect 147146 126873 147148 126882
rect 147094 126841 147146 126847
rect 146998 115059 147050 115065
rect 146998 115001 147050 115007
rect 148150 112469 148202 112475
rect 148150 112411 148202 112417
rect 148054 112395 148106 112401
rect 148054 112337 148106 112343
rect 147958 109583 148010 109589
rect 147958 109525 148010 109531
rect 147862 106697 147914 106703
rect 147862 106639 147914 106645
rect 146902 104847 146954 104853
rect 146902 104789 146954 104795
rect 146914 103669 146942 104789
rect 146902 103663 146954 103669
rect 146902 103605 146954 103611
rect 147766 100851 147818 100857
rect 147766 100793 147818 100799
rect 146818 66512 146942 66540
rect 146804 66406 146860 66415
rect 146804 66341 146860 66350
rect 146818 66299 146846 66341
rect 146806 66293 146858 66299
rect 146806 66235 146858 66241
rect 146914 66096 146942 66512
rect 146818 66068 146942 66096
rect 146818 65060 146846 66068
rect 146818 65032 146942 65060
rect 146914 64616 146942 65032
rect 146818 64588 146942 64616
rect 146710 52159 146762 52165
rect 146710 52101 146762 52107
rect 146614 50901 146666 50907
rect 146614 50843 146666 50849
rect 146818 50833 146846 64588
rect 146902 63407 146954 63413
rect 146902 63349 146954 63355
rect 146914 62419 146942 63349
rect 146900 62410 146956 62419
rect 146900 62345 146956 62354
rect 146900 60782 146956 60791
rect 146900 60717 146956 60726
rect 146914 60453 146942 60717
rect 146902 60447 146954 60453
rect 146902 60389 146954 60395
rect 146806 50827 146858 50833
rect 146806 50769 146858 50775
rect 146326 49939 146378 49945
rect 146326 49881 146378 49887
rect 147778 47725 147806 100793
rect 147766 47719 147818 47725
rect 147766 47661 147818 47667
rect 147874 47651 147902 106639
rect 147862 47645 147914 47651
rect 147862 47587 147914 47593
rect 147970 47577 147998 109525
rect 147958 47571 148010 47577
rect 147958 47513 148010 47519
rect 148066 47503 148094 112337
rect 148054 47497 148106 47503
rect 148054 47439 148106 47445
rect 148162 47429 148190 112411
rect 148150 47423 148202 47429
rect 148150 47365 148202 47371
rect 133618 46708 133646 46990
rect 133618 46680 133694 46708
rect 133666 42841 133694 46680
rect 148258 46245 148286 213125
rect 148354 74143 148382 237545
rect 149698 224511 149726 273065
rect 150274 272093 150302 277870
rect 150262 272087 150314 272093
rect 150262 272029 150314 272035
rect 151426 271427 151454 277870
rect 152674 273129 152702 277870
rect 153826 274609 153854 277870
rect 155088 277856 155486 277884
rect 153814 274603 153866 274609
rect 153814 274545 153866 274551
rect 152662 273123 152714 273129
rect 152662 273065 152714 273071
rect 155350 273123 155402 273129
rect 155350 273065 155402 273071
rect 151414 271421 151466 271427
rect 151414 271363 151466 271369
rect 152566 271421 152618 271427
rect 152566 271363 152618 271369
rect 151126 271125 151178 271131
rect 151126 271067 151178 271073
rect 151138 270835 151166 271067
rect 151126 270829 151178 270835
rect 151126 270771 151178 270777
rect 151126 230573 151178 230579
rect 151126 230515 151178 230521
rect 149686 224505 149738 224511
rect 149686 224447 149738 224453
rect 148438 204525 148490 204531
rect 148438 204467 148490 204473
rect 148342 74137 148394 74143
rect 148342 74079 148394 74085
rect 148342 60521 148394 60527
rect 148342 60463 148394 60469
rect 148354 54163 148382 60463
rect 148342 54157 148394 54163
rect 148342 54099 148394 54105
rect 148450 48613 148478 204467
rect 148534 184471 148586 184477
rect 148534 184413 148586 184419
rect 148438 48607 148490 48613
rect 148438 48549 148490 48555
rect 148546 46837 148574 184413
rect 148630 178699 148682 178705
rect 148630 178641 148682 178647
rect 148534 46831 148586 46837
rect 148534 46773 148586 46779
rect 148642 46541 148670 178641
rect 148726 161309 148778 161315
rect 148726 161251 148778 161257
rect 148738 46615 148766 161251
rect 148822 158497 148874 158503
rect 148822 158439 148874 158445
rect 148834 47133 148862 158439
rect 148918 155759 148970 155765
rect 148918 155701 148970 155707
rect 148822 47127 148874 47133
rect 148822 47069 148874 47075
rect 148930 46911 148958 155701
rect 149014 149913 149066 149919
rect 149014 149855 149066 149861
rect 148918 46905 148970 46911
rect 148918 46847 148970 46853
rect 149026 46689 149054 149855
rect 149108 149730 149164 149739
rect 149108 149665 149164 149674
rect 149122 48243 149150 149665
rect 149206 142587 149258 142593
rect 149206 142529 149258 142535
rect 149110 48237 149162 48243
rect 149110 48179 149162 48185
rect 149218 48169 149246 142529
rect 149302 136297 149354 136303
rect 149302 136239 149354 136245
rect 149206 48163 149258 48169
rect 149206 48105 149258 48111
rect 149314 48021 149342 136239
rect 149398 136001 149450 136007
rect 149398 135943 149450 135949
rect 149410 48095 149438 135943
rect 149494 126899 149546 126905
rect 149494 126841 149546 126847
rect 149398 48089 149450 48095
rect 149398 48031 149450 48037
rect 149302 48015 149354 48021
rect 149302 47957 149354 47963
rect 149506 47873 149534 126841
rect 149590 121127 149642 121133
rect 149590 121069 149642 121075
rect 149602 47947 149630 121069
rect 149686 115577 149738 115583
rect 149686 115519 149738 115525
rect 149590 47941 149642 47947
rect 149590 47883 149642 47889
rect 149494 47867 149546 47873
rect 149494 47809 149546 47815
rect 149698 47799 149726 115519
rect 151138 100561 151166 230515
rect 152578 224437 152606 271363
rect 155362 246975 155390 273065
rect 155348 246966 155404 246975
rect 155348 246901 155404 246910
rect 152566 224431 152618 224437
rect 152566 224373 152618 224379
rect 155458 221773 155486 277856
rect 156226 273129 156254 277870
rect 156884 273458 156940 273467
rect 156884 273393 156940 273402
rect 156214 273123 156266 273129
rect 156214 273065 156266 273071
rect 156898 272727 156926 273393
rect 157474 273351 157502 277870
rect 157462 273345 157514 273351
rect 156980 273310 157036 273319
rect 156980 273245 157036 273254
rect 157172 273310 157228 273319
rect 157462 273287 157514 273293
rect 157172 273245 157228 273254
rect 156692 272718 156748 272727
rect 156692 272653 156748 272662
rect 156884 272718 156940 272727
rect 156884 272653 156940 272662
rect 156706 271099 156734 272653
rect 156692 271090 156748 271099
rect 156692 271025 156748 271034
rect 156994 270951 157022 273245
rect 157186 271691 157214 273245
rect 158326 273123 158378 273129
rect 158326 273065 158378 273071
rect 157172 271682 157228 271691
rect 157172 271617 157228 271626
rect 156980 270942 157036 270951
rect 156980 270877 157036 270886
rect 156884 247706 156940 247715
rect 156884 247641 156940 247650
rect 156898 247271 156926 247641
rect 156884 247262 156940 247271
rect 156884 247197 156940 247206
rect 158338 245347 158366 273065
rect 158626 264545 158654 277870
rect 158806 273715 158858 273721
rect 158806 273657 158858 273663
rect 158818 272981 158846 273657
rect 158806 272975 158858 272981
rect 158806 272917 158858 272923
rect 159874 270021 159902 277870
rect 160726 273641 160778 273647
rect 160726 273583 160778 273589
rect 160738 272852 160766 273583
rect 161026 273425 161054 277870
rect 161206 274603 161258 274609
rect 161206 274545 161258 274551
rect 161014 273419 161066 273425
rect 161014 273361 161066 273367
rect 161218 273296 161246 274545
rect 161218 273268 161342 273296
rect 161314 273203 161342 273268
rect 161302 273197 161354 273203
rect 161302 273139 161354 273145
rect 162178 273129 162206 277870
rect 163440 277856 164030 277884
rect 162166 273123 162218 273129
rect 162166 273065 162218 273071
rect 161206 272901 161258 272907
rect 160738 272849 161206 272852
rect 160738 272843 161258 272849
rect 160738 272824 161246 272843
rect 160534 272753 160586 272759
rect 160534 272695 160586 272701
rect 161206 272753 161258 272759
rect 161206 272695 161258 272701
rect 160546 272556 160574 272695
rect 161218 272556 161246 272695
rect 160546 272528 161246 272556
rect 159862 270015 159914 270021
rect 159862 269957 159914 269963
rect 161110 270015 161162 270021
rect 161110 269957 161162 269963
rect 158614 264539 158666 264545
rect 158614 264481 158666 264487
rect 161122 247715 161150 269957
rect 161206 264539 161258 264545
rect 161206 264481 161258 264487
rect 161108 247706 161164 247715
rect 161108 247641 161164 247650
rect 158324 245338 158380 245347
rect 158324 245273 158380 245282
rect 161218 242387 161246 264481
rect 161302 246261 161354 246267
rect 161354 246209 161438 246212
rect 161302 246203 161438 246209
rect 161314 246193 161438 246203
rect 161314 246187 161450 246193
rect 161314 246184 161398 246187
rect 161398 246129 161450 246135
rect 164002 245939 164030 277856
rect 164278 273197 164330 273203
rect 164278 273139 164330 273145
rect 164086 273123 164138 273129
rect 164086 273065 164138 273071
rect 163988 245930 164044 245939
rect 163988 245865 164044 245874
rect 157940 242378 157996 242387
rect 157940 242313 157996 242322
rect 161204 242378 161260 242387
rect 161204 242313 161260 242322
rect 157954 242123 157982 242313
rect 161110 242265 161162 242271
rect 161110 242207 161162 242213
rect 157942 242117 157994 242123
rect 157942 242059 157994 242065
rect 161122 242049 161150 242207
rect 161204 242082 161260 242091
rect 161110 242043 161162 242049
rect 161204 242017 161260 242026
rect 161110 241985 161162 241991
rect 159766 228797 159818 228803
rect 159766 228739 159818 228745
rect 156886 226429 156938 226435
rect 156886 226371 156938 226377
rect 155446 221767 155498 221773
rect 155446 221709 155498 221715
rect 154006 213257 154058 213263
rect 154006 213199 154058 213205
rect 151222 190169 151274 190175
rect 151222 190111 151274 190117
rect 151126 100555 151178 100561
rect 151126 100497 151178 100503
rect 151234 94863 151262 190111
rect 151414 129711 151466 129717
rect 151414 129653 151466 129659
rect 151318 103811 151370 103817
rect 151318 103753 151370 103759
rect 151222 94857 151274 94863
rect 151222 94799 151274 94805
rect 151222 89455 151274 89461
rect 151222 89397 151274 89403
rect 151126 77911 151178 77917
rect 151126 77853 151178 77859
rect 149782 70289 149834 70295
rect 149782 70231 149834 70237
rect 149794 69037 149822 70231
rect 149782 69031 149834 69037
rect 149782 68973 149834 68979
rect 149782 62519 149834 62525
rect 149782 62461 149834 62467
rect 149794 60379 149822 62461
rect 149782 60373 149834 60379
rect 149782 60315 149834 60321
rect 151138 52461 151166 77853
rect 151234 71997 151262 89397
rect 151222 71991 151274 71997
rect 151222 71933 151274 71939
rect 151222 60595 151274 60601
rect 151222 60537 151274 60543
rect 151234 54681 151262 60537
rect 151222 54675 151274 54681
rect 151222 54617 151274 54623
rect 151330 52609 151358 103753
rect 151426 83541 151454 129653
rect 154018 97897 154046 213199
rect 154102 144363 154154 144369
rect 154102 144305 154154 144311
rect 154006 97891 154058 97897
rect 154006 97833 154058 97839
rect 154006 92267 154058 92273
rect 154006 92209 154058 92215
rect 151414 83535 151466 83541
rect 151414 83477 151466 83483
rect 154018 74883 154046 92209
rect 154114 86427 154142 144305
rect 156898 97823 156926 226371
rect 156982 167303 157034 167309
rect 156982 167245 157034 167251
rect 156886 97817 156938 97823
rect 156886 97759 156938 97765
rect 156994 89239 157022 167245
rect 157078 101591 157130 101597
rect 157078 101533 157130 101539
rect 156982 89233 157034 89239
rect 156982 89175 157034 89181
rect 154102 86421 154154 86427
rect 154102 86363 154154 86369
rect 157090 77769 157118 101533
rect 157078 77763 157130 77769
rect 157078 77705 157130 77711
rect 156982 75025 157034 75031
rect 156982 74967 157034 74973
rect 154006 74877 154058 74883
rect 154006 74819 154058 74825
rect 154678 72065 154730 72071
rect 154678 72007 154730 72013
rect 154690 68963 154718 72007
rect 154678 68957 154730 68963
rect 154678 68899 154730 68905
rect 156994 68889 157022 74967
rect 156982 68883 157034 68889
rect 156982 68825 157034 68831
rect 152662 67255 152714 67261
rect 152662 67197 152714 67203
rect 152674 66151 152702 67197
rect 158326 66441 158378 66447
rect 158326 66383 158378 66389
rect 152662 66145 152714 66151
rect 152662 66087 152714 66093
rect 158338 66077 158366 66383
rect 158326 66071 158378 66077
rect 158326 66013 158378 66019
rect 156310 60743 156362 60749
rect 156310 60685 156362 60691
rect 152662 60669 152714 60675
rect 152662 60611 152714 60617
rect 152674 56531 152702 60611
rect 156322 57123 156350 60685
rect 156310 57117 156362 57123
rect 156310 57059 156362 57065
rect 152662 56525 152714 56531
rect 152662 56467 152714 56473
rect 151318 52603 151370 52609
rect 151318 52545 151370 52551
rect 151126 52455 151178 52461
rect 151126 52397 151178 52403
rect 149686 47793 149738 47799
rect 149686 47735 149738 47741
rect 149014 46683 149066 46689
rect 149014 46625 149066 46631
rect 148726 46609 148778 46615
rect 148726 46551 148778 46557
rect 148630 46535 148682 46541
rect 148630 46477 148682 46483
rect 159778 46393 159806 228739
rect 161218 221699 161246 242017
rect 162742 240489 162794 240495
rect 162742 240431 162794 240437
rect 162754 237651 162782 240431
rect 162740 237642 162796 237651
rect 162740 237577 162796 237586
rect 162646 227687 162698 227693
rect 162646 227629 162698 227635
rect 161206 221693 161258 221699
rect 161206 221635 161258 221641
rect 159862 171299 159914 171305
rect 159862 171241 159914 171247
rect 159874 89165 159902 171241
rect 159958 104255 160010 104261
rect 159958 104197 160010 104203
rect 159862 89159 159914 89165
rect 159862 89101 159914 89107
rect 159970 77695 159998 104197
rect 159958 77689 160010 77695
rect 159958 77631 160010 77637
rect 160150 75099 160202 75105
rect 160150 75041 160202 75047
rect 160162 68815 160190 75041
rect 161494 74951 161546 74957
rect 161494 74893 161546 74899
rect 161506 71923 161534 74893
rect 161494 71917 161546 71923
rect 161494 71859 161546 71865
rect 160150 68809 160202 68815
rect 160150 68751 160202 68757
rect 160534 60817 160586 60823
rect 160534 60759 160586 60765
rect 160546 59639 160574 60759
rect 160534 59633 160586 59639
rect 160534 59575 160586 59581
rect 161300 52198 161356 52207
rect 161300 52133 161302 52142
rect 161354 52133 161356 52142
rect 161302 52101 161354 52107
rect 159766 46387 159818 46393
rect 159766 46329 159818 46335
rect 148246 46239 148298 46245
rect 148246 46181 148298 46187
rect 162658 46171 162686 227629
rect 164098 221625 164126 273065
rect 164290 272093 164318 273139
rect 164278 272087 164330 272093
rect 164278 272029 164330 272035
rect 164578 272019 164606 277870
rect 165826 272093 165854 277870
rect 165814 272087 165866 272093
rect 165814 272029 165866 272035
rect 164566 272013 164618 272019
rect 164566 271955 164618 271961
rect 166772 271682 166828 271691
rect 166772 271617 166828 271626
rect 166786 270803 166814 271617
rect 166772 270794 166828 270803
rect 166772 270729 166828 270738
rect 166882 246087 166910 277870
rect 166966 272087 167018 272093
rect 166966 272029 167018 272035
rect 166868 246078 166924 246087
rect 166868 246013 166924 246022
rect 165526 230499 165578 230505
rect 165526 230441 165578 230447
rect 164086 221619 164138 221625
rect 164086 221561 164138 221567
rect 162742 172853 162794 172859
rect 162742 172795 162794 172801
rect 162754 89091 162782 172795
rect 162838 106623 162890 106629
rect 162838 106565 162890 106571
rect 162742 89085 162794 89091
rect 162742 89027 162794 89033
rect 162850 77621 162878 106565
rect 162838 77615 162890 77621
rect 162838 77557 162890 77563
rect 165538 48211 165566 230441
rect 166978 221551 167006 272029
rect 168130 271353 168158 277870
rect 169296 277856 169886 277884
rect 168118 271347 168170 271353
rect 168118 271289 168170 271295
rect 168598 245373 168650 245379
rect 168596 245338 168598 245347
rect 168650 245338 168652 245347
rect 168596 245273 168652 245282
rect 168406 236271 168458 236277
rect 168406 236213 168458 236219
rect 166966 221545 167018 221551
rect 166966 221487 167018 221493
rect 165622 207485 165674 207491
rect 165622 207427 165674 207433
rect 165634 94789 165662 207427
rect 165718 132671 165770 132677
rect 165718 132613 165770 132619
rect 165622 94783 165674 94789
rect 165622 94725 165674 94731
rect 165622 89381 165674 89387
rect 165622 89323 165674 89329
rect 165634 71849 165662 89323
rect 165730 83467 165758 132613
rect 165718 83461 165770 83467
rect 165718 83403 165770 83409
rect 165622 71843 165674 71849
rect 165622 71785 165674 71791
rect 165524 48202 165580 48211
rect 165524 48137 165580 48146
rect 168418 47915 168446 236213
rect 169858 221477 169886 277856
rect 170530 272093 170558 277870
rect 170518 272087 170570 272093
rect 170518 272029 170570 272035
rect 171682 271723 171710 277870
rect 172726 272087 172778 272093
rect 172726 272029 172778 272035
rect 171670 271717 171722 271723
rect 171670 271659 171722 271665
rect 171668 247262 171724 247271
rect 171668 247197 171724 247206
rect 171682 245199 171710 247197
rect 171764 246226 171820 246235
rect 171764 246161 171820 246170
rect 171778 245347 171806 246161
rect 172738 245791 172766 272029
rect 172930 271945 172958 277870
rect 174082 272093 174110 277870
rect 174070 272087 174122 272093
rect 174070 272029 174122 272035
rect 172918 271939 172970 271945
rect 172918 271881 172970 271887
rect 175330 271649 175358 277870
rect 175510 272087 175562 272093
rect 175510 272029 175562 272035
rect 175318 271643 175370 271649
rect 175318 271585 175370 271591
rect 172724 245782 172780 245791
rect 172724 245717 172780 245726
rect 175522 245643 175550 272029
rect 176482 271945 176510 277870
rect 177044 273458 177100 273467
rect 177044 273393 177100 273402
rect 177058 272727 177086 273393
rect 177428 273310 177484 273319
rect 177428 273245 177484 273254
rect 177044 272718 177100 272727
rect 177044 272653 177100 272662
rect 177236 272718 177292 272727
rect 177236 272653 177292 272662
rect 175606 271939 175658 271945
rect 175606 271881 175658 271887
rect 176470 271939 176522 271945
rect 176470 271881 176522 271887
rect 175508 245634 175564 245643
rect 175508 245569 175564 245578
rect 171764 245338 171820 245347
rect 171764 245273 171820 245282
rect 171668 245190 171724 245199
rect 171668 245125 171724 245134
rect 174166 236197 174218 236203
rect 174166 236139 174218 236145
rect 171286 233311 171338 233317
rect 171286 233253 171338 233259
rect 169846 221471 169898 221477
rect 169846 221413 169898 221419
rect 168502 207411 168554 207417
rect 168502 207353 168554 207359
rect 168514 94715 168542 207353
rect 168598 138369 168650 138375
rect 168598 138311 168650 138317
rect 168502 94709 168554 94715
rect 168502 94651 168554 94657
rect 168502 89307 168554 89313
rect 168502 89249 168554 89255
rect 168514 71775 168542 89249
rect 168610 83393 168638 138311
rect 168598 83387 168650 83393
rect 168598 83329 168650 83335
rect 168502 71769 168554 71775
rect 168502 71711 168554 71717
rect 171298 48655 171326 233253
rect 171382 213331 171434 213337
rect 171382 213273 171434 213279
rect 171394 94641 171422 213273
rect 171478 141181 171530 141187
rect 171478 141123 171530 141129
rect 171382 94635 171434 94641
rect 171382 94577 171434 94583
rect 171490 83319 171518 141123
rect 171574 92193 171626 92199
rect 171574 92135 171626 92141
rect 171478 83313 171530 83319
rect 171478 83255 171530 83261
rect 171586 71701 171614 92135
rect 171574 71695 171626 71701
rect 171574 71637 171626 71643
rect 171284 48646 171340 48655
rect 171284 48581 171340 48590
rect 174178 48507 174206 236139
rect 175618 218887 175646 271881
rect 177046 271273 177098 271279
rect 177046 271215 177098 271221
rect 177058 270909 177086 271215
rect 177250 271099 177278 272653
rect 177442 271099 177470 273245
rect 177634 272093 177662 277870
rect 178294 273715 178346 273721
rect 178294 273657 178346 273663
rect 177716 273310 177772 273319
rect 177716 273245 177772 273254
rect 177622 272087 177674 272093
rect 177622 272029 177674 272035
rect 177236 271090 177292 271099
rect 177236 271025 177292 271034
rect 177428 271090 177484 271099
rect 177428 271025 177484 271034
rect 177730 270951 177758 273245
rect 178306 273000 178334 273657
rect 178486 273049 178538 273055
rect 178306 272997 178486 273000
rect 178306 272991 178538 272997
rect 178306 272972 178526 272991
rect 178390 272087 178442 272093
rect 178390 272029 178442 272035
rect 177716 270942 177772 270951
rect 177046 270903 177098 270909
rect 177716 270877 177772 270886
rect 177046 270845 177098 270851
rect 177044 246670 177100 246679
rect 177044 246605 177100 246614
rect 177058 245939 177086 246605
rect 177044 245930 177100 245939
rect 177044 245865 177100 245874
rect 178402 245791 178430 272029
rect 178486 271939 178538 271945
rect 178486 271881 178538 271887
rect 178388 245782 178444 245791
rect 178388 245717 178444 245726
rect 177046 242043 177098 242049
rect 177046 241985 177098 241991
rect 175606 218881 175658 218887
rect 175606 218823 175658 218829
rect 174262 216069 174314 216075
rect 174262 216011 174314 216017
rect 174274 97749 174302 216011
rect 174358 146953 174410 146959
rect 174358 146895 174410 146901
rect 174262 97743 174314 97749
rect 174262 97685 174314 97691
rect 174370 86353 174398 146895
rect 174454 95153 174506 95159
rect 174454 95095 174506 95101
rect 174358 86347 174410 86353
rect 174358 86289 174410 86295
rect 174466 74809 174494 95095
rect 174454 74803 174506 74809
rect 174454 74745 174506 74751
rect 174164 48498 174220 48507
rect 174164 48433 174220 48442
rect 177058 48359 177086 241985
rect 177142 218955 177194 218961
rect 177142 218897 177194 218903
rect 177154 97675 177182 218897
rect 178498 218813 178526 271881
rect 178882 271575 178910 277870
rect 180034 272093 180062 277870
rect 180022 272087 180074 272093
rect 180022 272029 180074 272035
rect 179446 271939 179498 271945
rect 179446 271881 179498 271887
rect 179458 271723 179486 271881
rect 179446 271717 179498 271723
rect 179446 271659 179498 271665
rect 178870 271569 178922 271575
rect 178870 271511 178922 271517
rect 178580 270202 178636 270211
rect 178580 270137 178636 270146
rect 178594 269767 178622 270137
rect 178580 269758 178636 269767
rect 178580 269693 178636 269702
rect 181282 245768 181310 277870
rect 181366 272087 181418 272093
rect 181366 272029 181418 272035
rect 181462 272087 181514 272093
rect 181462 272029 181514 272035
rect 181378 245897 181406 272029
rect 181474 271353 181502 272029
rect 182434 271575 182462 277870
rect 183600 277856 184286 277884
rect 287734 277933 287786 277939
rect 191446 277875 191498 277881
rect 182422 271569 182474 271575
rect 182422 271511 182474 271517
rect 181462 271347 181514 271353
rect 181462 271289 181514 271295
rect 181558 246261 181610 246267
rect 181474 246209 181558 246212
rect 181474 246203 181610 246209
rect 181474 246193 181598 246203
rect 181462 246187 181598 246193
rect 181514 246184 181598 246187
rect 181462 246129 181514 246135
rect 181366 245891 181418 245897
rect 181366 245833 181418 245839
rect 181282 245740 181406 245768
rect 181378 245643 181406 245740
rect 181364 245634 181420 245643
rect 181364 245569 181420 245578
rect 181366 245521 181418 245527
rect 181268 245486 181324 245495
rect 181366 245463 181418 245469
rect 181268 245421 181324 245430
rect 181282 245379 181310 245421
rect 181270 245373 181322 245379
rect 181270 245315 181322 245321
rect 179926 221915 179978 221921
rect 179926 221857 179978 221863
rect 178486 218807 178538 218813
rect 178486 218749 178538 218755
rect 177238 149839 177290 149845
rect 177238 149781 177290 149787
rect 177142 97669 177194 97675
rect 177142 97611 177194 97617
rect 177250 86279 177278 149781
rect 177334 95079 177386 95085
rect 177334 95021 177386 95027
rect 177238 86273 177290 86279
rect 177238 86215 177290 86221
rect 177346 74735 177374 95021
rect 177334 74729 177386 74735
rect 177334 74671 177386 74677
rect 177044 48350 177100 48359
rect 177044 48285 177100 48294
rect 168404 47906 168460 47915
rect 168404 47841 168460 47850
rect 179938 47355 179966 221857
rect 181378 218739 181406 245463
rect 182806 221841 182858 221847
rect 182806 221783 182858 221789
rect 181366 218733 181418 218739
rect 181366 218675 181418 218681
rect 180022 152799 180074 152805
rect 180022 152741 180074 152747
rect 180034 86205 180062 152741
rect 180118 98113 180170 98119
rect 180118 98055 180170 98061
rect 180022 86199 180074 86205
rect 180022 86141 180074 86147
rect 180130 74661 180158 98055
rect 182818 97601 182846 221783
rect 184258 218665 184286 277856
rect 184738 271279 184766 277870
rect 185986 271353 186014 277870
rect 185974 271347 186026 271353
rect 185974 271289 186026 271295
rect 184726 271273 184778 271279
rect 184726 271215 184778 271221
rect 187030 271273 187082 271279
rect 187030 271215 187082 271221
rect 187042 245495 187070 271215
rect 186836 245486 186892 245495
rect 186836 245421 186892 245430
rect 187028 245486 187084 245495
rect 187028 245421 187084 245430
rect 186850 245028 186878 245421
rect 187028 245042 187084 245051
rect 186850 245000 187028 245028
rect 187028 244977 187084 244986
rect 184246 218659 184298 218665
rect 184246 218601 184298 218607
rect 187138 216001 187166 277870
rect 187220 273606 187276 273615
rect 187220 273541 187276 273550
rect 187234 271691 187262 273541
rect 187220 271682 187276 271691
rect 187220 271617 187276 271626
rect 188386 267547 188414 277870
rect 189538 271057 189566 277870
rect 190786 271871 190814 277870
rect 190774 271865 190826 271871
rect 190774 271807 190826 271813
rect 190582 271791 190634 271797
rect 190582 271733 190634 271739
rect 190594 271427 190622 271733
rect 190582 271421 190634 271427
rect 190582 271363 190634 271369
rect 189622 271125 189674 271131
rect 189622 271067 189674 271073
rect 189526 271051 189578 271057
rect 189526 270993 189578 270999
rect 189634 270835 189662 271067
rect 189622 270829 189674 270835
rect 189622 270771 189674 270777
rect 188372 267538 188428 267547
rect 188372 267473 188428 267482
rect 191458 252483 191486 277875
rect 191938 270761 191966 277870
rect 193090 275127 193118 277870
rect 194338 276533 194366 277870
rect 194326 276527 194378 276533
rect 194326 276469 194378 276475
rect 193078 275121 193130 275127
rect 193078 275063 193130 275069
rect 194516 273458 194572 273467
rect 194516 273393 194572 273402
rect 192886 271865 192938 271871
rect 192886 271807 192938 271813
rect 191926 270755 191978 270761
rect 191926 270697 191978 270703
rect 191446 252477 191498 252483
rect 191446 252419 191498 252425
rect 188180 247262 188236 247271
rect 188098 247220 188180 247248
rect 187892 247114 187948 247123
rect 187892 247049 187948 247058
rect 187906 247007 187934 247049
rect 187894 247001 187946 247007
rect 187700 246966 187756 246975
rect 187894 246943 187946 246949
rect 187700 246901 187756 246910
rect 187604 246818 187660 246827
rect 187604 246753 187660 246762
rect 187618 245324 187646 246753
rect 187714 246656 187742 246901
rect 187988 246670 188044 246679
rect 187714 246628 187988 246656
rect 187988 246605 188044 246614
rect 187988 245338 188044 245347
rect 187618 245296 187988 245324
rect 187988 245273 188044 245282
rect 187700 245190 187756 245199
rect 188098 245176 188126 247220
rect 188180 247197 188236 247206
rect 187756 245148 188126 245176
rect 187700 245125 187756 245134
rect 187126 215995 187178 216001
rect 187126 215937 187178 215943
rect 192898 215927 192926 271807
rect 194530 270803 194558 273393
rect 195190 271273 195242 271279
rect 195190 271215 195242 271221
rect 195202 270909 195230 271215
rect 195490 270983 195518 277870
rect 196738 275275 196766 277870
rect 196726 275269 196778 275275
rect 196726 275211 196778 275217
rect 197588 273310 197644 273319
rect 197588 273245 197644 273254
rect 197204 272718 197260 272727
rect 197204 272653 197260 272662
rect 197218 271099 197246 272653
rect 197204 271090 197260 271099
rect 197204 271025 197260 271034
rect 195478 270977 195530 270983
rect 197602 270951 197630 273245
rect 195478 270919 195530 270925
rect 197588 270942 197644 270951
rect 195190 270903 195242 270909
rect 197588 270877 197644 270886
rect 195190 270845 195242 270851
rect 194516 270794 194572 270803
rect 194516 270729 194572 270738
rect 195874 270308 195998 270336
rect 195874 270211 195902 270308
rect 195860 270202 195916 270211
rect 195860 270137 195916 270146
rect 195970 270063 195998 270308
rect 195956 270054 196012 270063
rect 195956 269989 196012 269998
rect 197890 265063 197918 277870
rect 199138 270909 199166 277870
rect 200194 275423 200222 277870
rect 200182 275417 200234 275423
rect 200182 275359 200234 275365
rect 199126 270903 199178 270909
rect 199126 270845 199178 270851
rect 201442 266173 201470 277870
rect 202594 270835 202622 277870
rect 202582 270829 202634 270835
rect 202582 270771 202634 270777
rect 203842 269133 203870 277870
rect 204994 275867 205022 277870
rect 204982 275861 205034 275867
rect 204982 275803 205034 275809
rect 205846 271791 205898 271797
rect 205846 271733 205898 271739
rect 203830 269127 203882 269133
rect 203830 269069 203882 269075
rect 201430 266167 201482 266173
rect 201430 266109 201482 266115
rect 197878 265057 197930 265063
rect 197878 264999 197930 265005
rect 193270 252477 193322 252483
rect 193270 252419 193322 252425
rect 193282 244861 193310 252419
rect 205858 247451 205886 271733
rect 206242 270761 206270 277870
rect 207394 274165 207422 277870
rect 207382 274159 207434 274165
rect 207382 274101 207434 274107
rect 207284 273606 207340 273615
rect 207284 273541 207340 273550
rect 207298 271691 207326 273541
rect 207284 271682 207340 271691
rect 207284 271617 207340 271626
rect 206998 271421 207050 271427
rect 206998 271363 207050 271369
rect 207094 271421 207146 271427
rect 207094 271363 207146 271369
rect 206230 270755 206282 270761
rect 206230 270697 206282 270703
rect 205942 269275 205994 269281
rect 205942 269217 205994 269223
rect 205846 247445 205898 247451
rect 205846 247387 205898 247393
rect 201526 247001 201578 247007
rect 201524 246966 201526 246975
rect 201578 246966 201580 246975
rect 201524 246901 201580 246910
rect 204982 246927 205034 246933
rect 204982 246869 205034 246875
rect 204694 246853 204746 246859
rect 204694 246795 204746 246801
rect 202100 246522 202156 246531
rect 202100 246457 202156 246466
rect 193270 244855 193322 244861
rect 193270 244797 193322 244803
rect 198934 244781 198986 244787
rect 202114 244755 202142 246457
rect 202582 246261 202634 246267
rect 202582 246203 202634 246209
rect 202594 245749 202622 246203
rect 202582 245743 202634 245749
rect 202582 245685 202634 245691
rect 202198 245447 202250 245453
rect 202198 245389 202250 245395
rect 202210 245347 202238 245389
rect 202196 245338 202252 245347
rect 202196 245273 202252 245282
rect 198934 244723 198986 244729
rect 202100 244746 202156 244755
rect 198946 240019 198974 244723
rect 202100 244681 202156 244690
rect 204502 244189 204554 244195
rect 204502 244131 204554 244137
rect 198932 240010 198988 240019
rect 198932 239945 198988 239954
rect 204514 227735 204542 244131
rect 204598 243967 204650 243973
rect 204598 243909 204650 243915
rect 204500 227726 204556 227735
rect 204500 227661 204556 227670
rect 202966 227613 203018 227619
rect 202966 227555 203018 227561
rect 200086 224727 200138 224733
rect 200086 224669 200138 224675
rect 192886 215921 192938 215927
rect 192886 215863 192938 215869
rect 197206 201639 197258 201645
rect 197206 201581 197258 201587
rect 188566 198901 188618 198907
rect 188566 198843 188618 198849
rect 185686 195867 185738 195873
rect 185686 195809 185738 195815
rect 182902 152725 182954 152731
rect 182902 152667 182954 152673
rect 182806 97595 182858 97601
rect 182806 97537 182858 97543
rect 182914 86131 182942 152667
rect 182998 98039 183050 98045
rect 182998 97981 183050 97987
rect 182902 86125 182954 86131
rect 182902 86067 182954 86073
rect 180118 74655 180170 74661
rect 180118 74597 180170 74603
rect 183010 74587 183038 97981
rect 182998 74581 183050 74587
rect 182998 74523 183050 74529
rect 181364 52198 181420 52207
rect 181364 52133 181366 52142
rect 181418 52133 181420 52142
rect 181366 52101 181418 52107
rect 179926 47349 179978 47355
rect 179926 47291 179978 47297
rect 185698 47281 185726 195809
rect 185782 175739 185834 175745
rect 185782 175681 185834 175687
rect 185794 89017 185822 175681
rect 185878 109509 185930 109515
rect 185878 109451 185930 109457
rect 185782 89011 185834 89017
rect 185782 88953 185834 88959
rect 185890 77547 185918 109451
rect 185878 77541 185930 77547
rect 185878 77483 185930 77489
rect 188578 48465 188606 198843
rect 191446 198827 191498 198833
rect 191446 198769 191498 198775
rect 188662 181511 188714 181517
rect 188662 181453 188714 181459
rect 188674 91829 188702 181453
rect 188758 118315 188810 118321
rect 188758 118257 188810 118263
rect 188662 91823 188714 91829
rect 188662 91765 188714 91771
rect 188770 80359 188798 118257
rect 191458 100487 191486 198769
rect 194326 198753 194378 198759
rect 194326 198695 194378 198701
rect 191542 178625 191594 178631
rect 191542 178567 191594 178573
rect 191446 100481 191498 100487
rect 191446 100423 191498 100429
rect 191554 88943 191582 178567
rect 191638 112691 191690 112697
rect 191638 112633 191690 112639
rect 191542 88937 191594 88943
rect 191542 88879 191594 88885
rect 188758 80353 188810 80359
rect 188758 80295 188810 80301
rect 189910 77763 189962 77769
rect 189910 77705 189962 77711
rect 189922 77473 189950 77705
rect 189910 77467 189962 77473
rect 189910 77409 189962 77415
rect 191650 77399 191678 112633
rect 191638 77393 191690 77399
rect 191638 77335 191690 77341
rect 188566 48459 188618 48465
rect 188566 48401 188618 48407
rect 185686 47275 185738 47281
rect 185686 47217 185738 47223
rect 194338 46985 194366 198695
rect 194422 184397 194474 184403
rect 194422 184339 194474 184345
rect 194434 91903 194462 184339
rect 194518 118611 194570 118617
rect 194518 118553 194570 118559
rect 194422 91897 194474 91903
rect 194422 91839 194474 91845
rect 194530 80433 194558 118553
rect 194518 80427 194570 80433
rect 194518 80369 194570 80375
rect 197218 48317 197246 201581
rect 197302 187283 197354 187289
rect 197302 187225 197354 187231
rect 197314 91977 197342 187225
rect 197398 124087 197450 124093
rect 197398 124029 197450 124035
rect 197302 91971 197354 91977
rect 197302 91913 197354 91919
rect 197410 80507 197438 124029
rect 197398 80501 197450 80507
rect 197398 80443 197450 80449
rect 197206 48311 197258 48317
rect 197206 48253 197258 48259
rect 200098 47059 200126 224669
rect 200182 155685 200234 155691
rect 200182 155627 200234 155633
rect 200194 92051 200222 155627
rect 200278 123939 200330 123945
rect 200278 123881 200330 123887
rect 200182 92045 200234 92051
rect 200182 91987 200234 91993
rect 200290 80581 200318 123881
rect 200278 80575 200330 80581
rect 200278 80517 200330 80523
rect 202978 47207 203006 227555
rect 204610 225492 204638 243909
rect 204706 230991 204734 246795
rect 204790 246779 204842 246785
rect 204790 246721 204842 246727
rect 204802 231583 204830 246721
rect 204886 246409 204938 246415
rect 204886 246351 204938 246357
rect 204898 232175 204926 246351
rect 204884 232166 204940 232175
rect 204994 232133 205022 246869
rect 205750 244633 205802 244639
rect 205750 244575 205802 244581
rect 205462 244485 205514 244491
rect 205462 244427 205514 244433
rect 205270 244411 205322 244417
rect 205270 244353 205322 244359
rect 205078 244337 205130 244343
rect 205078 244279 205130 244285
rect 204884 232101 204940 232110
rect 204982 232127 205034 232133
rect 204982 232069 205034 232075
rect 205090 232004 205118 244279
rect 205174 243449 205226 243455
rect 205174 243391 205226 243397
rect 204898 231976 205118 232004
rect 204788 231574 204844 231583
rect 204788 231509 204844 231518
rect 204692 230982 204748 230991
rect 204692 230917 204748 230926
rect 204898 226699 204926 231976
rect 205186 228327 205214 243391
rect 205172 228318 205228 228327
rect 205172 228253 205228 228262
rect 205078 227465 205130 227471
rect 205078 227407 205130 227413
rect 204884 226690 204940 226699
rect 204884 226625 204940 226634
rect 204610 225464 204926 225492
rect 204502 224653 204554 224659
rect 204502 224595 204554 224601
rect 204514 224035 204542 224595
rect 204598 224505 204650 224511
rect 204598 224447 204650 224453
rect 204500 224026 204556 224035
rect 204500 223961 204556 223970
rect 204610 222851 204638 224447
rect 204596 222842 204652 222851
rect 204596 222777 204652 222786
rect 204502 221767 204554 221773
rect 204502 221709 204554 221715
rect 204514 221223 204542 221709
rect 204598 221471 204650 221477
rect 204598 221413 204650 221419
rect 204500 221214 204556 221223
rect 204500 221149 204556 221158
rect 204610 219447 204638 221413
rect 204596 219438 204652 219447
rect 204596 219373 204652 219382
rect 204502 218881 204554 218887
rect 204502 218823 204554 218829
rect 204514 218559 204542 218823
rect 204598 218807 204650 218813
rect 204598 218749 204650 218755
rect 204500 218550 204556 218559
rect 204500 218485 204556 218494
rect 204610 217967 204638 218749
rect 204694 218733 204746 218739
rect 204694 218675 204746 218681
rect 204596 217958 204652 217967
rect 204596 217893 204652 217902
rect 204706 217819 204734 218675
rect 204692 217810 204748 217819
rect 204692 217745 204748 217754
rect 204790 215995 204842 216001
rect 204790 215937 204842 215943
rect 204502 215921 204554 215927
rect 204802 215895 204830 215937
rect 204502 215863 204554 215869
rect 204788 215886 204844 215895
rect 204514 215303 204542 215863
rect 204788 215821 204844 215830
rect 204500 215294 204556 215303
rect 204500 215229 204556 215238
rect 204898 212935 204926 225464
rect 204982 221693 205034 221699
rect 204982 221635 205034 221641
rect 204994 221075 205022 221635
rect 204980 221066 205036 221075
rect 204980 221001 205036 221010
rect 204884 212926 204940 212935
rect 204884 212861 204940 212870
rect 205090 212764 205118 227407
rect 205282 226107 205310 244353
rect 205268 226098 205324 226107
rect 205268 226033 205324 226042
rect 205474 225663 205502 244427
rect 205654 244263 205706 244269
rect 205654 244205 205706 244211
rect 205556 232314 205612 232323
rect 205556 232249 205612 232258
rect 205570 232133 205598 232249
rect 205558 232127 205610 232133
rect 205558 232069 205610 232075
rect 205460 225654 205516 225663
rect 205460 225589 205516 225598
rect 205462 224579 205514 224585
rect 205462 224521 205514 224527
rect 205474 223443 205502 224521
rect 205460 223434 205516 223443
rect 205460 223369 205516 223378
rect 205366 221619 205418 221625
rect 205366 221561 205418 221567
rect 205378 220187 205406 221561
rect 205364 220178 205420 220187
rect 205364 220113 205420 220122
rect 205366 218659 205418 218665
rect 205366 218601 205418 218607
rect 205378 216931 205406 218601
rect 205364 216922 205420 216931
rect 205364 216857 205420 216866
rect 205570 213189 205598 232069
rect 205666 227291 205694 244205
rect 205652 227282 205708 227291
rect 205652 227217 205708 227226
rect 205762 224479 205790 244575
rect 205846 242043 205898 242049
rect 205846 241985 205898 241991
rect 205748 224470 205804 224479
rect 205748 224405 205804 224414
rect 205858 224308 205886 241985
rect 205954 236425 205982 269217
rect 207010 266659 207038 271363
rect 207106 271057 207134 271363
rect 207094 271051 207146 271057
rect 207094 270993 207146 270999
rect 207190 271051 207242 271057
rect 207190 270993 207242 270999
rect 207202 270687 207230 270993
rect 207190 270681 207242 270687
rect 207190 270623 207242 270629
rect 206996 266650 207052 266659
rect 206996 266585 207052 266594
rect 208546 266321 208574 277870
rect 209794 273499 209822 277870
rect 209686 273493 209738 273499
rect 209686 273435 209738 273441
rect 209782 273493 209834 273499
rect 209782 273435 209834 273441
rect 209698 271871 209726 273435
rect 209686 271865 209738 271871
rect 209686 271807 209738 271813
rect 210946 268393 210974 277870
rect 212194 276607 212222 277870
rect 212182 276601 212234 276607
rect 212182 276543 212234 276549
rect 211606 273567 211658 273573
rect 211606 273509 211658 273515
rect 210934 268387 210986 268393
rect 210934 268329 210986 268335
rect 208534 266315 208586 266321
rect 208534 266257 208586 266263
rect 211508 261904 211564 261913
rect 211508 261839 211564 261848
rect 207284 255402 207340 255411
rect 207284 255337 207340 255346
rect 206806 252033 206858 252039
rect 206806 251975 206858 251981
rect 206422 244115 206474 244121
rect 206422 244057 206474 244063
rect 206230 244041 206282 244047
rect 206230 243983 206282 243989
rect 206038 243671 206090 243677
rect 206038 243613 206090 243619
rect 205942 236419 205994 236425
rect 205942 236361 205994 236367
rect 205942 236197 205994 236203
rect 205942 236139 205994 236145
rect 205954 230547 205982 236139
rect 205940 230538 205996 230547
rect 205940 230473 205996 230482
rect 206050 229192 206078 243613
rect 206134 243375 206186 243381
rect 206134 243317 206186 243323
rect 206146 229363 206174 243317
rect 206132 229354 206188 229363
rect 206132 229289 206188 229298
rect 206050 229164 206174 229192
rect 206146 224881 206174 229164
rect 206134 224875 206186 224881
rect 206134 224817 206186 224823
rect 206134 224653 206186 224659
rect 206134 224595 206186 224601
rect 205666 224280 205886 224308
rect 205558 213183 205610 213189
rect 205558 213125 205610 213131
rect 204898 212736 205118 212764
rect 204898 210271 204926 212736
rect 204884 210262 204940 210271
rect 204884 210197 204940 210206
rect 205076 210262 205132 210271
rect 205076 210197 205132 210206
rect 205090 190175 205118 210197
rect 205666 202723 205694 224280
rect 206146 214711 206174 224595
rect 206132 214702 206188 214711
rect 206132 214637 206188 214646
rect 206242 212047 206270 243983
rect 206326 243745 206378 243751
rect 206326 243687 206378 243693
rect 206338 214563 206366 243687
rect 206434 224585 206462 244057
rect 206614 243893 206666 243899
rect 206614 243835 206666 243841
rect 206518 243819 206570 243825
rect 206518 243761 206570 243767
rect 206422 224579 206474 224585
rect 206422 224521 206474 224527
rect 206422 224431 206474 224437
rect 206422 224373 206474 224379
rect 206434 221815 206462 224373
rect 206420 221806 206476 221815
rect 206420 221741 206476 221750
rect 206324 214554 206380 214563
rect 206324 214489 206380 214498
rect 206530 213675 206558 243761
rect 206516 213666 206572 213675
rect 206516 213601 206572 213610
rect 206626 213083 206654 243835
rect 206710 243597 206762 243603
rect 206710 243539 206762 243545
rect 206722 216339 206750 243539
rect 206818 229955 206846 251975
rect 206900 249926 206956 249935
rect 206900 249861 206956 249870
rect 206914 244732 206942 249861
rect 206914 244704 207134 244732
rect 206998 244559 207050 244565
rect 206998 244501 207050 244507
rect 206902 243523 206954 243529
rect 206902 243465 206954 243471
rect 206804 229946 206860 229955
rect 206804 229881 206860 229890
rect 206806 224579 206858 224585
rect 206806 224521 206858 224527
rect 206708 216330 206764 216339
rect 206708 216265 206764 216274
rect 206612 213074 206668 213083
rect 206612 213009 206668 213018
rect 206228 212038 206284 212047
rect 206228 211973 206284 211982
rect 206818 211455 206846 224521
rect 206914 222407 206942 243465
rect 207010 225071 207038 244501
rect 207106 237609 207134 244704
rect 207298 243423 207326 255337
rect 210646 252107 210698 252113
rect 210646 252049 210698 252055
rect 210166 246705 210218 246711
rect 210166 246647 210218 246653
rect 209686 246335 209738 246341
rect 209686 246277 209738 246283
rect 209698 244861 209726 246277
rect 210178 244935 210206 246647
rect 210550 246483 210602 246489
rect 210550 246425 210602 246431
rect 210562 245495 210590 246425
rect 210548 245486 210604 245495
rect 210548 245421 210604 245430
rect 210166 244929 210218 244935
rect 210166 244871 210218 244877
rect 209686 244855 209738 244861
rect 209686 244797 209738 244803
rect 207284 243414 207340 243423
rect 207284 243349 207340 243358
rect 208724 240010 208780 240019
rect 208724 239945 208780 239954
rect 208738 239131 208766 239945
rect 208724 239122 208780 239131
rect 208724 239057 208780 239066
rect 209876 239122 209932 239131
rect 209876 239057 209932 239066
rect 207094 237603 207146 237609
rect 207094 237545 207146 237551
rect 209780 236754 209836 236763
rect 209780 236689 209836 236698
rect 209684 236606 209740 236615
rect 209684 236541 209740 236550
rect 208054 233607 208106 233613
rect 208054 233549 208106 233555
rect 207380 232166 207436 232175
rect 207380 232101 207436 232110
rect 207092 229946 207148 229955
rect 207092 229881 207148 229890
rect 206996 225062 207052 225071
rect 206996 224997 207052 225006
rect 206900 222398 206956 222407
rect 206900 222333 206956 222342
rect 206902 221545 206954 221551
rect 206902 221487 206954 221493
rect 206914 219595 206942 221487
rect 206900 219586 206956 219595
rect 206900 219521 206956 219530
rect 206804 211446 206860 211455
rect 206804 211381 206860 211390
rect 205652 202714 205708 202723
rect 205652 202649 205708 202658
rect 204886 190169 204938 190175
rect 204886 190111 204938 190117
rect 205078 190169 205130 190175
rect 205078 190111 205130 190117
rect 204898 187215 204926 190111
rect 204886 187209 204938 187215
rect 204886 187151 204938 187157
rect 205078 187209 205130 187215
rect 205078 187151 205130 187157
rect 206998 187209 207050 187215
rect 206998 187151 207050 187157
rect 203062 155611 203114 155617
rect 203062 155553 203114 155559
rect 203074 92125 203102 155553
rect 205090 152676 205118 187151
rect 207010 162943 207038 187151
rect 206998 162937 207050 162943
rect 206998 162879 207050 162885
rect 204994 152648 205118 152676
rect 204994 145424 205022 152648
rect 204898 145396 205022 145424
rect 203158 126825 203210 126831
rect 203158 126767 203210 126773
rect 203062 92119 203114 92125
rect 203062 92061 203114 92067
rect 203170 80655 203198 126767
rect 204898 126683 204926 145396
rect 204790 126677 204842 126683
rect 204790 126619 204842 126625
rect 204886 126677 204938 126683
rect 204886 126619 204938 126625
rect 204802 106629 204830 126619
rect 204790 106623 204842 106629
rect 204790 106565 204842 106571
rect 204982 106623 205034 106629
rect 204982 106565 205034 106571
rect 204502 103589 204554 103595
rect 204502 103531 204554 103537
rect 204514 102083 204542 103531
rect 204500 102074 204556 102083
rect 204500 102009 204556 102018
rect 204694 100777 204746 100783
rect 204694 100719 204746 100725
rect 204598 100629 204650 100635
rect 204598 100571 204650 100577
rect 204502 100555 204554 100561
rect 204502 100497 204554 100503
rect 204514 100455 204542 100497
rect 204500 100446 204556 100455
rect 204500 100381 204556 100390
rect 204610 100307 204638 100571
rect 204596 100298 204652 100307
rect 204596 100233 204652 100242
rect 204706 98679 204734 100719
rect 204790 100481 204842 100487
rect 204790 100423 204842 100429
rect 204802 99419 204830 100423
rect 204788 99410 204844 99419
rect 204788 99345 204844 99354
rect 204692 98670 204748 98679
rect 204692 98605 204748 98614
rect 204502 97817 204554 97823
rect 204500 97782 204502 97791
rect 204554 97782 204556 97791
rect 204500 97717 204556 97726
rect 204502 97595 204554 97601
rect 204502 97537 204554 97543
rect 204514 97199 204542 97537
rect 204500 97190 204556 97199
rect 204500 97125 204556 97134
rect 204598 94857 204650 94863
rect 204598 94799 204650 94805
rect 204500 94674 204556 94683
rect 204500 94609 204502 94618
rect 204554 94609 204556 94618
rect 204502 94577 204554 94583
rect 204610 93795 204638 94799
rect 204596 93786 204652 93795
rect 204596 93721 204652 93730
rect 204598 92119 204650 92125
rect 204598 92061 204650 92067
rect 204502 92045 204554 92051
rect 204610 92019 204638 92061
rect 204502 91987 204554 91993
rect 204596 92010 204652 92019
rect 204514 91279 204542 91987
rect 204596 91945 204652 91954
rect 204694 91971 204746 91977
rect 204694 91913 204746 91919
rect 204598 91897 204650 91903
rect 204598 91839 204650 91845
rect 204500 91270 204556 91279
rect 204500 91205 204556 91214
rect 204610 90095 204638 91839
rect 204706 90687 204734 91913
rect 204790 91823 204842 91829
rect 204790 91765 204842 91771
rect 204692 90678 204748 90687
rect 204692 90613 204748 90622
rect 204596 90086 204652 90095
rect 204596 90021 204652 90030
rect 204802 89651 204830 91765
rect 204788 89642 204844 89651
rect 204788 89577 204844 89586
rect 204994 89387 205022 106565
rect 206710 103663 206762 103669
rect 206710 103605 206762 103611
rect 206230 103515 206282 103521
rect 206230 103457 206282 103463
rect 206242 101047 206270 103457
rect 206722 101639 206750 103605
rect 206708 101630 206764 101639
rect 206708 101565 206764 101574
rect 206228 101038 206284 101047
rect 206228 100973 206284 100982
rect 206902 100703 206954 100709
rect 206902 100645 206954 100651
rect 206914 98827 206942 100645
rect 206900 98818 206956 98827
rect 206900 98753 206956 98762
rect 206518 97891 206570 97897
rect 206518 97833 206570 97839
rect 205270 97743 205322 97749
rect 205270 97685 205322 97691
rect 205282 96163 205310 97685
rect 206134 97669 206186 97675
rect 206134 97611 206186 97617
rect 206146 97051 206174 97611
rect 206132 97042 206188 97051
rect 206132 96977 206188 96986
rect 205268 96154 205324 96163
rect 205268 96089 205324 96098
rect 206530 95571 206558 97833
rect 206516 95562 206572 95571
rect 206516 95497 206572 95506
rect 206326 95005 206378 95011
rect 206326 94947 206378 94953
rect 205846 94783 205898 94789
rect 205846 94725 205898 94731
rect 205750 94709 205802 94715
rect 205750 94651 205802 94657
rect 205762 94535 205790 94651
rect 205748 94526 205804 94535
rect 205748 94461 205804 94470
rect 205858 93943 205886 94725
rect 205844 93934 205900 93943
rect 205844 93869 205900 93878
rect 206338 92315 206366 94947
rect 206902 94931 206954 94937
rect 206902 94873 206954 94879
rect 206914 92907 206942 94873
rect 206900 92898 206956 92907
rect 206900 92833 206956 92842
rect 206324 92306 206380 92315
rect 206324 92241 206380 92250
rect 204982 89381 205034 89387
rect 204982 89323 205034 89329
rect 205078 89307 205130 89313
rect 205078 89249 205130 89255
rect 204694 89233 204746 89239
rect 204694 89175 204746 89181
rect 204598 89085 204650 89091
rect 204598 89027 204650 89033
rect 204502 89011 204554 89017
rect 204502 88953 204554 88959
rect 204514 88467 204542 88953
rect 204500 88458 204556 88467
rect 204500 88393 204556 88402
rect 204610 88023 204638 89027
rect 204596 88014 204652 88023
rect 204596 87949 204652 87958
rect 204706 86839 204734 89175
rect 204788 89050 204844 89059
rect 204788 88985 204844 88994
rect 204802 88943 204830 88985
rect 204790 88937 204842 88943
rect 204790 88879 204842 88885
rect 204692 86830 204748 86839
rect 204692 86765 204748 86774
rect 204694 86421 204746 86427
rect 204500 86386 204556 86395
rect 204694 86363 204746 86369
rect 204500 86321 204556 86330
rect 204514 86131 204542 86321
rect 204598 86273 204650 86279
rect 204598 86215 204650 86221
rect 204502 86125 204554 86131
rect 204502 86067 204554 86073
rect 204500 85794 204556 85803
rect 204500 85729 204556 85738
rect 204514 85021 204542 85729
rect 204502 85015 204554 85021
rect 204502 84957 204554 84963
rect 204610 84767 204638 86215
rect 204596 84758 204652 84767
rect 204596 84693 204652 84702
rect 204706 83583 204734 86363
rect 204692 83574 204748 83583
rect 204692 83509 204748 83518
rect 204502 83313 204554 83319
rect 204502 83255 204554 83261
rect 204514 83139 204542 83255
rect 204500 83130 204556 83139
rect 204500 83065 204556 83074
rect 204502 82129 204554 82135
rect 204502 82071 204554 82077
rect 204514 81955 204542 82071
rect 204500 81946 204556 81955
rect 204500 81881 204556 81890
rect 203158 80649 203210 80655
rect 203158 80591 203210 80597
rect 204502 80575 204554 80581
rect 204502 80517 204554 80523
rect 204514 80179 204542 80517
rect 204598 80501 204650 80507
rect 204598 80443 204650 80449
rect 204500 80170 204556 80179
rect 204500 80105 204556 80114
rect 204610 79291 204638 80443
rect 204694 80427 204746 80433
rect 204694 80369 204746 80375
rect 204596 79282 204652 79291
rect 204596 79217 204652 79226
rect 204706 78699 204734 80369
rect 205090 80008 205118 89249
rect 206998 89233 207050 89239
rect 206998 89175 207050 89181
rect 205270 89159 205322 89165
rect 205270 89101 205322 89107
rect 205282 87431 205310 89101
rect 205268 87422 205324 87431
rect 205268 87357 205324 87366
rect 206614 86347 206666 86353
rect 206614 86289 206666 86295
rect 205558 86199 205610 86205
rect 205558 86141 205610 86147
rect 205570 85211 205598 86141
rect 205556 85202 205612 85211
rect 205556 85137 205612 85146
rect 206626 84175 206654 86289
rect 206612 84166 206668 84175
rect 206612 84101 206668 84110
rect 206230 83535 206282 83541
rect 206230 83477 206282 83483
rect 205750 83387 205802 83393
rect 205750 83329 205802 83335
rect 205762 82547 205790 83329
rect 205748 82538 205804 82547
rect 205748 82473 205804 82482
rect 206242 80919 206270 83477
rect 206710 83461 206762 83467
rect 206710 83403 206762 83409
rect 206722 81511 206750 83403
rect 206708 81502 206764 81511
rect 206708 81437 206764 81446
rect 206228 80910 206284 80919
rect 206228 80845 206284 80854
rect 205270 80649 205322 80655
rect 205270 80591 205322 80597
rect 205282 80327 205310 80591
rect 205268 80318 205324 80327
rect 205268 80253 205324 80262
rect 205090 79980 205310 80008
rect 204692 78690 204748 78699
rect 204692 78625 204748 78634
rect 204598 77763 204650 77769
rect 204598 77705 204650 77711
rect 204502 77615 204554 77621
rect 204502 77557 204554 77563
rect 204514 76035 204542 77557
rect 204610 77071 204638 77705
rect 204788 77654 204844 77663
rect 204788 77589 204844 77598
rect 204694 77467 204746 77473
rect 204694 77409 204746 77415
rect 204596 77062 204652 77071
rect 204596 76997 204652 77006
rect 204500 76026 204556 76035
rect 204500 75961 204556 75970
rect 204706 75295 204734 77409
rect 204802 77399 204830 77589
rect 204790 77393 204842 77399
rect 204790 77335 204842 77341
rect 204692 75286 204748 75295
rect 204692 75221 204748 75230
rect 204694 74877 204746 74883
rect 204694 74819 204746 74825
rect 204598 74729 204650 74735
rect 204598 74671 204650 74677
rect 204502 74581 204554 74587
rect 204502 74523 204554 74529
rect 204514 74407 204542 74523
rect 204500 74398 204556 74407
rect 204500 74333 204556 74342
rect 204610 73667 204638 74671
rect 204596 73658 204652 73667
rect 204596 73593 204652 73602
rect 204706 72187 204734 74819
rect 204692 72178 204748 72187
rect 204692 72113 204748 72122
rect 204982 71917 205034 71923
rect 204982 71859 205034 71865
rect 204598 71769 204650 71775
rect 204500 71734 204556 71743
rect 204598 71711 204650 71717
rect 204500 71669 204502 71678
rect 204554 71669 204556 71678
rect 204502 71637 204554 71643
rect 204610 71151 204638 71711
rect 204596 71142 204652 71151
rect 204596 71077 204652 71086
rect 204994 69523 205022 71859
rect 204980 69514 205036 69523
rect 204980 69449 205036 69458
rect 205282 69204 205310 79980
rect 206518 77689 206570 77695
rect 206518 77631 206570 77637
rect 205942 77541 205994 77547
rect 205942 77483 205994 77489
rect 205954 76923 205982 77483
rect 205940 76914 205996 76923
rect 205940 76849 205996 76858
rect 206530 75443 206558 77631
rect 206516 75434 206572 75443
rect 206516 75369 206572 75378
rect 206806 74803 206858 74809
rect 206806 74745 206858 74751
rect 205750 74655 205802 74661
rect 205750 74597 205802 74603
rect 205762 73815 205790 74597
rect 205748 73806 205804 73815
rect 205748 73741 205804 73750
rect 206818 72779 206846 74745
rect 206804 72770 206860 72779
rect 206804 72705 206860 72714
rect 206806 71991 206858 71997
rect 206806 71933 206858 71939
rect 205462 71843 205514 71849
rect 205462 71785 205514 71791
rect 205474 70559 205502 71785
rect 205460 70550 205516 70559
rect 205460 70485 205516 70494
rect 206818 69967 206846 71933
rect 206804 69958 206860 69967
rect 206804 69893 206860 69902
rect 205186 69176 205310 69204
rect 207010 69185 207038 89175
rect 206998 69179 207050 69185
rect 205186 69037 205214 69176
rect 206998 69121 207050 69127
rect 206518 69105 206570 69111
rect 206518 69047 206570 69053
rect 204118 69031 204170 69037
rect 204118 68973 204170 68979
rect 205174 69031 205226 69037
rect 205174 68973 205226 68979
rect 204130 67303 204158 68973
rect 204598 68957 204650 68963
rect 204500 68922 204556 68931
rect 204598 68899 204650 68905
rect 204500 68857 204556 68866
rect 204514 68815 204542 68857
rect 204502 68809 204554 68815
rect 204502 68751 204554 68757
rect 204610 67895 204638 68899
rect 206422 68883 206474 68889
rect 206422 68825 206474 68831
rect 206434 68339 206462 68825
rect 206420 68330 206476 68339
rect 206420 68265 206476 68274
rect 204596 67886 204652 67895
rect 204596 67821 204652 67830
rect 204116 67294 204172 67303
rect 204116 67229 204172 67238
rect 206530 66711 206558 69047
rect 206516 66702 206572 66711
rect 206516 66637 206572 66646
rect 204500 66258 204556 66267
rect 204500 66193 204556 66202
rect 205462 66219 205514 66225
rect 204514 66077 204542 66193
rect 205462 66161 205514 66167
rect 204502 66071 204554 66077
rect 204502 66013 204554 66019
rect 205474 65083 205502 66161
rect 206326 66145 206378 66151
rect 206326 66087 206378 66093
rect 206338 65675 206366 66087
rect 206324 65666 206380 65675
rect 206324 65601 206380 65610
rect 205460 65074 205516 65083
rect 205460 65009 205516 65018
rect 204598 64887 204650 64893
rect 204598 64829 204650 64835
rect 204502 64813 204554 64819
rect 204502 64755 204554 64761
rect 204514 64639 204542 64755
rect 204500 64630 204556 64639
rect 204500 64565 204556 64574
rect 204610 64047 204638 64829
rect 204596 64038 204652 64047
rect 204596 63973 204652 63982
rect 204500 63446 204556 63455
rect 204500 63381 204502 63390
rect 204554 63381 204556 63390
rect 204502 63349 204554 63355
rect 204596 63002 204652 63011
rect 204596 62937 204652 62946
rect 204610 60823 204638 62937
rect 204692 62410 204748 62419
rect 204692 62345 204748 62354
rect 204598 60817 204650 60823
rect 204500 60782 204556 60791
rect 204598 60759 204650 60765
rect 204706 60749 204734 62345
rect 204884 61818 204940 61827
rect 204884 61753 204940 61762
rect 204788 61374 204844 61383
rect 204788 61309 204844 61318
rect 204500 60717 204556 60726
rect 204694 60743 204746 60749
rect 204514 60675 204542 60717
rect 204694 60685 204746 60691
rect 204502 60669 204554 60675
rect 204502 60611 204554 60617
rect 204802 60527 204830 61309
rect 204898 60601 204926 61753
rect 204886 60595 204938 60601
rect 204886 60537 204938 60543
rect 204790 60521 204842 60527
rect 204790 60463 204842 60469
rect 206806 60447 206858 60453
rect 206806 60389 206858 60395
rect 204598 60373 204650 60379
rect 204598 60315 204650 60321
rect 204500 60190 204556 60199
rect 204500 60125 204556 60134
rect 204514 59047 204542 60125
rect 204610 59163 204638 60315
rect 206818 60051 206846 60389
rect 206804 60042 206860 60051
rect 206804 59977 206860 59986
rect 204596 59154 204652 59163
rect 204596 59089 204652 59098
rect 204502 59041 204554 59047
rect 204502 58983 204554 58989
rect 206900 55898 206956 55907
rect 206900 55833 206956 55842
rect 202966 47201 203018 47207
rect 202966 47143 203018 47149
rect 200086 47053 200138 47059
rect 200086 46995 200138 47001
rect 194326 46979 194378 46985
rect 194326 46921 194378 46927
rect 162646 46165 162698 46171
rect 162646 46107 162698 46113
rect 133654 42835 133706 42841
rect 133654 42777 133706 42783
rect 136534 42835 136586 42841
rect 136534 42777 136586 42783
rect 136546 40219 136574 42777
rect 206914 42175 206942 55833
rect 207106 53243 207134 229881
rect 207394 227471 207422 232101
rect 207956 230982 208012 230991
rect 207956 230917 208012 230926
rect 207382 227465 207434 227471
rect 207382 227407 207434 227413
rect 207190 213183 207242 213189
rect 207190 213125 207242 213131
rect 207202 210271 207230 213125
rect 207188 210262 207244 210271
rect 207188 210197 207244 210206
rect 207284 190134 207340 190143
rect 207284 190069 207340 190078
rect 207298 187215 207326 190069
rect 207286 187209 207338 187215
rect 207286 187151 207338 187157
rect 207382 162937 207434 162943
rect 207382 162879 207434 162885
rect 207394 112401 207422 162879
rect 207190 112395 207242 112401
rect 207190 112337 207242 112343
rect 207382 112395 207434 112401
rect 207382 112337 207434 112343
rect 207202 89239 207230 112337
rect 207190 89233 207242 89239
rect 207190 89175 207242 89181
rect 207286 69179 207338 69185
rect 207286 69121 207338 69127
rect 207298 64801 207326 69121
rect 207478 69031 207530 69037
rect 207478 68973 207530 68979
rect 207202 64773 207326 64801
rect 207202 53275 207230 64773
rect 207284 57674 207340 57683
rect 207284 57609 207340 57618
rect 207190 53269 207242 53275
rect 207092 53234 207148 53243
rect 207190 53211 207242 53217
rect 207092 53169 207148 53178
rect 207298 52905 207326 57609
rect 207490 54237 207518 68973
rect 207766 60373 207818 60379
rect 207766 60315 207818 60321
rect 207478 54231 207530 54237
rect 207478 54173 207530 54179
rect 207286 52899 207338 52905
rect 207286 52841 207338 52847
rect 207778 46319 207806 60315
rect 207862 60299 207914 60305
rect 207862 60241 207914 60247
rect 207874 46763 207902 60241
rect 207970 53053 207998 230917
rect 208066 53867 208094 233549
rect 209588 231574 209644 231583
rect 209588 231509 209644 231518
rect 209396 230538 209452 230547
rect 209396 230473 209452 230482
rect 209300 202714 209356 202723
rect 209300 202649 209356 202658
rect 208726 164195 208778 164201
rect 208726 164137 208778 164143
rect 208630 126751 208682 126757
rect 208630 126693 208682 126699
rect 208534 121053 208586 121059
rect 208534 120995 208586 121001
rect 208438 118167 208490 118173
rect 208438 118109 208490 118115
rect 208342 115281 208394 115287
rect 208342 115223 208394 115229
rect 208246 103737 208298 103743
rect 208246 103679 208298 103685
rect 208150 97965 208202 97971
rect 208150 97907 208202 97913
rect 208054 53861 208106 53867
rect 208054 53803 208106 53809
rect 208162 53127 208190 97907
rect 208150 53121 208202 53127
rect 208150 53063 208202 53069
rect 207958 53047 208010 53053
rect 207958 52989 208010 52995
rect 208258 50389 208286 103679
rect 208150 50383 208202 50389
rect 208150 50325 208202 50331
rect 208246 50383 208298 50389
rect 208246 50325 208298 50331
rect 207958 50309 208010 50315
rect 207958 50251 208010 50257
rect 207970 49723 207998 50251
rect 208162 49797 208190 50325
rect 208150 49791 208202 49797
rect 208150 49733 208202 49739
rect 207958 49717 208010 49723
rect 207958 49659 208010 49665
rect 208354 49649 208382 115223
rect 208450 53941 208478 118109
rect 208438 53935 208490 53941
rect 208438 53877 208490 53883
rect 208342 49643 208394 49649
rect 208342 49585 208394 49591
rect 208546 48909 208574 120995
rect 208534 48903 208586 48909
rect 208534 48845 208586 48851
rect 208642 48761 208670 126693
rect 208738 60379 208766 164137
rect 208822 144067 208874 144073
rect 208822 144009 208874 144015
rect 208726 60373 208778 60379
rect 208726 60315 208778 60321
rect 208834 60305 208862 144009
rect 208918 138295 208970 138301
rect 208918 138237 208970 138243
rect 208822 60299 208874 60305
rect 208822 60241 208874 60247
rect 208930 60176 208958 138237
rect 209110 132745 209162 132751
rect 209110 132687 209162 132693
rect 209014 132597 209066 132603
rect 209014 132539 209066 132545
rect 208738 60148 208958 60176
rect 208630 48755 208682 48761
rect 208630 48697 208682 48703
rect 208738 48391 208766 60148
rect 208822 60003 208874 60009
rect 208822 59945 208874 59951
rect 208834 48539 208862 59945
rect 209026 57660 209054 132539
rect 209122 60009 209150 132687
rect 209206 129637 209258 129643
rect 209206 129579 209258 129585
rect 209110 60003 209162 60009
rect 209110 59945 209162 59951
rect 208930 57632 209054 57660
rect 208930 48687 208958 57632
rect 209218 57512 209246 129579
rect 209026 57484 209246 57512
rect 209026 48835 209054 57484
rect 209314 57364 209342 202649
rect 209122 57336 209342 57364
rect 209122 49871 209150 57336
rect 209204 57230 209260 57239
rect 209204 57165 209260 57174
rect 209218 54089 209246 57165
rect 209300 56638 209356 56647
rect 209300 56573 209356 56582
rect 209206 54083 209258 54089
rect 209206 54025 209258 54031
rect 209314 54015 209342 56573
rect 209302 54009 209354 54015
rect 209302 53951 209354 53957
rect 209410 53349 209438 230473
rect 209494 60003 209546 60009
rect 209494 59945 209546 59951
rect 209398 53343 209450 53349
rect 209398 53285 209450 53291
rect 209110 49865 209162 49871
rect 209110 49807 209162 49813
rect 209506 48951 209534 59945
rect 209602 53423 209630 231509
rect 209590 53417 209642 53423
rect 209590 53359 209642 53365
rect 209698 51795 209726 236541
rect 209794 53201 209822 236689
rect 209782 53195 209834 53201
rect 209782 53137 209834 53143
rect 209686 51789 209738 51795
rect 209686 51731 209738 51737
rect 209890 51721 209918 239057
rect 210658 236203 210686 252049
rect 211126 246705 211178 246711
rect 211126 246647 211178 246653
rect 211030 246631 211082 246637
rect 211030 246573 211082 246579
rect 210742 246409 210794 246415
rect 210742 246351 210794 246357
rect 210754 245643 210782 246351
rect 211042 245939 211070 246573
rect 211138 246087 211166 246647
rect 211412 246374 211468 246383
rect 211318 246335 211370 246341
rect 211412 246309 211468 246318
rect 211318 246277 211370 246283
rect 211330 246235 211358 246277
rect 211316 246226 211372 246235
rect 211316 246161 211372 246170
rect 211124 246078 211180 246087
rect 211124 246013 211180 246022
rect 211028 245930 211084 245939
rect 211028 245865 211084 245874
rect 210740 245634 210796 245643
rect 210740 245569 210796 245578
rect 211426 244755 211454 246309
rect 211220 244746 211276 244755
rect 211412 244746 211468 244755
rect 211276 244704 211358 244732
rect 211220 244681 211276 244690
rect 211030 239009 211082 239015
rect 211030 238951 211082 238957
rect 210932 236310 210988 236319
rect 210932 236245 210988 236254
rect 210262 236197 210314 236203
rect 210262 236139 210314 236145
rect 210646 236197 210698 236203
rect 210646 236139 210698 236145
rect 210164 234830 210220 234839
rect 210164 234765 210220 234774
rect 210070 233533 210122 233539
rect 210070 233475 210122 233481
rect 209974 233459 210026 233465
rect 209974 233401 210026 233407
rect 209986 60009 210014 233401
rect 209974 60003 210026 60009
rect 209974 59945 210026 59951
rect 209972 56046 210028 56055
rect 209972 55981 210028 55990
rect 209986 54903 210014 55981
rect 209974 54897 210026 54903
rect 209974 54839 210026 54845
rect 209972 54788 210028 54797
rect 209972 54723 210028 54732
rect 209986 53645 210014 54723
rect 210082 54163 210110 233475
rect 210178 228919 210206 234765
rect 210164 228910 210220 228919
rect 210164 228845 210220 228854
rect 210164 172670 210220 172679
rect 210164 172605 210220 172614
rect 210178 152699 210206 172605
rect 210164 152690 210220 152699
rect 210164 152625 210220 152634
rect 210164 119094 210220 119103
rect 210164 119029 210220 119038
rect 210178 94239 210206 119029
rect 210164 94230 210220 94239
rect 210164 94165 210220 94174
rect 210166 80353 210218 80359
rect 210166 80295 210218 80301
rect 210178 78181 210206 80295
rect 210164 78172 210220 78181
rect 210164 78107 210220 78116
rect 210274 55144 210302 236139
rect 210358 233681 210410 233687
rect 210358 233623 210410 233629
rect 210178 55116 210302 55144
rect 210178 54311 210206 55116
rect 210260 55010 210316 55019
rect 210260 54945 210316 54954
rect 210166 54305 210218 54311
rect 210166 54247 210218 54253
rect 210070 54157 210122 54163
rect 210070 54099 210122 54105
rect 210274 53719 210302 54945
rect 210262 53713 210314 53719
rect 210262 53655 210314 53661
rect 209974 53639 210026 53645
rect 209974 53581 210026 53587
rect 210370 53497 210398 233623
rect 210946 233484 210974 236245
rect 211042 233655 211070 238951
rect 211330 233655 211358 244704
rect 211412 244681 211468 244690
rect 211522 244195 211550 261839
rect 211618 247377 211646 273509
rect 212564 273458 212620 273467
rect 212564 273393 212620 273402
rect 212374 273271 212426 273277
rect 212374 273213 212426 273219
rect 212182 271495 212234 271501
rect 212182 271437 212234 271443
rect 211796 271386 211852 271395
rect 211796 271321 211852 271330
rect 211702 271199 211754 271205
rect 211702 271141 211754 271147
rect 211606 247371 211658 247377
rect 211606 247313 211658 247319
rect 211714 247100 211742 271141
rect 211810 247303 211838 271321
rect 211894 271273 211946 271279
rect 211894 271215 211946 271221
rect 211988 271238 212044 271247
rect 211798 247297 211850 247303
rect 211798 247239 211850 247245
rect 211714 247072 211838 247100
rect 211606 246853 211658 246859
rect 211606 246795 211658 246801
rect 211618 246679 211646 246795
rect 211604 246670 211660 246679
rect 211604 246605 211660 246614
rect 211810 245231 211838 247072
rect 211906 246360 211934 271215
rect 211988 271173 212044 271182
rect 212002 247155 212030 271173
rect 212086 271125 212138 271131
rect 212086 271067 212138 271073
rect 211990 247149 212042 247155
rect 211990 247091 212042 247097
rect 211906 246332 212030 246360
rect 211894 246261 211946 246267
rect 211894 246203 211946 246209
rect 211798 245225 211850 245231
rect 211798 245167 211850 245173
rect 211510 244189 211562 244195
rect 211510 244131 211562 244137
rect 211906 233803 211934 246203
rect 212002 245157 212030 246332
rect 211990 245151 212042 245157
rect 211990 245093 212042 245099
rect 212098 244607 212126 271067
rect 212194 247229 212222 271437
rect 212386 265142 212414 273213
rect 212578 270803 212606 273393
rect 213346 273277 213374 277870
rect 214594 274091 214622 277870
rect 214582 274085 214634 274091
rect 214582 274027 214634 274033
rect 213334 273271 213386 273277
rect 213334 273213 213386 273219
rect 213044 272866 213100 272875
rect 213044 272801 213100 272810
rect 213058 271131 213086 272801
rect 213238 271865 213290 271871
rect 213238 271807 213290 271813
rect 213046 271125 213098 271131
rect 213046 271067 213098 271073
rect 212564 270794 212620 270803
rect 212564 270729 212620 270738
rect 212756 270794 212812 270803
rect 212756 270729 212812 270738
rect 212770 265142 212798 270729
rect 213250 265142 213278 271807
rect 213814 271051 213866 271057
rect 213814 270993 213866 270999
rect 213826 265156 213854 270993
rect 214486 270977 214538 270983
rect 214486 270919 214538 270925
rect 213826 265128 214080 265156
rect 214498 265142 214526 270919
rect 214966 270903 215018 270909
rect 214966 270845 215018 270851
rect 214978 265142 215006 270845
rect 215446 270829 215498 270835
rect 215446 270771 215498 270777
rect 215458 265142 215486 270771
rect 215542 270755 215594 270761
rect 215542 270697 215594 270703
rect 215554 265156 215582 270697
rect 215746 266543 215774 277870
rect 216118 273493 216170 273499
rect 216118 273435 216170 273441
rect 216022 269941 216074 269947
rect 216020 269906 216022 269915
rect 216074 269906 216076 269915
rect 216020 269841 216076 269850
rect 215734 266537 215786 266543
rect 215734 266479 215786 266485
rect 216130 265156 216158 273435
rect 216694 273271 216746 273277
rect 216694 273213 216746 273219
rect 215554 265128 215808 265156
rect 216130 265128 216288 265156
rect 216706 265142 216734 273213
rect 216898 265156 216926 277870
rect 217364 273310 217420 273319
rect 217364 273245 217420 273254
rect 217558 273271 217610 273277
rect 217378 270951 217406 273245
rect 217558 273213 217610 273219
rect 217364 270942 217420 270951
rect 217364 270877 217420 270886
rect 216898 265128 217200 265156
rect 217570 265142 217598 273213
rect 218050 268319 218078 277870
rect 218230 273493 218282 273499
rect 218230 273435 218282 273441
rect 218038 268313 218090 268319
rect 218038 268255 218090 268261
rect 218242 265156 218270 273435
rect 220450 273277 220478 277870
rect 220438 273271 220490 273277
rect 220438 273213 220490 273219
rect 220822 271791 220874 271797
rect 220822 271733 220874 271739
rect 220342 271273 220394 271279
rect 220342 271215 220394 271221
rect 219766 271199 219818 271205
rect 219766 271141 219818 271147
rect 219286 271125 219338 271131
rect 219286 271067 219338 271073
rect 218902 271051 218954 271057
rect 218902 270993 218954 270999
rect 218710 270977 218762 270983
rect 218710 270919 218762 270925
rect 218722 265156 218750 270919
rect 218016 265128 218270 265156
rect 218496 265128 218750 265156
rect 218914 265142 218942 270993
rect 219298 265142 219326 271067
rect 219778 265142 219806 271141
rect 220354 265156 220382 271215
rect 220834 265156 220862 271733
rect 221014 270903 221066 270909
rect 221014 270845 221066 270851
rect 220224 265128 220382 265156
rect 220608 265128 220862 265156
rect 221026 265142 221054 270845
rect 221494 269275 221546 269281
rect 221494 269217 221546 269223
rect 221506 265142 221534 269217
rect 221698 265211 221726 277870
rect 222864 277856 223166 277884
rect 223030 273789 223082 273795
rect 223030 273731 223082 273737
rect 222550 268017 222602 268023
rect 222550 267959 222602 267965
rect 221974 267869 222026 267875
rect 221974 267811 222026 267817
rect 221686 265205 221738 265211
rect 221686 265147 221738 265153
rect 221986 265142 222014 267811
rect 222562 265156 222590 267959
rect 223042 265156 223070 273731
rect 222336 265128 222590 265156
rect 222816 265128 223070 265156
rect 223138 265137 223166 277856
rect 224002 273499 224030 277870
rect 225264 277856 225374 277884
rect 225238 273937 225290 273943
rect 225238 273879 225290 273885
rect 224086 273863 224138 273869
rect 224086 273805 224138 273811
rect 223990 273493 224042 273499
rect 223990 273435 224042 273441
rect 223702 268239 223754 268245
rect 223702 268181 223754 268187
rect 223222 268165 223274 268171
rect 223222 268107 223274 268113
rect 223234 265142 223262 268107
rect 223714 265142 223742 268181
rect 224098 265142 224126 273805
rect 224566 273493 224618 273499
rect 224566 273435 224618 273441
rect 224578 265156 224606 273435
rect 225250 265156 225278 273879
rect 225346 265285 225374 277856
rect 226294 275565 226346 275571
rect 226294 275507 226346 275513
rect 225430 274011 225482 274017
rect 225430 273953 225482 273959
rect 225334 265279 225386 265285
rect 225334 265221 225386 265227
rect 223126 265131 223178 265137
rect 224544 265128 224606 265156
rect 225024 265128 225278 265156
rect 225442 265142 225470 273953
rect 225814 268461 225866 268467
rect 225814 268403 225866 268409
rect 225826 265142 225854 268403
rect 226306 265142 226334 275507
rect 227446 275491 227498 275497
rect 227446 275433 227498 275439
rect 226966 269867 227018 269873
rect 226966 269809 227018 269815
rect 226978 265156 227006 269809
rect 227458 265156 227486 275433
rect 227540 271682 227596 271691
rect 227540 271617 227596 271626
rect 227554 271099 227582 271617
rect 227540 271090 227596 271099
rect 227540 271025 227596 271034
rect 227650 270983 227678 277870
rect 228022 275195 228074 275201
rect 228022 275137 228074 275143
rect 227638 270977 227690 270983
rect 227638 270919 227690 270925
rect 227542 269571 227594 269577
rect 227542 269513 227594 269519
rect 226752 265128 227006 265156
rect 227232 265128 227486 265156
rect 227554 265142 227582 269513
rect 228034 265142 228062 275137
rect 228802 273573 228830 277870
rect 229078 275047 229130 275053
rect 229078 274989 229130 274995
rect 228790 273567 228842 273573
rect 228790 273509 228842 273515
rect 228502 269423 228554 269429
rect 228502 269365 228554 269371
rect 228514 265142 228542 269365
rect 229090 265156 229118 274989
rect 229750 273271 229802 273277
rect 229750 273213 229802 273219
rect 229558 269349 229610 269355
rect 229558 269291 229610 269297
rect 229570 265156 229598 269291
rect 228864 265128 229118 265156
rect 229344 265128 229598 265156
rect 229762 265142 229790 273213
rect 230050 266691 230078 277870
rect 230230 274307 230282 274313
rect 230230 274249 230282 274255
rect 230038 266685 230090 266691
rect 230038 266627 230090 266633
rect 230242 265142 230270 274249
rect 230614 274233 230666 274239
rect 230614 274175 230666 274181
rect 230626 265142 230654 274175
rect 231202 271057 231230 277870
rect 231766 276453 231818 276459
rect 231766 276395 231818 276401
rect 231190 271051 231242 271057
rect 231190 270993 231242 270999
rect 231286 270681 231338 270687
rect 231286 270623 231338 270629
rect 231298 265156 231326 270623
rect 231778 265156 231806 276395
rect 232342 276379 232394 276385
rect 232342 276321 232394 276327
rect 231958 270533 232010 270539
rect 231958 270475 232010 270481
rect 231072 265128 231326 265156
rect 231552 265128 231806 265156
rect 231970 265142 231998 270475
rect 232354 265142 232382 276321
rect 232450 271871 232478 277870
rect 233398 276157 233450 276163
rect 233398 276099 233450 276105
rect 232438 271865 232490 271871
rect 232438 271807 232490 271813
rect 232822 270385 232874 270391
rect 232822 270327 232874 270333
rect 232834 265142 232862 270327
rect 233410 265156 233438 276099
rect 233506 274831 233534 277870
rect 234070 276009 234122 276015
rect 234070 275951 234122 275957
rect 233494 274825 233546 274831
rect 233494 274767 233546 274773
rect 233974 270311 234026 270317
rect 233974 270253 234026 270259
rect 233986 265156 234014 270253
rect 233280 265128 233438 265156
rect 233760 265128 234014 265156
rect 234082 265142 234110 275951
rect 234658 271131 234686 277870
rect 235030 275713 235082 275719
rect 235030 275655 235082 275661
rect 234646 271125 234698 271131
rect 234646 271067 234698 271073
rect 234550 270163 234602 270169
rect 234550 270105 234602 270111
rect 234562 265142 234590 270105
rect 235042 265142 235070 275655
rect 235702 270089 235754 270095
rect 235702 270031 235754 270037
rect 235714 265156 235742 270031
rect 235906 268097 235934 277870
rect 237168 277856 237470 277884
rect 235990 275639 236042 275645
rect 235990 275581 236042 275587
rect 235894 268091 235946 268097
rect 235894 268033 235946 268039
rect 236002 265156 236030 275581
rect 236758 275343 236810 275349
rect 236758 275285 236810 275291
rect 236278 269497 236330 269503
rect 236278 269439 236330 269445
rect 235488 265128 235742 265156
rect 235872 265128 236030 265156
rect 236290 265142 236318 269439
rect 236770 265142 236798 275285
rect 237142 268905 237194 268911
rect 237142 268847 237194 268853
rect 237154 265142 237182 268847
rect 237442 266987 237470 277856
rect 237814 274381 237866 274387
rect 237814 274323 237866 274329
rect 237620 273458 237676 273467
rect 237620 273393 237676 273402
rect 237524 272866 237580 272875
rect 237524 272801 237580 272810
rect 237538 271395 237566 272801
rect 237524 271386 237580 271395
rect 237524 271321 237580 271330
rect 237634 271247 237662 273393
rect 237716 273310 237772 273319
rect 237716 273245 237772 273254
rect 237730 271395 237758 273245
rect 237716 271386 237772 271395
rect 237716 271321 237772 271330
rect 237620 271238 237676 271247
rect 237620 271173 237676 271182
rect 237430 266981 237482 266987
rect 237430 266923 237482 266929
rect 237826 265156 237854 274323
rect 238306 271205 238334 277870
rect 239458 276681 239486 277870
rect 240706 277347 240734 277870
rect 240694 277341 240746 277347
rect 240694 277283 240746 277289
rect 239446 276675 239498 276681
rect 239446 276617 239498 276623
rect 241078 274677 241130 274683
rect 241078 274619 241130 274625
rect 240502 274603 240554 274609
rect 240502 274545 240554 274551
rect 239350 274529 239402 274535
rect 239350 274471 239402 274477
rect 238486 274455 238538 274461
rect 238486 274397 238538 274403
rect 238294 271199 238346 271205
rect 238294 271141 238346 271147
rect 238294 268683 238346 268689
rect 238294 268625 238346 268631
rect 238306 265156 238334 268625
rect 237600 265128 237854 265156
rect 238080 265128 238334 265156
rect 238498 265142 238526 274397
rect 238870 268609 238922 268615
rect 238870 268551 238922 268557
rect 238882 265142 238910 268551
rect 239362 265142 239390 274471
rect 240022 268535 240074 268541
rect 240022 268477 240074 268483
rect 240034 265156 240062 268477
rect 240514 265156 240542 274545
rect 240886 268757 240938 268763
rect 240886 268699 240938 268705
rect 240898 265156 240926 268699
rect 239808 265128 240062 265156
rect 240288 265128 240542 265156
rect 240672 265128 240926 265156
rect 241090 265142 241118 274619
rect 241858 271279 241886 277870
rect 242998 274899 243050 274905
rect 242998 274841 243050 274847
rect 242230 274751 242282 274757
rect 242230 274693 242282 274699
rect 241846 271273 241898 271279
rect 241846 271215 241898 271221
rect 241558 268831 241610 268837
rect 241558 268773 241610 268779
rect 241570 265142 241598 268773
rect 242242 265156 242270 274693
rect 242614 268979 242666 268985
rect 242614 268921 242666 268927
rect 242626 265156 242654 268921
rect 243010 265156 243038 274841
rect 243106 267949 243134 277870
rect 243766 274973 243818 274979
rect 243766 274915 243818 274921
rect 243286 269941 243338 269947
rect 243284 269906 243286 269915
rect 243338 269906 243340 269915
rect 243284 269841 243340 269850
rect 243286 269053 243338 269059
rect 243286 268995 243338 269001
rect 243094 267943 243146 267949
rect 243094 267885 243146 267891
rect 242016 265128 242270 265156
rect 242400 265128 242654 265156
rect 242880 265128 243038 265156
rect 243298 265142 243326 268995
rect 243778 265142 243806 274915
rect 244150 269201 244202 269207
rect 244150 269143 244202 269149
rect 244162 265142 244190 269143
rect 244258 267061 244286 277870
rect 244726 276305 244778 276311
rect 244726 276247 244778 276253
rect 244246 267055 244298 267061
rect 244246 266997 244298 267003
rect 244738 265156 244766 276247
rect 245398 276231 245450 276237
rect 245398 276173 245450 276179
rect 245302 270607 245354 270613
rect 245302 270549 245354 270555
rect 245314 265156 245342 270549
rect 244608 265128 244766 265156
rect 245088 265128 245342 265156
rect 245410 265142 245438 276173
rect 245506 271797 245534 277870
rect 246358 276083 246410 276089
rect 246358 276025 246410 276031
rect 245494 271791 245546 271797
rect 245494 271733 245546 271739
rect 245878 270459 245930 270465
rect 245878 270401 245930 270407
rect 245890 265142 245918 270401
rect 246370 265142 246398 276025
rect 246658 271501 246686 277870
rect 247906 276755 247934 277870
rect 247894 276749 247946 276755
rect 247894 276691 247946 276697
rect 247414 275935 247466 275941
rect 247414 275877 247466 275883
rect 246646 271495 246698 271501
rect 246646 271437 246698 271443
rect 247030 270237 247082 270243
rect 247030 270179 247082 270185
rect 247042 265156 247070 270179
rect 247426 265156 247454 275877
rect 248086 275787 248138 275793
rect 248086 275729 248138 275735
rect 247604 271682 247660 271691
rect 247604 271617 247660 271626
rect 247618 271099 247646 271617
rect 247604 271090 247660 271099
rect 247604 271025 247660 271034
rect 247606 270015 247658 270021
rect 247606 269957 247658 269963
rect 246816 265128 247070 265156
rect 247200 265128 247454 265156
rect 247618 265142 247646 269957
rect 248098 265142 248126 275729
rect 248180 273606 248236 273615
rect 248180 273541 248236 273550
rect 248194 272727 248222 273541
rect 248180 272718 248236 272727
rect 248180 272653 248236 272662
rect 249058 270909 249086 277870
rect 249812 274050 249868 274059
rect 249812 273985 249868 273994
rect 249140 273902 249196 273911
rect 249140 273837 249196 273846
rect 249046 270903 249098 270909
rect 249046 270845 249098 270851
rect 248566 269941 248618 269947
rect 248566 269883 248618 269889
rect 248578 265142 248606 269883
rect 249154 265156 249182 273837
rect 249622 269793 249674 269799
rect 249622 269735 249674 269741
rect 249634 265156 249662 269735
rect 248928 265128 249182 265156
rect 249408 265128 249662 265156
rect 249826 265142 249854 273985
rect 250210 271797 250238 277870
rect 251376 277856 251678 277884
rect 250676 274198 250732 274207
rect 250676 274133 250732 274142
rect 250580 273310 250636 273319
rect 250580 273245 250636 273254
rect 250198 271791 250250 271797
rect 250198 271733 250250 271739
rect 250594 271395 250622 273245
rect 250580 271386 250636 271395
rect 250580 271321 250636 271330
rect 250294 269719 250346 269725
rect 250294 269661 250346 269667
rect 250306 265142 250334 269661
rect 250690 265142 250718 274133
rect 251350 269645 251402 269651
rect 251350 269587 251402 269593
rect 251362 265156 251390 269587
rect 251650 267209 251678 277856
rect 252310 276675 252362 276681
rect 252310 276617 252362 276623
rect 251828 274346 251884 274355
rect 251828 274281 251884 274290
rect 251638 267203 251690 267209
rect 251638 267145 251690 267151
rect 251842 265156 251870 274281
rect 252322 274091 252350 276617
rect 252404 274494 252460 274503
rect 252404 274429 252460 274438
rect 252214 274085 252266 274091
rect 252214 274027 252266 274033
rect 252310 274085 252362 274091
rect 252310 274027 252362 274033
rect 252226 273795 252254 274027
rect 252214 273789 252266 273795
rect 252214 273731 252266 273737
rect 252020 268870 252076 268879
rect 252020 268805 252076 268814
rect 251136 265128 251390 265156
rect 251616 265128 251870 265156
rect 252034 265142 252062 268805
rect 252418 265142 252446 274429
rect 252514 269281 252542 277870
rect 253762 271057 253790 277870
rect 254914 277051 254942 277870
rect 254902 277045 254954 277051
rect 254902 276987 254954 276993
rect 253940 274642 253996 274651
rect 253940 274577 253996 274586
rect 253750 271051 253802 271057
rect 253750 270993 253802 270999
rect 253462 270903 253514 270909
rect 253462 270845 253514 270851
rect 253364 269906 253420 269915
rect 253364 269841 253420 269850
rect 253378 269767 253406 269841
rect 253364 269758 253420 269767
rect 253364 269693 253420 269702
rect 252502 269275 252554 269281
rect 252502 269217 252554 269223
rect 253364 269166 253420 269175
rect 253364 269101 253420 269110
rect 252884 269018 252940 269027
rect 252884 268953 252940 268962
rect 252898 265142 252926 268953
rect 253378 265156 253406 269101
rect 253474 268023 253502 270845
rect 253462 268017 253514 268023
rect 253462 267959 253514 267965
rect 253954 265156 253982 274577
rect 255092 273754 255148 273763
rect 255092 273689 255148 273698
rect 254612 270350 254668 270359
rect 254612 270285 254668 270294
rect 254134 269275 254186 269281
rect 254134 269217 254186 269223
rect 253344 265128 253406 265156
rect 253728 265128 253982 265156
rect 254146 265142 254174 269217
rect 254626 265142 254654 270285
rect 255106 265142 255134 273689
rect 256162 267875 256190 277870
rect 257314 270835 257342 277870
rect 258576 277856 258878 277884
rect 257506 275340 257918 275368
rect 257506 275201 257534 275340
rect 257590 275269 257642 275275
rect 257642 275217 257822 275220
rect 257590 275211 257822 275217
rect 257494 275195 257546 275201
rect 257602 275192 257822 275211
rect 257890 275201 257918 275340
rect 257494 275137 257546 275143
rect 257794 275127 257822 275192
rect 257878 275195 257930 275201
rect 257878 275137 257930 275143
rect 257590 275121 257642 275127
rect 257590 275063 257642 275069
rect 257782 275121 257834 275127
rect 257782 275063 257834 275069
rect 257302 270829 257354 270835
rect 257302 270771 257354 270777
rect 256436 270646 256492 270655
rect 256436 270581 256492 270590
rect 256340 269462 256396 269471
rect 256450 269448 256478 270581
rect 256396 269420 256478 269448
rect 256340 269397 256396 269406
rect 256150 267869 256202 267875
rect 256150 267811 256202 267817
rect 255670 267721 255722 267727
rect 255670 267663 255722 267669
rect 256148 267686 256204 267695
rect 255682 265156 255710 267663
rect 256148 267621 256204 267630
rect 256162 265156 256190 267621
rect 256340 267390 256396 267399
rect 256340 267325 256396 267334
rect 255456 265128 255710 265156
rect 255936 265128 256190 265156
rect 256354 265142 256382 267325
rect 256820 267242 256876 267251
rect 256820 267177 256876 267186
rect 256834 265142 256862 267177
rect 257204 267094 257260 267103
rect 257204 267029 257260 267038
rect 257218 265142 257246 267029
rect 257602 265581 257630 275063
rect 257684 273458 257740 273467
rect 257684 273393 257740 273402
rect 257698 271247 257726 273393
rect 257684 271238 257740 271247
rect 257684 271173 257740 271182
rect 257876 270498 257932 270507
rect 257876 270433 257932 270442
rect 257590 265575 257642 265581
rect 257590 265517 257642 265523
rect 257890 265156 257918 270433
rect 258548 268574 258604 268583
rect 258548 268509 258604 268518
rect 258356 267982 258412 267991
rect 258356 267917 258412 267926
rect 258370 265156 258398 267917
rect 257664 265128 257918 265156
rect 258144 265128 258398 265156
rect 258562 265142 258590 268509
rect 258850 267357 258878 277856
rect 259412 274790 259468 274799
rect 259412 274725 259468 274734
rect 258932 268130 258988 268139
rect 258932 268065 258988 268074
rect 258838 267351 258890 267357
rect 258838 267293 258890 267299
rect 258946 265142 258974 268065
rect 259426 265142 259454 274725
rect 259714 270909 259742 277870
rect 260084 272866 260140 272875
rect 260084 272801 260140 272810
rect 259702 270903 259754 270909
rect 259702 270845 259754 270851
rect 260098 265156 260126 272801
rect 260962 270909 260990 277870
rect 262114 276829 262142 277870
rect 262102 276823 262154 276829
rect 262102 276765 262154 276771
rect 262676 276418 262732 276427
rect 262676 276353 262732 276362
rect 262004 274938 262060 274947
rect 262004 274873 262060 274882
rect 261140 271090 261196 271099
rect 261140 271025 261196 271034
rect 260950 270903 261002 270909
rect 260950 270845 261002 270851
rect 260564 269610 260620 269619
rect 260564 269545 260620 269554
rect 260578 265156 260606 269545
rect 260660 268278 260716 268287
rect 260660 268213 260716 268222
rect 259872 265128 260126 265156
rect 260352 265128 260606 265156
rect 260674 265142 260702 268213
rect 261154 265142 261182 271025
rect 261620 269314 261676 269323
rect 261620 269249 261676 269258
rect 261634 265142 261662 269249
rect 262018 265156 262046 274873
rect 262690 265156 262718 276353
rect 262868 276122 262924 276131
rect 262868 276057 262924 276066
rect 261984 265128 262046 265156
rect 262464 265128 262718 265156
rect 262882 265142 262910 276057
rect 263362 273721 263390 277870
rect 263636 275974 263692 275983
rect 263636 275909 263692 275918
rect 263350 273715 263402 273721
rect 263350 273657 263402 273663
rect 263650 265156 263678 275909
rect 263732 275826 263788 275835
rect 263732 275761 263788 275770
rect 263376 265128 263678 265156
rect 263746 265142 263774 275761
rect 264404 275678 264460 275687
rect 264404 275613 264460 275622
rect 264418 265156 264446 275613
rect 264514 271131 264542 277870
rect 265460 275530 265516 275539
rect 265460 275465 265516 275474
rect 264502 271125 264554 271131
rect 264502 271067 264554 271073
rect 264884 270942 264940 270951
rect 264884 270877 264940 270886
rect 264898 265156 264926 270877
rect 265076 268426 265132 268435
rect 265076 268361 265132 268370
rect 264192 265128 264446 265156
rect 264672 265128 264926 265156
rect 265090 265142 265118 268361
rect 265474 265142 265502 275465
rect 265762 267505 265790 277870
rect 266530 277856 266832 277884
rect 265940 275234 265996 275243
rect 265940 275169 265996 275178
rect 265750 267499 265802 267505
rect 265750 267441 265802 267447
rect 265954 265142 265982 275169
rect 266530 268171 266558 277856
rect 267670 275417 267722 275423
rect 267668 275382 267670 275391
rect 267766 275417 267818 275423
rect 267722 275382 267724 275391
rect 267766 275359 267818 275365
rect 267860 275382 267916 275391
rect 267668 275317 267724 275326
rect 267778 275220 267806 275359
rect 267860 275317 267916 275326
rect 267682 275192 267806 275220
rect 267682 275127 267710 275192
rect 267670 275121 267722 275127
rect 266900 275086 266956 275095
rect 267670 275063 267722 275069
rect 267766 275121 267818 275127
rect 267766 275063 267818 275069
rect 266900 275021 266956 275030
rect 266518 268165 266570 268171
rect 266518 268107 266570 268113
rect 266614 267943 266666 267949
rect 266614 267885 266666 267891
rect 266626 265156 266654 267885
rect 266914 265452 266942 275021
rect 267778 273795 267806 275063
rect 267766 273789 267818 273795
rect 267766 273731 267818 273737
rect 267190 273715 267242 273721
rect 267190 273657 267242 273663
rect 266400 265128 266654 265156
rect 266866 265424 266942 265452
rect 266866 265142 266894 265424
rect 267202 265142 267230 273657
rect 267874 273647 267902 275317
rect 267862 273641 267914 273647
rect 267862 273583 267914 273589
rect 268066 271797 268094 277870
rect 269218 276903 269246 277870
rect 269206 276897 269258 276903
rect 269206 276839 269258 276845
rect 268148 275678 268204 275687
rect 268148 275613 268204 275622
rect 268162 275516 268190 275613
rect 268820 275530 268876 275539
rect 268162 275488 268820 275516
rect 268820 275465 268876 275474
rect 270262 275417 270314 275423
rect 270262 275359 270314 275365
rect 269398 273789 269450 273795
rect 269398 273731 269450 273737
rect 267958 271791 268010 271797
rect 267958 271733 268010 271739
rect 268054 271791 268106 271797
rect 268054 271733 268106 271739
rect 267860 271682 267916 271691
rect 267860 271617 267916 271626
rect 267874 271395 267902 271617
rect 267860 271386 267916 271395
rect 267860 271321 267916 271330
rect 267970 271205 267998 271733
rect 267958 271199 268010 271205
rect 267958 271141 268010 271147
rect 268726 270977 268778 270983
rect 268726 270919 268778 270925
rect 268148 269462 268204 269471
rect 268148 269397 268204 269406
rect 267670 267869 267722 267875
rect 267670 267811 267722 267817
rect 267572 267390 267628 267399
rect 267572 267325 267628 267334
rect 267586 267283 267614 267325
rect 267574 267277 267626 267283
rect 267574 267219 267626 267225
rect 267682 265142 267710 267811
rect 267766 267721 267818 267727
rect 267764 267686 267766 267695
rect 267818 267686 267820 267695
rect 267764 267621 267820 267630
rect 267862 267573 267914 267579
rect 267860 267538 267862 267547
rect 267914 267538 267916 267547
rect 267860 267473 267916 267482
rect 268052 267538 268108 267547
rect 268052 267473 268108 267482
rect 268066 267283 268094 267473
rect 268054 267277 268106 267283
rect 268054 267219 268106 267225
rect 268162 265142 268190 269397
rect 268738 265156 268766 270919
rect 269204 268722 269260 268731
rect 269204 268657 269260 268666
rect 269218 265156 269246 268657
rect 268512 265128 268766 265156
rect 268992 265128 269246 265156
rect 269410 265142 269438 273731
rect 269878 265575 269930 265581
rect 269878 265517 269930 265523
rect 269890 265142 269918 265517
rect 270274 265142 270302 275359
rect 270370 268245 270398 277870
rect 271318 274159 271370 274165
rect 271318 274101 271370 274107
rect 270562 273712 270878 273740
rect 270562 270983 270590 273712
rect 270850 273647 270878 273712
rect 270742 273641 270794 273647
rect 270742 273583 270794 273589
rect 270838 273641 270890 273647
rect 270838 273583 270890 273589
rect 270644 271534 270700 271543
rect 270644 271469 270700 271478
rect 270550 270977 270602 270983
rect 270550 270919 270602 270925
rect 270358 268239 270410 268245
rect 270358 268181 270410 268187
rect 270658 266469 270686 271469
rect 270646 266463 270698 266469
rect 270646 266405 270698 266411
rect 270754 265156 270782 273583
rect 271222 271865 271274 271871
rect 271222 271807 271274 271813
rect 271234 271279 271262 271807
rect 271222 271273 271274 271279
rect 271222 271215 271274 271221
rect 270934 269127 270986 269133
rect 270934 269069 270986 269075
rect 270720 265128 270782 265156
rect 270946 265156 270974 269069
rect 271330 265156 271358 274101
rect 271618 271871 271646 277870
rect 272470 275121 272522 275127
rect 272470 275063 272522 275069
rect 271606 271865 271658 271871
rect 271606 271807 271658 271813
rect 271990 268387 272042 268393
rect 271990 268329 272042 268335
rect 270946 265128 271200 265156
rect 271330 265128 271632 265156
rect 272002 265142 272030 268329
rect 272482 265142 272510 275063
rect 272770 269133 272798 277870
rect 274018 273869 274046 277870
rect 274006 273863 274058 273869
rect 274006 273805 274058 273811
rect 274102 273863 274154 273869
rect 274102 273805 274154 273811
rect 274114 273647 274142 273805
rect 274102 273641 274154 273647
rect 274102 273583 274154 273589
rect 275170 273573 275198 277870
rect 276418 274165 276446 277870
rect 276406 274159 276458 274165
rect 276406 274101 276458 274107
rect 275254 274085 275306 274091
rect 275254 274027 275306 274033
rect 274198 273567 274250 273573
rect 274198 273509 274250 273515
rect 275158 273567 275210 273573
rect 275158 273509 275210 273515
rect 272758 269127 272810 269133
rect 272758 269069 272810 269075
rect 272662 268313 272714 268319
rect 272662 268255 272714 268261
rect 272674 265156 272702 268255
rect 273622 265279 273674 265285
rect 273622 265221 273674 265227
rect 273142 265205 273194 265211
rect 272674 265128 272928 265156
rect 273634 265156 273662 265221
rect 273194 265153 273408 265156
rect 273142 265147 273408 265153
rect 273154 265128 273408 265147
rect 273634 265128 273792 265156
rect 274210 265142 274238 273509
rect 274678 271273 274730 271279
rect 274678 271215 274730 271221
rect 274690 265142 274718 271215
rect 274870 268091 274922 268097
rect 274870 268033 274922 268039
rect 274882 265156 274910 268033
rect 275266 265156 275294 274027
rect 277570 273499 277598 277870
rect 278818 273499 278846 277870
rect 279670 273567 279722 273573
rect 279670 273509 279722 273515
rect 277558 273493 277610 273499
rect 277558 273435 277610 273441
rect 278806 273493 278858 273499
rect 278806 273435 278858 273441
rect 279394 272981 279614 273000
rect 279382 272975 279626 272981
rect 279434 272972 279574 272975
rect 279382 272917 279434 272923
rect 279574 272917 279626 272923
rect 279478 271865 279530 271871
rect 279478 271807 279530 271813
rect 278998 271791 279050 271797
rect 278998 271733 279050 271739
rect 276118 271495 276170 271501
rect 276118 271437 276170 271443
rect 275734 268017 275786 268023
rect 275734 267959 275786 267965
rect 275746 265156 275774 267959
rect 276130 265156 276158 271437
rect 276790 271199 276842 271205
rect 276790 271141 276842 271147
rect 276308 270646 276364 270655
rect 276308 270581 276364 270590
rect 276322 269915 276350 270581
rect 276596 270202 276652 270211
rect 276596 270137 276652 270146
rect 276308 269906 276364 269915
rect 276308 269841 276364 269850
rect 276500 269906 276556 269915
rect 276610 269892 276638 270137
rect 276556 269864 276638 269892
rect 276500 269841 276556 269850
rect 274882 265128 275136 265156
rect 275266 265128 275520 265156
rect 275746 265128 276000 265156
rect 276130 265128 276432 265156
rect 276802 265142 276830 271141
rect 278518 271125 278570 271131
rect 278518 271067 278570 271073
rect 277270 271051 277322 271057
rect 277270 270993 277322 270999
rect 277282 265142 277310 270993
rect 277942 270903 277994 270909
rect 277942 270845 277994 270851
rect 277462 270829 277514 270835
rect 277462 270771 277514 270777
rect 277474 265156 277502 270771
rect 277954 265156 277982 270845
rect 277474 265128 277728 265156
rect 277954 265128 278208 265156
rect 278530 265142 278558 271067
rect 279010 265142 279038 271733
rect 279490 265142 279518 271807
rect 279682 265156 279710 273509
rect 279970 270909 279998 277870
rect 281122 273943 281150 277870
rect 281110 273937 281162 273943
rect 281110 273879 281162 273885
rect 282370 273499 282398 277870
rect 283536 277865 283838 277884
rect 287734 277875 287786 277881
rect 283536 277859 283850 277865
rect 283536 277856 283798 277859
rect 283798 277801 283850 277807
rect 284674 274017 284702 277870
rect 284950 275121 285002 275127
rect 284950 275063 285002 275069
rect 284662 274011 284714 274017
rect 284662 273953 284714 273959
rect 280054 273493 280106 273499
rect 280054 273435 280106 273441
rect 280726 273493 280778 273499
rect 280726 273435 280778 273441
rect 282358 273493 282410 273499
rect 282358 273435 282410 273441
rect 284470 273493 284522 273499
rect 284470 273435 284522 273441
rect 279958 270903 280010 270909
rect 279958 270845 280010 270851
rect 280066 265156 280094 273435
rect 279682 265128 279936 265156
rect 280066 265128 280320 265156
rect 280738 265142 280766 273435
rect 283798 271865 283850 271871
rect 283798 271807 283850 271813
rect 283414 271791 283466 271797
rect 283414 271733 283466 271739
rect 282742 271495 282794 271501
rect 282742 271437 282794 271443
rect 281206 271199 281258 271205
rect 281206 271141 281258 271147
rect 281218 265142 281246 271141
rect 282166 271051 282218 271057
rect 282166 270993 282218 270999
rect 281686 270977 281738 270983
rect 281686 270919 281738 270925
rect 281698 265142 281726 270919
rect 282178 265156 282206 270993
rect 282754 265156 282782 271437
rect 282934 271273 282986 271279
rect 282934 271215 282986 271221
rect 282048 265128 282206 265156
rect 282528 265128 282782 265156
rect 282946 265142 282974 271215
rect 283426 265142 283454 271733
rect 283810 265142 283838 271807
rect 284482 265156 284510 273435
rect 284854 270903 284906 270909
rect 284854 270845 284906 270851
rect 284866 268393 284894 270845
rect 284854 268387 284906 268393
rect 284854 268329 284906 268335
rect 284962 265156 284990 275063
rect 285526 273493 285578 273499
rect 285526 273435 285578 273441
rect 285046 268239 285098 268245
rect 285046 268181 285098 268187
rect 284256 265128 284510 265156
rect 284736 265128 284990 265156
rect 285058 265142 285086 268181
rect 285538 265142 285566 273435
rect 285826 271205 285854 277870
rect 287074 274091 287102 277870
rect 287062 274085 287114 274091
rect 287062 274027 287114 274033
rect 286678 273863 286730 273869
rect 286678 273805 286730 273811
rect 286006 273789 286058 273795
rect 286006 273731 286058 273737
rect 286018 273647 286046 273731
rect 286006 273641 286058 273647
rect 286006 273583 286058 273589
rect 285814 271199 285866 271205
rect 285814 271141 285866 271147
rect 286006 268165 286058 268171
rect 286006 268107 286058 268113
rect 286018 265142 286046 268107
rect 286690 265156 286718 273805
rect 287062 268313 287114 268319
rect 287062 268255 287114 268261
rect 287074 265156 287102 268255
rect 287636 266798 287692 266807
rect 287636 266733 287638 266742
rect 287690 266733 287692 266742
rect 287638 266701 287690 266707
rect 287636 266650 287692 266659
rect 287636 266585 287692 266594
rect 287650 266395 287678 266585
rect 287638 266389 287690 266395
rect 287638 266331 287690 266337
rect 287254 265797 287306 265803
rect 287254 265739 287306 265745
rect 286464 265128 286718 265156
rect 286848 265128 287102 265156
rect 287266 265142 287294 265739
rect 287746 265142 287774 277875
rect 288226 268467 288254 277870
rect 288406 277785 288458 277791
rect 288406 277727 288458 277733
rect 288214 268461 288266 268467
rect 288214 268403 288266 268409
rect 287926 267573 287978 267579
rect 287926 267515 287978 267521
rect 287938 266807 287966 267515
rect 287924 266798 287980 266807
rect 287924 266733 287980 266742
rect 287924 266650 287980 266659
rect 287924 266585 287980 266594
rect 287938 266469 287966 266585
rect 287926 266463 287978 266469
rect 287926 266405 287978 266411
rect 288418 265156 288446 277727
rect 289270 277711 289322 277717
rect 289270 277653 289322 277659
rect 288790 265871 288842 265877
rect 288790 265813 288842 265819
rect 288802 265156 288830 265813
rect 289282 265156 289310 277653
rect 289474 270983 289502 277870
rect 289942 277563 289994 277569
rect 289942 277505 289994 277511
rect 289462 270977 289514 270983
rect 289462 270919 289514 270925
rect 289462 267647 289514 267653
rect 289462 267589 289514 267595
rect 288240 265128 288446 265156
rect 288576 265128 288830 265156
rect 289056 265128 289310 265156
rect 289474 265142 289502 267589
rect 289954 265142 289982 277505
rect 290626 267801 290654 277870
rect 290806 276675 290858 276681
rect 290806 276617 290858 276623
rect 290614 267795 290666 267801
rect 290614 267737 290666 267743
rect 290326 267573 290378 267579
rect 290326 267515 290378 267521
rect 290338 265142 290366 267515
rect 290818 265156 290846 276617
rect 291478 267425 291530 267431
rect 291478 267367 291530 267373
rect 291490 265156 291518 267367
rect 290784 265128 290846 265156
rect 291264 265128 291518 265156
rect 291682 265142 291710 277949
rect 291874 275571 291902 277870
rect 291862 275565 291914 275571
rect 291862 275507 291914 275513
rect 292066 265142 292094 278319
rect 293206 278229 293258 278235
rect 293206 278171 293258 278177
rect 293026 271057 293054 277870
rect 293014 271051 293066 271057
rect 293014 270993 293066 270999
rect 292534 267277 292586 267283
rect 292534 267219 292586 267225
rect 292546 265142 292574 267219
rect 293218 265156 293246 278171
rect 294274 268467 294302 277870
rect 294742 277637 294794 277643
rect 294742 277579 294794 277585
rect 294262 268461 294314 268467
rect 294262 268403 294314 268409
rect 293590 267129 293642 267135
rect 293590 267071 293642 267077
rect 293602 265156 293630 267071
rect 293782 266907 293834 266913
rect 293782 266849 293834 266855
rect 292992 265128 293246 265156
rect 293376 265128 293630 265156
rect 293794 265142 293822 266849
rect 294262 266833 294314 266839
rect 294262 266775 294314 266781
rect 294274 265142 294302 266775
rect 294754 265142 294782 277579
rect 295426 269873 295454 277870
rect 295798 277489 295850 277495
rect 295798 277431 295850 277437
rect 295414 269867 295466 269873
rect 295414 269809 295466 269815
rect 295510 269867 295562 269873
rect 295510 269809 295562 269815
rect 295522 269577 295550 269809
rect 295510 269571 295562 269577
rect 295510 269513 295562 269519
rect 295318 266611 295370 266617
rect 295318 266553 295370 266559
rect 295330 265156 295358 266553
rect 295810 265156 295838 277431
rect 296470 277415 296522 277421
rect 296470 277357 296522 277363
rect 295990 266463 296042 266469
rect 295990 266405 296042 266411
rect 295104 265128 295358 265156
rect 295584 265128 295838 265156
rect 296002 265142 296030 266405
rect 296482 265142 296510 277357
rect 296674 271501 296702 277870
rect 297526 277267 297578 277273
rect 297526 277209 297578 277215
rect 296662 271495 296714 271501
rect 296662 271437 296714 271443
rect 296758 270903 296810 270909
rect 296758 270845 296810 270851
rect 296564 270202 296620 270211
rect 296564 270137 296620 270146
rect 296578 269915 296606 270137
rect 296564 269906 296620 269915
rect 296564 269841 296620 269850
rect 296662 268017 296714 268023
rect 296662 267959 296714 267965
rect 296674 266765 296702 267959
rect 296662 266759 296714 266765
rect 296662 266701 296714 266707
rect 296770 266395 296798 270845
rect 296758 266389 296810 266395
rect 296758 266331 296810 266337
rect 296854 266389 296906 266395
rect 296854 266331 296906 266337
rect 296866 265142 296894 266331
rect 297538 265156 297566 277209
rect 297826 276977 297854 277870
rect 298198 277119 298250 277125
rect 298198 277061 298250 277067
rect 297814 276971 297866 276977
rect 297814 276913 297866 276919
rect 297910 269571 297962 269577
rect 297910 269513 297962 269519
rect 297922 269355 297950 269513
rect 297910 269349 297962 269355
rect 297910 269291 297962 269297
rect 298102 267721 298154 267727
rect 298102 267663 298154 267669
rect 298006 266241 298058 266247
rect 298006 266183 298058 266189
rect 298018 265156 298046 266183
rect 298114 265803 298142 267663
rect 298102 265797 298154 265803
rect 298102 265739 298154 265745
rect 297312 265128 297566 265156
rect 297792 265128 298046 265156
rect 298210 265142 298238 277061
rect 298978 275497 299006 277870
rect 298966 275491 299018 275497
rect 298966 275433 299018 275439
rect 298582 266093 298634 266099
rect 298582 266035 298634 266041
rect 298594 265142 298622 266035
rect 299266 265156 299294 278541
rect 299506 278476 299534 278541
rect 329782 278525 329834 278531
rect 304532 278490 304588 278499
rect 299506 278448 299678 278476
rect 299650 276279 299678 278448
rect 329782 278467 329834 278473
rect 304532 278425 304588 278434
rect 326518 278451 326570 278457
rect 302806 278303 302858 278309
rect 302806 278245 302858 278251
rect 300790 278155 300842 278161
rect 300790 278097 300842 278103
rect 299636 276270 299692 276279
rect 299636 276205 299692 276214
rect 300130 271279 300158 277870
rect 300118 271273 300170 271279
rect 300118 271215 300170 271221
rect 300214 271051 300266 271057
rect 300214 270993 300266 270999
rect 299506 270012 299774 270040
rect 299506 269915 299534 270012
rect 299492 269906 299548 269915
rect 299492 269841 299548 269850
rect 299746 269767 299774 270012
rect 299732 269758 299788 269767
rect 299732 269693 299788 269702
rect 300022 267573 300074 267579
rect 300022 267515 300074 267521
rect 300034 267431 300062 267515
rect 299926 267425 299978 267431
rect 299926 267367 299978 267373
rect 300022 267425 300074 267431
rect 300022 267367 300074 267373
rect 299938 267283 299966 267367
rect 299830 267277 299882 267283
rect 299830 267219 299882 267225
rect 299926 267277 299978 267283
rect 299926 267219 299978 267225
rect 299842 267135 299870 267219
rect 299734 267129 299786 267135
rect 299734 267071 299786 267077
rect 299830 267129 299882 267135
rect 299830 267071 299882 267077
rect 299746 266913 299774 267071
rect 299734 266907 299786 266913
rect 299734 266849 299786 266855
rect 299734 266019 299786 266025
rect 299734 265961 299786 265967
rect 299746 265156 299774 265961
rect 300226 265156 300254 270993
rect 300406 267647 300458 267653
rect 300406 267589 300458 267595
rect 300310 265945 300362 265951
rect 300310 265887 300362 265893
rect 299088 265128 299294 265156
rect 299520 265128 299774 265156
rect 300000 265128 300254 265156
rect 300322 265142 300350 265887
rect 300418 265877 300446 267589
rect 300406 265871 300458 265877
rect 300406 265813 300458 265819
rect 300802 265142 300830 278097
rect 301846 278081 301898 278087
rect 301846 278023 301898 278029
rect 301282 273943 301310 277870
rect 301270 273937 301322 273943
rect 301270 273879 301322 273885
rect 301270 265871 301322 265877
rect 301270 265813 301322 265819
rect 301282 265142 301310 265813
rect 301858 265156 301886 278023
rect 302422 273049 302474 273055
rect 302422 272991 302474 272997
rect 302434 271691 302462 272991
rect 302420 271682 302476 271691
rect 302420 271617 302476 271626
rect 302530 269873 302558 277870
rect 302518 269867 302570 269873
rect 302518 269809 302570 269815
rect 302326 265797 302378 265803
rect 302326 265739 302378 265745
rect 302338 265156 302366 265739
rect 302818 265156 302846 278245
rect 303380 276566 303436 276575
rect 303380 276501 303436 276510
rect 302998 265723 303050 265729
rect 302998 265665 303050 265671
rect 301632 265128 301886 265156
rect 302112 265128 302366 265156
rect 302544 265128 302846 265156
rect 303010 265142 303038 265665
rect 303394 265142 303422 276501
rect 303682 271797 303710 277870
rect 303670 271791 303722 271797
rect 303670 271733 303722 271739
rect 304054 265649 304106 265655
rect 304054 265591 304106 265597
rect 304066 265156 304094 265591
rect 304546 265156 304574 278425
rect 326518 278393 326570 278399
rect 305204 278342 305260 278351
rect 305204 278277 305260 278286
rect 304930 269429 304958 277870
rect 304918 269423 304970 269429
rect 304918 269365 304970 269371
rect 304726 265575 304778 265581
rect 304726 265517 304778 265523
rect 303840 265128 304094 265156
rect 304320 265128 304574 265156
rect 304738 265142 304766 265517
rect 305218 265156 305246 278277
rect 305588 278194 305644 278203
rect 305588 278129 305644 278138
rect 305136 265128 305246 265156
rect 305602 265142 305630 278129
rect 306356 278046 306412 278055
rect 306356 277981 306412 277990
rect 306082 275201 306110 277870
rect 306070 275195 306122 275201
rect 306070 275137 306122 275143
rect 306370 265156 306398 277981
rect 307028 277898 307084 277907
rect 307028 277833 307084 277842
rect 306742 265501 306794 265507
rect 306742 265443 306794 265449
rect 306754 265156 306782 265443
rect 307042 265156 307070 277833
rect 307330 271871 307358 277870
rect 307796 277750 307852 277759
rect 307796 277685 307852 277694
rect 307318 271865 307370 271871
rect 307318 271807 307370 271813
rect 307318 265427 307370 265433
rect 307318 265369 307370 265375
rect 306048 265128 306398 265156
rect 306528 265128 306782 265156
rect 306912 265128 307070 265156
rect 307330 265142 307358 265369
rect 307810 265142 307838 277685
rect 308482 271501 308510 277870
rect 309524 277602 309580 277611
rect 309524 277537 309580 277546
rect 308470 271495 308522 271501
rect 308470 271437 308522 271443
rect 308182 269867 308234 269873
rect 308182 269809 308234 269815
rect 308194 269577 308222 269809
rect 308182 269571 308234 269577
rect 308182 269513 308234 269519
rect 308278 269571 308330 269577
rect 308278 269513 308330 269519
rect 308290 268023 308318 269513
rect 308278 268017 308330 268023
rect 308278 267959 308330 267965
rect 308230 265353 308282 265359
rect 308230 265295 308282 265301
rect 308242 265142 308270 265295
rect 308854 265279 308906 265285
rect 308854 265221 308906 265227
rect 308866 265156 308894 265221
rect 309334 265205 309386 265211
rect 308640 265128 308894 265156
rect 309120 265153 309334 265156
rect 309120 265147 309386 265153
rect 309120 265128 309374 265147
rect 309538 265142 309566 277537
rect 309730 269355 309758 277870
rect 310388 277454 310444 277463
rect 310388 277389 310444 277398
rect 309718 269349 309770 269355
rect 309718 269291 309770 269297
rect 309814 266537 309866 266543
rect 309814 266479 309866 266485
rect 310006 266537 310058 266543
rect 310006 266479 310058 266485
rect 223126 265073 223178 265079
rect 309826 264989 309854 266479
rect 310018 266321 310046 266479
rect 310006 266315 310058 266321
rect 310006 266257 310058 266263
rect 310102 266315 310154 266321
rect 310102 266257 310154 266263
rect 310114 266173 310142 266257
rect 310102 266167 310154 266173
rect 310102 266109 310154 266115
rect 310198 266167 310250 266173
rect 310198 266109 310250 266115
rect 310210 265156 310238 266109
rect 309936 265128 310238 265156
rect 310402 265142 310430 277389
rect 310882 273573 310910 277870
rect 311540 277306 311596 277315
rect 311540 277241 311596 277250
rect 310870 273567 310922 273573
rect 310870 273509 310922 273515
rect 310966 268091 311018 268097
rect 310966 268033 311018 268039
rect 310978 265156 311006 268033
rect 311554 265156 311582 277241
rect 311636 277158 311692 277167
rect 311636 277093 311692 277102
rect 310848 265128 311006 265156
rect 311328 265128 311582 265156
rect 311650 265142 311678 277093
rect 312130 271871 312158 277870
rect 313172 277010 313228 277019
rect 313172 276945 313228 276954
rect 312118 271865 312170 271871
rect 312118 271807 312170 271813
rect 312116 270646 312172 270655
rect 312116 270581 312172 270590
rect 311926 269867 311978 269873
rect 311926 269809 311978 269815
rect 312022 269867 312074 269873
rect 312022 269809 312074 269815
rect 311938 269355 311966 269809
rect 311926 269349 311978 269355
rect 311926 269291 311978 269297
rect 312034 268319 312062 269809
rect 312022 268313 312074 268319
rect 312022 268255 312074 268261
rect 312130 265142 312158 270581
rect 312884 270054 312940 270063
rect 312884 269989 312940 269998
rect 312214 268313 312266 268319
rect 312214 268255 312266 268261
rect 312226 265729 312254 268255
rect 312898 268245 312926 269989
rect 312886 268239 312938 268245
rect 312886 268181 312938 268187
rect 312598 268017 312650 268023
rect 312598 267959 312650 267965
rect 312214 265723 312266 265729
rect 312214 265665 312266 265671
rect 312610 265142 312638 267959
rect 312982 266537 313034 266543
rect 312982 266479 313034 266485
rect 312994 266173 313022 266479
rect 312886 266167 312938 266173
rect 312886 266109 312938 266115
rect 312982 266167 313034 266173
rect 312982 266109 313034 266115
rect 312898 265729 312926 266109
rect 312886 265723 312938 265729
rect 312886 265665 312938 265671
rect 313186 265156 313214 276945
rect 313282 275053 313310 277870
rect 314326 275195 314378 275201
rect 314326 275137 314378 275143
rect 313270 275047 313322 275053
rect 313270 274989 313322 274995
rect 313654 271791 313706 271797
rect 313654 271733 313706 271739
rect 313666 265156 313694 271733
rect 313846 270977 313898 270983
rect 313846 270919 313898 270925
rect 313056 265128 313214 265156
rect 313440 265128 313694 265156
rect 313858 265142 313886 270919
rect 314338 265142 314366 275137
rect 314434 275127 314462 277870
rect 315382 275491 315434 275497
rect 315382 275433 315434 275439
rect 314422 275121 314474 275127
rect 314422 275063 314474 275069
rect 314806 268239 314858 268245
rect 314806 268181 314858 268187
rect 314818 265142 314846 268181
rect 315094 267795 315146 267801
rect 315094 267737 315146 267743
rect 315190 267795 315242 267801
rect 315190 267737 315242 267743
rect 315106 266543 315134 267737
rect 315202 267209 315230 267737
rect 315190 267203 315242 267209
rect 315190 267145 315242 267151
rect 315094 266537 315146 266543
rect 315094 266479 315146 266485
rect 315394 265156 315422 275433
rect 315682 271131 315710 277870
rect 316066 277856 316752 277884
rect 317506 277856 318000 277884
rect 315958 275417 316010 275423
rect 315958 275359 316010 275365
rect 315764 271534 315820 271543
rect 315764 271469 315820 271478
rect 315670 271125 315722 271131
rect 315670 271067 315722 271073
rect 315778 268171 315806 271469
rect 315970 269152 315998 275359
rect 316066 269355 316094 277856
rect 317014 274011 317066 274017
rect 317014 273953 317066 273959
rect 316342 271273 316394 271279
rect 316342 271215 316394 271221
rect 316354 269873 316382 271215
rect 316822 271199 316874 271205
rect 316822 271141 316874 271147
rect 316342 269867 316394 269873
rect 316342 269809 316394 269815
rect 316438 269867 316490 269873
rect 316438 269809 316490 269815
rect 316054 269349 316106 269355
rect 316054 269291 316106 269297
rect 316150 269349 316202 269355
rect 316150 269291 316202 269297
rect 315970 269124 316094 269152
rect 316162 269133 316190 269291
rect 315766 268165 315818 268171
rect 315766 268107 315818 268113
rect 315862 268165 315914 268171
rect 315862 268107 315914 268113
rect 315874 265156 315902 268107
rect 315168 265128 315422 265156
rect 315648 265128 315902 265156
rect 316066 265142 316094 269124
rect 316150 269127 316202 269133
rect 316150 269069 316202 269075
rect 316246 269127 316298 269133
rect 316246 269069 316298 269075
rect 316258 268393 316286 269069
rect 316246 268387 316298 268393
rect 316246 268329 316298 268335
rect 316450 265142 316478 269809
rect 316834 269577 316862 271141
rect 316822 269571 316874 269577
rect 316822 269513 316874 269519
rect 317026 267727 317054 273953
rect 317206 270829 317258 270835
rect 317206 270771 317258 270777
rect 317014 267721 317066 267727
rect 317014 267663 317066 267669
rect 317218 267505 317246 270771
rect 317506 270063 317534 277856
rect 317974 277193 318026 277199
rect 317974 277135 318026 277141
rect 317590 275861 317642 275867
rect 317590 275803 317642 275809
rect 317686 275861 317738 275867
rect 317686 275803 317738 275809
rect 317602 275571 317630 275803
rect 317590 275565 317642 275571
rect 317590 275507 317642 275513
rect 317590 275269 317642 275275
rect 317590 275211 317642 275217
rect 317492 270054 317548 270063
rect 317492 269989 317548 269998
rect 317492 269906 317548 269915
rect 317492 269841 317548 269850
rect 317302 267721 317354 267727
rect 317302 267663 317354 267669
rect 317206 267499 317258 267505
rect 317206 267441 317258 267447
rect 317110 267203 317162 267209
rect 317110 267145 317162 267151
rect 317122 266321 317150 267145
rect 317314 267061 317342 267663
rect 317302 267055 317354 267061
rect 317302 266997 317354 267003
rect 317110 266315 317162 266321
rect 317110 266257 317162 266263
rect 317206 266315 317258 266321
rect 317206 266257 317258 266263
rect 317218 265156 317246 266257
rect 317506 265156 317534 269841
rect 317602 266321 317630 275211
rect 317698 275201 317726 275803
rect 317686 275195 317738 275201
rect 317686 275137 317738 275143
rect 317986 271057 318014 277135
rect 318646 275195 318698 275201
rect 318646 275137 318698 275143
rect 318166 275047 318218 275053
rect 318166 274989 318218 274995
rect 318178 274831 318206 274989
rect 318166 274825 318218 274831
rect 318166 274767 318218 274773
rect 318262 274825 318314 274831
rect 318262 274767 318314 274773
rect 318274 274165 318302 274767
rect 318262 274159 318314 274165
rect 318262 274101 318314 274107
rect 318454 274159 318506 274165
rect 318454 274101 318506 274107
rect 317974 271051 318026 271057
rect 317974 270993 318026 270999
rect 318166 269571 318218 269577
rect 318166 269513 318218 269519
rect 318178 269471 318206 269513
rect 318164 269462 318220 269471
rect 318164 269397 318220 269406
rect 317878 268165 317930 268171
rect 317878 268107 317930 268113
rect 317686 268091 317738 268097
rect 317686 268033 317738 268039
rect 317698 267505 317726 268033
rect 317890 268023 317918 268107
rect 317878 268017 317930 268023
rect 317878 267959 317930 267965
rect 318466 267820 318494 274101
rect 318274 267792 318494 267820
rect 317686 267499 317738 267505
rect 317686 267441 317738 267447
rect 317782 267203 317834 267209
rect 318166 267203 318218 267209
rect 317834 267163 318014 267191
rect 317782 267145 317834 267151
rect 317986 267061 318014 267163
rect 318166 267145 318218 267151
rect 317974 267055 318026 267061
rect 317974 266997 318026 267003
rect 318178 266691 318206 267145
rect 318166 266685 318218 266691
rect 318166 266627 318218 266633
rect 318274 266321 318302 267792
rect 318454 267721 318506 267727
rect 318454 267663 318506 267669
rect 318550 267721 318602 267727
rect 318550 267663 318602 267669
rect 318466 266987 318494 267663
rect 318358 266981 318410 266987
rect 318358 266923 318410 266929
rect 318454 266981 318506 266987
rect 318454 266923 318506 266929
rect 318370 266784 318398 266923
rect 318562 266784 318590 267663
rect 318370 266756 318590 266784
rect 318550 266685 318602 266691
rect 318550 266627 318602 266633
rect 317590 266315 317642 266321
rect 317590 266257 317642 266263
rect 317974 266315 318026 266321
rect 317974 266257 318026 266263
rect 318262 266315 318314 266321
rect 318262 266257 318314 266263
rect 317986 265156 318014 266257
rect 318166 266241 318218 266247
rect 318454 266241 318506 266247
rect 318218 266189 318454 266192
rect 318166 266183 318506 266189
rect 318178 266164 318494 266183
rect 318562 265156 318590 266627
rect 316944 265128 317246 265156
rect 317376 265128 317534 265156
rect 317856 265128 318014 265156
rect 318370 265128 318590 265156
rect 318658 265142 318686 275137
rect 319138 273573 319166 277870
rect 320180 276418 320236 276427
rect 320180 276353 320236 276362
rect 319798 275121 319850 275127
rect 319798 275063 319850 275069
rect 319126 273567 319178 273573
rect 319126 273509 319178 273515
rect 319124 270202 319180 270211
rect 319124 270137 319180 270146
rect 318740 270054 318796 270063
rect 318740 269989 318796 269998
rect 318370 264989 318398 265128
rect 318754 264989 318782 269989
rect 318838 266981 318890 266987
rect 318838 266923 318890 266929
rect 318934 266981 318986 266987
rect 318934 266923 318986 266929
rect 318850 266173 318878 266923
rect 318946 266321 318974 266923
rect 318934 266315 318986 266321
rect 318934 266257 318986 266263
rect 318838 266167 318890 266173
rect 318838 266109 318890 266115
rect 319138 265142 319166 270137
rect 319810 265156 319838 275063
rect 320194 265156 320222 276353
rect 320386 273277 320414 277870
rect 321538 273499 321566 277870
rect 322800 277856 323102 277884
rect 322484 276270 322540 276279
rect 322484 276205 322540 276214
rect 322676 276270 322732 276279
rect 322676 276205 322732 276214
rect 321526 273493 321578 273499
rect 321526 273435 321578 273441
rect 321622 273493 321674 273499
rect 321622 273435 321674 273441
rect 320374 273271 320426 273277
rect 320374 273213 320426 273219
rect 320470 273271 320522 273277
rect 320470 273213 320522 273219
rect 320374 271051 320426 271057
rect 320374 270993 320426 270999
rect 319584 265128 319838 265156
rect 319968 265128 320222 265156
rect 320386 265142 320414 270993
rect 320482 270983 320510 273213
rect 321634 271871 321662 273435
rect 322498 273055 322526 276205
rect 322486 273049 322538 273055
rect 322486 272991 322538 272997
rect 321622 271865 321674 271871
rect 321622 271807 321674 271813
rect 321814 271791 321866 271797
rect 321814 271733 321866 271739
rect 321826 271501 321854 271733
rect 321814 271495 321866 271501
rect 321814 271437 321866 271443
rect 322498 271492 322622 271520
rect 322498 271395 322526 271492
rect 322484 271386 322540 271395
rect 322484 271321 322540 271330
rect 322594 271247 322622 271492
rect 322580 271238 322636 271247
rect 322580 271173 322636 271182
rect 320470 270977 320522 270983
rect 320470 270919 320522 270925
rect 320566 270977 320618 270983
rect 320566 270919 320618 270925
rect 320578 270655 320606 270919
rect 320564 270646 320620 270655
rect 320564 270581 320620 270590
rect 322484 270646 322540 270655
rect 322484 270581 322540 270590
rect 320852 269462 320908 269471
rect 320852 269397 320908 269406
rect 320866 265142 320894 269397
rect 321910 268461 321962 268467
rect 321910 268403 321962 268409
rect 321430 268091 321482 268097
rect 321430 268033 321482 268039
rect 321442 267357 321470 268033
rect 321430 267351 321482 267357
rect 321430 267293 321482 267299
rect 321526 267351 321578 267357
rect 321526 267293 321578 267299
rect 321538 265156 321566 267293
rect 321922 265156 321950 268403
rect 322498 268245 322526 270581
rect 322486 268239 322538 268245
rect 322210 268199 322430 268227
rect 322210 268171 322238 268199
rect 322198 268165 322250 268171
rect 322198 268107 322250 268113
rect 322294 268165 322346 268171
rect 322294 268107 322346 268113
rect 322306 267801 322334 268107
rect 322402 267801 322430 268199
rect 322486 268181 322538 268187
rect 322294 267795 322346 267801
rect 322294 267737 322346 267743
rect 322390 267795 322442 267801
rect 322390 267737 322442 267743
rect 322486 266315 322538 266321
rect 322486 266257 322538 266263
rect 322498 265156 322526 266257
rect 322690 265156 322718 276205
rect 323074 271501 323102 277856
rect 323650 277856 323952 277884
rect 324994 277856 325200 277884
rect 323650 274313 323678 277856
rect 324022 275861 324074 275867
rect 324022 275803 324074 275809
rect 324502 275861 324554 275867
rect 324502 275803 324554 275809
rect 324034 274313 324062 275803
rect 323638 274307 323690 274313
rect 323638 274249 323690 274255
rect 324022 274307 324074 274313
rect 324022 274249 324074 274255
rect 323734 273567 323786 273573
rect 323734 273509 323786 273515
rect 323830 273567 323882 273573
rect 323830 273509 323882 273515
rect 323746 273277 323774 273509
rect 323638 273271 323690 273277
rect 323638 273213 323690 273219
rect 323734 273271 323786 273277
rect 323734 273213 323786 273219
rect 323650 273148 323678 273213
rect 323842 273148 323870 273509
rect 323650 273120 323870 273148
rect 324404 271682 324460 271691
rect 324404 271617 324460 271626
rect 323062 271495 323114 271501
rect 323062 271437 323114 271443
rect 323252 271386 323308 271395
rect 323252 271321 323308 271330
rect 323158 270163 323210 270169
rect 323158 270105 323210 270111
rect 323170 269767 323198 270105
rect 323266 270063 323294 271321
rect 323350 270163 323402 270169
rect 323350 270105 323402 270111
rect 323252 270054 323308 270063
rect 323252 269989 323308 269998
rect 323156 269758 323212 269767
rect 323156 269693 323212 269702
rect 322772 268722 322828 268731
rect 322772 268657 322828 268666
rect 322786 268245 322814 268657
rect 322774 268239 322826 268245
rect 322774 268181 322826 268187
rect 323362 265156 323390 270105
rect 323444 270054 323500 270063
rect 323444 269989 323500 269998
rect 321360 265128 321566 265156
rect 321696 265128 321950 265156
rect 322176 265128 322526 265156
rect 322608 265128 322718 265156
rect 323088 265128 323390 265156
rect 323458 265142 323486 269989
rect 324418 269471 324446 271617
rect 324404 269462 324460 269471
rect 324404 269397 324460 269406
rect 324514 265156 324542 275803
rect 324994 271543 325022 277856
rect 325750 276527 325802 276533
rect 325750 276469 325802 276475
rect 325282 271640 325694 271668
rect 324980 271534 325036 271543
rect 325282 271520 325310 271640
rect 324980 271469 325036 271478
rect 325186 271492 325310 271520
rect 325364 271534 325420 271543
rect 325186 271224 325214 271492
rect 325666 271501 325694 271640
rect 325364 271469 325420 271478
rect 325558 271495 325610 271501
rect 324610 271196 325214 271224
rect 324610 271131 324638 271196
rect 324598 271125 324650 271131
rect 324598 271067 324650 271073
rect 324694 271125 324746 271131
rect 324694 271067 324746 271073
rect 324706 269915 324734 271067
rect 325378 271057 325406 271469
rect 325558 271437 325610 271443
rect 325654 271495 325706 271501
rect 325654 271437 325706 271443
rect 325460 271090 325516 271099
rect 325366 271051 325418 271057
rect 325570 271057 325598 271437
rect 325654 271125 325706 271131
rect 325652 271090 325654 271099
rect 325706 271090 325708 271099
rect 325460 271025 325516 271034
rect 325558 271051 325610 271057
rect 325366 270993 325418 270999
rect 324692 269906 324748 269915
rect 324692 269841 324748 269850
rect 325474 269471 325502 271025
rect 325652 271025 325708 271034
rect 325558 270993 325610 270999
rect 325460 269462 325516 269471
rect 325460 269397 325516 269406
rect 324596 268722 324652 268731
rect 324596 268657 324652 268666
rect 324610 268467 324638 268657
rect 324598 268461 324650 268467
rect 324598 268403 324650 268409
rect 324694 268461 324746 268467
rect 324694 268403 324746 268409
rect 324384 265128 324542 265156
rect 324706 265142 324734 268403
rect 325762 265156 325790 276469
rect 326338 271131 326366 277870
rect 326326 271125 326378 271131
rect 326326 271067 326378 271073
rect 326326 267795 326378 267801
rect 326326 267737 326378 267743
rect 326422 267795 326474 267801
rect 326422 267737 326474 267743
rect 326338 267061 326366 267737
rect 326230 267055 326282 267061
rect 326230 266997 326282 267003
rect 326326 267055 326378 267061
rect 326326 266997 326378 267003
rect 325680 265128 325790 265156
rect 326242 265156 326270 266997
rect 326434 266691 326462 267737
rect 326530 266691 326558 278393
rect 327382 276601 327434 276607
rect 327382 276543 327434 276549
rect 326998 275565 327050 275571
rect 326998 275507 327050 275513
rect 327094 275565 327146 275571
rect 327094 275507 327146 275513
rect 326806 269571 326858 269577
rect 326806 269513 326858 269519
rect 326818 268245 326846 269513
rect 326710 268239 326762 268245
rect 326710 268181 326762 268187
rect 326806 268239 326858 268245
rect 326806 268181 326858 268187
rect 326722 268097 326750 268181
rect 326614 268091 326666 268097
rect 326614 268033 326666 268039
rect 326710 268091 326762 268097
rect 326710 268033 326762 268039
rect 326422 266685 326474 266691
rect 326422 266627 326474 266633
rect 326518 266685 326570 266691
rect 326518 266627 326570 266633
rect 326242 265128 326496 265156
rect 326626 265063 326654 268033
rect 327010 265156 327038 275507
rect 327106 274313 327134 275507
rect 327094 274307 327146 274313
rect 327094 274249 327146 274255
rect 327190 271199 327242 271205
rect 327190 271141 327242 271147
rect 327202 270835 327230 271141
rect 327094 270829 327146 270835
rect 327094 270771 327146 270777
rect 327190 270829 327242 270835
rect 327190 270771 327242 270777
rect 327106 269915 327134 270771
rect 327092 269906 327148 269915
rect 327092 269841 327148 269850
rect 327394 268116 327422 276543
rect 327490 274239 327518 277870
rect 327478 274233 327530 274239
rect 327478 274175 327530 274181
rect 328738 273869 328766 277870
rect 328726 273863 328778 273869
rect 328726 273805 328778 273811
rect 328820 271682 328876 271691
rect 327970 271640 328190 271668
rect 327970 271247 327998 271640
rect 328162 271501 328190 271640
rect 328820 271617 328876 271626
rect 329012 271682 329068 271691
rect 329012 271617 329068 271626
rect 328054 271495 328106 271501
rect 328054 271437 328106 271443
rect 328150 271495 328202 271501
rect 328150 271437 328202 271443
rect 327956 271238 328012 271247
rect 327956 271173 328012 271182
rect 328066 270983 328094 271437
rect 328148 271238 328204 271247
rect 328148 271173 328204 271182
rect 328342 271199 328394 271205
rect 327958 270977 328010 270983
rect 327958 270919 328010 270925
rect 328054 270977 328106 270983
rect 328054 270919 328106 270925
rect 327970 269873 327998 270919
rect 328162 270687 328190 271173
rect 328342 271141 328394 271147
rect 328150 270681 328202 270687
rect 328052 270646 328108 270655
rect 328150 270623 328202 270629
rect 328246 270681 328298 270687
rect 328246 270623 328298 270629
rect 328052 270581 328108 270590
rect 327862 269867 327914 269873
rect 327862 269809 327914 269815
rect 327958 269867 328010 269873
rect 327958 269809 328010 269815
rect 327874 269355 327902 269809
rect 328066 269577 328094 270581
rect 328054 269571 328106 269577
rect 328054 269513 328106 269519
rect 328258 269448 328286 270623
rect 328354 270539 328382 271141
rect 328834 271099 328862 271617
rect 329026 271501 329054 271617
rect 329014 271495 329066 271501
rect 329014 271437 329066 271443
rect 328628 271090 328684 271099
rect 328628 271025 328684 271034
rect 328820 271090 328876 271099
rect 328820 271025 328876 271034
rect 328642 270655 328670 271025
rect 328628 270646 328684 270655
rect 328628 270581 328684 270590
rect 328342 270533 328394 270539
rect 328342 270475 328394 270481
rect 328342 270385 328394 270391
rect 328342 270327 328394 270333
rect 328438 270385 328490 270391
rect 328438 270327 328490 270333
rect 328354 269744 328382 270327
rect 328450 269915 328478 270327
rect 329012 270054 329068 270063
rect 329012 269989 329068 269998
rect 328436 269906 328492 269915
rect 328436 269841 328492 269850
rect 328354 269716 328574 269744
rect 327970 269429 328286 269448
rect 327958 269423 328286 269429
rect 328010 269420 328286 269423
rect 328438 269423 328490 269429
rect 327958 269365 328010 269371
rect 328438 269365 328490 269371
rect 327574 269349 327626 269355
rect 327574 269291 327626 269297
rect 327862 269349 327914 269355
rect 327862 269291 327914 269297
rect 327586 268264 327614 269291
rect 327586 268236 328286 268264
rect 328258 268171 328286 268236
rect 328054 268165 328106 268171
rect 327394 268088 327710 268116
rect 328054 268107 328106 268113
rect 328246 268165 328298 268171
rect 328246 268107 328298 268113
rect 327574 267795 327626 267801
rect 327574 267737 327626 267743
rect 327586 267061 327614 267737
rect 327574 267055 327626 267061
rect 327574 266997 327626 267003
rect 327382 266981 327434 266987
rect 327382 266923 327434 266929
rect 326928 265128 327038 265156
rect 327394 265142 327422 266923
rect 327682 265156 327710 268088
rect 328066 267801 328094 268107
rect 328450 268023 328478 269365
rect 328546 268023 328574 269716
rect 329026 269471 329054 269989
rect 328820 269462 328876 269471
rect 328820 269397 328876 269406
rect 329012 269462 329068 269471
rect 329012 269397 329068 269406
rect 328834 268731 328862 269397
rect 328628 268722 328684 268731
rect 328628 268657 328684 268666
rect 328820 268722 328876 268731
rect 328820 268657 328876 268666
rect 328642 268560 328670 268657
rect 328642 268532 329150 268560
rect 328438 268017 328490 268023
rect 328438 267959 328490 267965
rect 328534 268017 328586 268023
rect 328534 267959 328586 267965
rect 328436 267834 328492 267843
rect 328054 267795 328106 267801
rect 328492 267792 329054 267820
rect 328436 267769 328492 267778
rect 328054 267737 328106 267743
rect 328918 267721 328970 267727
rect 328642 267681 328918 267709
rect 327766 267499 327818 267505
rect 328642 267487 328670 267681
rect 328918 267663 328970 267669
rect 328726 267647 328778 267653
rect 328778 267607 328862 267635
rect 328726 267589 328778 267595
rect 327818 267459 328670 267487
rect 327766 267441 327818 267447
rect 327958 267425 328010 267431
rect 328342 267425 328394 267431
rect 328010 267385 328342 267413
rect 327958 267367 328010 267373
rect 328342 267367 328394 267373
rect 328246 267351 328298 267357
rect 328066 267311 328246 267339
rect 328066 267103 328094 267311
rect 328246 267293 328298 267299
rect 328246 267203 328298 267209
rect 328246 267145 328298 267151
rect 328438 267203 328490 267209
rect 328438 267145 328490 267151
rect 328052 267094 328108 267103
rect 327958 267055 328010 267061
rect 328258 267061 328286 267145
rect 328340 267094 328396 267103
rect 328052 267029 328108 267038
rect 328246 267055 328298 267061
rect 327958 266997 328010 267003
rect 328340 267029 328396 267038
rect 328246 266997 328298 267003
rect 327970 265156 327998 266997
rect 328354 266987 328382 267029
rect 328342 266981 328394 266987
rect 328450 266955 328478 267145
rect 328342 266923 328394 266929
rect 328436 266946 328492 266955
rect 328436 266881 328492 266890
rect 328628 266946 328684 266955
rect 328628 266881 328684 266890
rect 328054 266685 328106 266691
rect 328054 266627 328106 266633
rect 328532 266650 328588 266659
rect 328066 265304 328094 266627
rect 328246 266611 328298 266617
rect 328532 266585 328588 266594
rect 328246 266553 328298 266559
rect 328258 266192 328286 266553
rect 328546 266543 328574 266585
rect 328534 266537 328586 266543
rect 328534 266479 328586 266485
rect 328642 266321 328670 266881
rect 328834 266321 328862 267607
rect 329026 267135 329054 267792
rect 329122 267709 329150 268532
rect 329314 267940 329726 267968
rect 329314 267801 329342 267940
rect 329302 267795 329354 267801
rect 329302 267737 329354 267743
rect 329398 267795 329450 267801
rect 329398 267737 329450 267743
rect 329410 267709 329438 267737
rect 329122 267681 329438 267709
rect 329014 267129 329066 267135
rect 329014 267071 329066 267077
rect 329300 266650 329356 266659
rect 328918 266611 328970 266617
rect 329300 266585 329356 266594
rect 328918 266553 328970 266559
rect 328630 266315 328682 266321
rect 328630 266257 328682 266263
rect 328822 266315 328874 266321
rect 328822 266257 328874 266263
rect 328930 266192 328958 266553
rect 328258 266164 328958 266192
rect 328066 265276 328382 265304
rect 327682 265128 327888 265156
rect 327970 265128 328224 265156
rect 325846 265057 325898 265063
rect 323904 264989 324158 265008
rect 325200 264994 325502 265008
rect 326614 265057 326666 265063
rect 325898 265005 326112 265008
rect 325846 264999 326112 265005
rect 326614 264999 326666 265005
rect 309814 264983 309866 264989
rect 309814 264925 309866 264931
rect 318358 264983 318410 264989
rect 318358 264925 318410 264931
rect 318454 264983 318506 264989
rect 318454 264925 318506 264931
rect 318742 264983 318794 264989
rect 323904 264983 324170 264989
rect 323904 264980 324118 264983
rect 318742 264925 318794 264931
rect 325200 264985 325516 264994
rect 325200 264980 325460 264985
rect 324118 264925 324170 264931
rect 325858 264980 326112 264999
rect 318466 264860 318494 264925
rect 325460 264920 325516 264929
rect 318192 264832 318494 264860
rect 328354 264860 328382 265276
rect 329026 265137 329136 265156
rect 329014 265131 329136 265137
rect 329066 265128 329136 265131
rect 329014 265073 329066 265079
rect 329314 264989 329342 266585
rect 329698 265137 329726 267940
rect 329686 265131 329738 265137
rect 329686 265073 329738 265079
rect 329794 265008 329822 278467
rect 339094 277933 339146 277939
rect 329986 271797 330014 277870
rect 330850 277856 331152 277884
rect 330166 275047 330218 275053
rect 330166 274989 330218 274995
rect 329878 271791 329930 271797
rect 329878 271733 329930 271739
rect 329974 271791 330026 271797
rect 329974 271733 330026 271739
rect 329890 271501 329918 271733
rect 329878 271495 329930 271501
rect 329878 271437 329930 271443
rect 330070 268313 330122 268319
rect 330070 268255 330122 268261
rect 330082 266987 330110 268255
rect 329974 266981 330026 266987
rect 329974 266923 330026 266929
rect 330070 266981 330122 266987
rect 330070 266923 330122 266929
rect 329986 265142 330014 266923
rect 330178 265156 330206 274989
rect 330850 271247 330878 277856
rect 331318 277341 331370 277347
rect 331318 277283 331370 277289
rect 330836 271238 330892 271247
rect 330836 271173 330892 271182
rect 331222 271199 331274 271205
rect 331222 271141 331274 271147
rect 331234 270539 331262 271141
rect 331222 270533 331274 270539
rect 331222 270475 331274 270481
rect 330646 267647 330698 267653
rect 330646 267589 330698 267595
rect 330658 265156 330686 267589
rect 330178 265128 330432 265156
rect 330658 265128 330912 265156
rect 331330 265142 331358 277283
rect 332182 276749 332234 276755
rect 332182 276691 332234 276697
rect 331894 267129 331946 267135
rect 331894 267071 331946 267077
rect 331906 266173 331934 267071
rect 331702 266167 331754 266173
rect 331702 266109 331754 266115
rect 331894 266167 331946 266173
rect 331894 266109 331946 266115
rect 331714 265142 331742 266109
rect 332194 265142 332222 276691
rect 332290 271279 332318 277870
rect 332758 277045 332810 277051
rect 332758 276987 332810 276993
rect 332278 271273 332330 271279
rect 332278 271215 332330 271221
rect 332566 267795 332618 267801
rect 332566 267737 332618 267743
rect 332578 267653 332606 267737
rect 332566 267647 332618 267653
rect 332566 267589 332618 267595
rect 332770 265156 332798 276987
rect 333442 268319 333470 277870
rect 334486 276897 334538 276903
rect 334486 276839 334538 276845
rect 333910 276823 333962 276829
rect 333910 276765 333962 276771
rect 333430 268313 333482 268319
rect 333430 268255 333482 268261
rect 332386 265137 332640 265156
rect 332374 265131 332640 265137
rect 332426 265128 332640 265131
rect 332770 265128 333024 265156
rect 333922 265142 333950 276765
rect 334102 273493 334154 273499
rect 334102 273435 334154 273441
rect 334114 271279 334142 273435
rect 334102 271273 334154 271279
rect 334102 271215 334154 271221
rect 334102 270385 334154 270391
rect 334102 270327 334154 270333
rect 334114 265156 334142 270327
rect 334498 265156 334526 276839
rect 334594 276459 334622 277870
rect 335458 277856 335856 277884
rect 339146 277881 339408 277884
rect 339094 277875 339408 277881
rect 336310 277859 336362 277865
rect 334582 276453 334634 276459
rect 334582 276395 334634 276401
rect 335458 274017 335486 277856
rect 336310 277801 336362 277807
rect 335638 274825 335690 274831
rect 335638 274767 335690 274773
rect 335446 274011 335498 274017
rect 335446 273953 335498 273959
rect 334966 268165 335018 268171
rect 334966 268107 335018 268113
rect 334978 265156 335006 268107
rect 334114 265128 334416 265156
rect 334498 265128 334752 265156
rect 334978 265128 335232 265156
rect 335650 265142 335678 274767
rect 336214 269645 336266 269651
rect 336214 269587 336266 269593
rect 336226 269133 336254 269587
rect 336118 269127 336170 269133
rect 336118 269069 336170 269075
rect 336214 269127 336266 269133
rect 336214 269069 336266 269075
rect 336130 265142 336158 269069
rect 336322 265156 336350 277801
rect 336694 274085 336746 274091
rect 336694 274027 336746 274033
rect 336598 270311 336650 270317
rect 336598 270253 336650 270259
rect 336610 269767 336638 270253
rect 336596 269758 336652 269767
rect 336596 269693 336652 269702
rect 336706 265156 336734 274027
rect 336994 273499 337022 277870
rect 338134 276971 338186 276977
rect 338134 276913 338186 276919
rect 336982 273493 337034 273499
rect 336982 273435 337034 273441
rect 336980 271386 337036 271395
rect 336980 271321 337036 271330
rect 336994 270211 337022 271321
rect 336980 270202 337036 270211
rect 336886 270163 336938 270169
rect 336980 270137 337036 270146
rect 336886 270105 336938 270111
rect 336898 267801 336926 270105
rect 338038 268461 338090 268467
rect 338038 268403 338090 268409
rect 337846 268387 337898 268393
rect 337846 268329 337898 268335
rect 336886 267795 336938 267801
rect 336886 267737 336938 267743
rect 337654 267647 337706 267653
rect 337654 267589 337706 267595
rect 337462 267499 337514 267505
rect 337462 267441 337514 267447
rect 337174 267055 337226 267061
rect 337174 266997 337226 267003
rect 337186 265729 337214 266997
rect 337474 266987 337502 267441
rect 337366 266981 337418 266987
rect 337366 266923 337418 266929
rect 337462 266981 337514 266987
rect 337462 266923 337514 266929
rect 337378 266784 337406 266923
rect 337378 266756 337598 266784
rect 337270 266685 337322 266691
rect 337270 266627 337322 266633
rect 337174 265723 337226 265729
rect 337174 265665 337226 265671
rect 337282 265156 337310 266627
rect 337570 265729 337598 266756
rect 337666 266691 337694 267589
rect 337654 266685 337706 266691
rect 337654 266627 337706 266633
rect 337558 265723 337610 265729
rect 337558 265665 337610 265671
rect 336322 265128 336528 265156
rect 336706 265128 336960 265156
rect 337282 265128 337440 265156
rect 337858 265142 337886 268329
rect 337942 267425 337994 267431
rect 337942 267367 337994 267373
rect 337954 267209 337982 267367
rect 338050 267209 338078 268403
rect 337942 267203 337994 267209
rect 337942 267145 337994 267151
rect 338038 267203 338090 267209
rect 338038 267145 338090 267151
rect 338146 265156 338174 276913
rect 338242 270539 338270 277870
rect 339106 277856 339408 277875
rect 338422 275195 338474 275201
rect 338422 275137 338474 275143
rect 338434 274313 338462 275137
rect 338422 274307 338474 274313
rect 338422 274249 338474 274255
rect 338710 273937 338762 273943
rect 338710 273879 338762 273885
rect 338230 270533 338282 270539
rect 338230 270475 338282 270481
rect 338326 270533 338378 270539
rect 338326 270475 338378 270481
rect 338338 269873 338366 270475
rect 338326 269867 338378 269873
rect 338326 269809 338378 269815
rect 338146 265128 338256 265156
rect 338722 265142 338750 273879
rect 339586 273055 339614 278596
rect 339874 278457 339902 278596
rect 374324 278638 374380 278647
rect 372884 278573 372940 278582
rect 374146 278596 374324 278624
rect 372898 278531 372926 278573
rect 350326 278525 350378 278531
rect 350326 278467 350378 278473
rect 351766 278525 351818 278531
rect 351766 278467 351818 278473
rect 372502 278525 372554 278531
rect 372502 278467 372554 278473
rect 372886 278525 372938 278531
rect 372886 278467 372938 278473
rect 339862 278451 339914 278457
rect 339862 278393 339914 278399
rect 340642 273277 340670 277870
rect 341794 276385 341822 277870
rect 342754 277856 342960 277884
rect 342754 277791 342782 277856
rect 342742 277785 342794 277791
rect 342742 277727 342794 277733
rect 341782 276379 341834 276385
rect 341782 276321 341834 276327
rect 343126 273863 343178 273869
rect 343126 273805 343178 273811
rect 343030 273493 343082 273499
rect 343030 273435 343082 273441
rect 340534 273271 340586 273277
rect 340534 273213 340586 273219
rect 340630 273271 340682 273277
rect 340630 273213 340682 273219
rect 339574 273049 339626 273055
rect 339574 272991 339626 272997
rect 339766 273049 339818 273055
rect 339766 272991 339818 272997
rect 339382 271495 339434 271501
rect 339382 271437 339434 271443
rect 338902 270681 338954 270687
rect 338902 270623 338954 270629
rect 338806 267499 338858 267505
rect 338806 267441 338858 267447
rect 338818 266543 338846 267441
rect 338806 266537 338858 266543
rect 338806 266479 338858 266485
rect 338914 265156 338942 270623
rect 339394 265156 339422 271437
rect 339778 271247 339806 272991
rect 339862 271273 339914 271279
rect 339764 271238 339820 271247
rect 339862 271215 339914 271221
rect 339764 271173 339820 271182
rect 339874 265156 339902 271215
rect 340438 270977 340490 270983
rect 340438 270919 340490 270925
rect 338914 265128 339168 265156
rect 339394 265128 339648 265156
rect 339874 265128 340032 265156
rect 340450 265142 340478 270919
rect 340546 265156 340574 273213
rect 341782 271791 341834 271797
rect 341782 271733 341834 271739
rect 341494 271125 341546 271131
rect 341494 271067 341546 271073
rect 341302 271051 341354 271057
rect 341302 270993 341354 270999
rect 340546 265128 340944 265156
rect 341314 265142 341342 270993
rect 341506 265156 341534 271067
rect 341794 265304 341822 271733
rect 342452 271090 342508 271099
rect 342452 271025 342508 271034
rect 341974 270681 342026 270687
rect 341974 270623 342026 270629
rect 341878 270089 341930 270095
rect 341878 270031 341930 270037
rect 341890 269725 341918 270031
rect 341878 269719 341930 269725
rect 341878 269661 341930 269667
rect 341986 269503 342014 270623
rect 342166 270163 342218 270169
rect 342166 270105 342218 270111
rect 342178 269873 342206 270105
rect 342466 269892 342494 271025
rect 342548 269906 342604 269915
rect 342166 269867 342218 269873
rect 342466 269864 342548 269892
rect 342548 269841 342604 269850
rect 342166 269809 342218 269815
rect 342550 269793 342602 269799
rect 342602 269753 342782 269781
rect 342550 269735 342602 269741
rect 341974 269497 342026 269503
rect 341974 269439 342026 269445
rect 342082 269281 342494 269300
rect 342070 269275 342506 269281
rect 342122 269272 342454 269275
rect 342070 269217 342122 269223
rect 342454 269217 342506 269223
rect 341974 269201 342026 269207
rect 342550 269201 342602 269207
rect 342026 269149 342550 269152
rect 341974 269143 342602 269149
rect 341986 269124 342590 269143
rect 342754 269133 342782 269753
rect 342838 269645 342890 269651
rect 342838 269587 342890 269593
rect 342646 269127 342698 269133
rect 342646 269069 342698 269075
rect 342742 269127 342794 269133
rect 342742 269069 342794 269075
rect 342658 269004 342686 269069
rect 342850 269004 342878 269587
rect 342658 268976 342878 269004
rect 342646 268313 342698 268319
rect 342646 268255 342698 268261
rect 341794 265276 341918 265304
rect 341890 265156 341918 265276
rect 341506 265128 341760 265156
rect 341890 265128 342240 265156
rect 342658 265142 342686 268255
rect 343042 265142 343070 273435
rect 343138 270317 343166 273805
rect 343510 273271 343562 273277
rect 343510 273213 343562 273219
rect 343126 270311 343178 270317
rect 343126 270253 343178 270259
rect 343522 265142 343550 273213
rect 343702 267425 343754 267431
rect 343702 267367 343754 267373
rect 332374 265073 332426 265079
rect 329302 264983 329354 264989
rect 329616 264980 329822 265008
rect 333142 265057 333194 265063
rect 333194 265005 333456 265008
rect 333142 264999 333456 265005
rect 333154 264980 333456 264999
rect 329302 264925 329354 264931
rect 343714 264915 343742 267367
rect 344194 265156 344222 277870
rect 344662 273271 344714 273277
rect 344662 273213 344714 273219
rect 344674 265156 344702 273213
rect 345238 271125 345290 271131
rect 345238 271067 345290 271073
rect 344758 271051 344810 271057
rect 344758 270993 344810 270999
rect 343968 265128 344222 265156
rect 344448 265128 344702 265156
rect 344770 265142 344798 270993
rect 345250 265142 345278 271067
rect 345346 268023 345374 277870
rect 345718 271199 345770 271205
rect 345718 271141 345770 271147
rect 345334 268017 345386 268023
rect 345334 267959 345386 267965
rect 345730 265142 345758 271141
rect 346390 270977 346442 270983
rect 346390 270919 346442 270925
rect 346402 265156 346430 270919
rect 346594 266321 346622 277870
rect 347446 273493 347498 273499
rect 347446 273435 347498 273441
rect 347254 271791 347306 271797
rect 347254 271733 347306 271739
rect 346774 271495 346826 271501
rect 346774 271437 346826 271443
rect 346582 266315 346634 266321
rect 346582 266257 346634 266263
rect 346786 265156 346814 271437
rect 347158 268091 347210 268097
rect 347158 268033 347210 268039
rect 347170 267579 347198 268033
rect 347158 267573 347210 267579
rect 347158 267515 347210 267521
rect 347266 265156 347294 271733
rect 346176 265128 346430 265156
rect 346560 265128 346814 265156
rect 346992 265128 347294 265156
rect 347458 265142 347486 273435
rect 347746 273277 347774 277870
rect 348994 276163 349022 277870
rect 350050 277717 350078 277870
rect 350038 277711 350090 277717
rect 350038 277653 350090 277659
rect 349174 276749 349226 276755
rect 349174 276691 349226 276697
rect 348982 276157 349034 276163
rect 348982 276099 349034 276105
rect 347734 273271 347786 273277
rect 347734 273213 347786 273219
rect 347926 273271 347978 273277
rect 347926 273213 347978 273219
rect 347830 267573 347882 267579
rect 347830 267515 347882 267521
rect 347842 267357 347870 267515
rect 347830 267351 347882 267357
rect 347830 267293 347882 267299
rect 347828 266946 347884 266955
rect 347828 266881 347884 266890
rect 347732 266650 347788 266659
rect 347732 266585 347788 266594
rect 347746 264989 347774 266585
rect 347842 266543 347870 266881
rect 347830 266537 347882 266543
rect 347830 266479 347882 266485
rect 347938 265142 347966 273213
rect 348214 270533 348266 270539
rect 348214 270475 348266 270481
rect 348406 270533 348458 270539
rect 348406 270475 348458 270481
rect 348118 270089 348170 270095
rect 348118 270031 348170 270037
rect 348130 269725 348158 270031
rect 348226 269873 348254 270475
rect 348310 270237 348362 270243
rect 348310 270179 348362 270185
rect 348322 270095 348350 270179
rect 348310 270089 348362 270095
rect 348310 270031 348362 270037
rect 348214 269867 348266 269873
rect 348214 269809 348266 269815
rect 348118 269719 348170 269725
rect 348118 269661 348170 269667
rect 348214 267425 348266 267431
rect 348214 267367 348266 267373
rect 348226 267209 348254 267367
rect 348214 267203 348266 267209
rect 348214 267145 348266 267151
rect 348022 266981 348074 266987
rect 348022 266923 348074 266929
rect 348034 266321 348062 266923
rect 348022 266315 348074 266321
rect 348022 266257 348074 266263
rect 348418 265156 348446 270475
rect 348788 267834 348844 267843
rect 348788 267769 348844 267778
rect 348980 267834 349036 267843
rect 348980 267769 349036 267778
rect 348502 267499 348554 267505
rect 348502 267441 348554 267447
rect 348514 267357 348542 267441
rect 348694 267425 348746 267431
rect 348694 267367 348746 267373
rect 348502 267351 348554 267357
rect 348502 267293 348554 267299
rect 348706 267283 348734 267367
rect 348694 267277 348746 267283
rect 348694 267219 348746 267225
rect 348598 267203 348650 267209
rect 348598 267145 348650 267151
rect 348500 266946 348556 266955
rect 348610 266932 348638 267145
rect 348802 266955 348830 267769
rect 348994 267579 349022 267769
rect 348982 267573 349034 267579
rect 348982 267515 349034 267521
rect 348982 267203 349034 267209
rect 348982 267145 349034 267151
rect 348556 266904 348638 266932
rect 348788 266946 348844 266955
rect 348500 266881 348556 266890
rect 348788 266881 348844 266890
rect 348692 266798 348748 266807
rect 348610 266756 348692 266784
rect 348610 266543 348638 266756
rect 348692 266733 348748 266742
rect 348598 266537 348650 266543
rect 348598 266479 348650 266485
rect 348994 265156 349022 267145
rect 349076 266650 349132 266659
rect 349076 266585 349132 266594
rect 349090 266543 349118 266585
rect 349078 266537 349130 266543
rect 349078 266479 349130 266485
rect 348288 265128 348446 265156
rect 348768 265128 349022 265156
rect 349186 265142 349214 276691
rect 349846 273493 349898 273499
rect 349846 273435 349898 273441
rect 349858 273277 349886 273435
rect 349750 273271 349802 273277
rect 349750 273213 349802 273219
rect 349846 273271 349898 273277
rect 349846 273213 349898 273219
rect 349762 271501 349790 273213
rect 349654 271495 349706 271501
rect 349654 271437 349706 271443
rect 349750 271495 349802 271501
rect 349750 271437 349802 271443
rect 349558 271273 349610 271279
rect 349558 271215 349610 271221
rect 349570 270983 349598 271215
rect 349666 270983 349694 271437
rect 349558 270977 349610 270983
rect 349558 270919 349610 270925
rect 349654 270977 349706 270983
rect 349654 270919 349706 270925
rect 349846 268017 349898 268023
rect 349846 267959 349898 267965
rect 349858 267727 349886 267959
rect 349846 267721 349898 267727
rect 349846 267663 349898 267669
rect 349846 267499 349898 267505
rect 349846 267441 349898 267447
rect 349364 267094 349420 267103
rect 349858 267061 349886 267441
rect 349364 267029 349420 267038
rect 349846 267055 349898 267061
rect 349378 266987 349406 267029
rect 349846 266997 349898 267003
rect 349366 266981 349418 266987
rect 349366 266923 349418 266929
rect 349844 266650 349900 266659
rect 349844 266585 349900 266594
rect 349858 266321 349886 266585
rect 349846 266315 349898 266321
rect 349846 266257 349898 266263
rect 349942 266315 349994 266321
rect 349942 266257 349994 266263
rect 349954 266173 349982 266257
rect 349942 266167 349994 266173
rect 349942 266109 349994 266115
rect 350338 265156 350366 278467
rect 351010 277856 351312 277884
rect 351010 271057 351038 277856
rect 351094 277341 351146 277347
rect 351094 277283 351146 277289
rect 350998 271051 351050 271057
rect 350998 270993 351050 270999
rect 350710 267499 350762 267505
rect 350710 267441 350762 267447
rect 350722 265156 350750 267441
rect 351106 265156 351134 277283
rect 351190 273493 351242 273499
rect 351190 273435 351242 273441
rect 351202 271279 351230 273435
rect 351190 271273 351242 271279
rect 351190 271215 351242 271221
rect 351286 271273 351338 271279
rect 351286 271215 351338 271221
rect 351298 270951 351326 271215
rect 351284 270942 351340 270951
rect 351284 270877 351340 270886
rect 351286 266167 351338 266173
rect 351286 266109 351338 266115
rect 349584 265137 349886 265156
rect 349584 265131 349898 265137
rect 349584 265128 349846 265131
rect 350064 265128 350366 265156
rect 350496 265128 350750 265156
rect 350976 265128 351134 265156
rect 351298 265142 351326 266109
rect 351778 265142 351806 278467
rect 366358 278451 366410 278457
rect 366358 278393 366410 278399
rect 352918 277933 352970 277939
rect 352918 277875 352970 277881
rect 352450 270391 352478 277870
rect 352438 270385 352490 270391
rect 352438 270327 352490 270333
rect 352246 267721 352298 267727
rect 352246 267663 352298 267669
rect 352258 265142 352286 267663
rect 352930 265156 352958 277875
rect 353494 274085 353546 274091
rect 353494 274027 353546 274033
rect 353302 270385 353354 270391
rect 353302 270327 353354 270333
rect 353314 265156 353342 270327
rect 352704 265128 352958 265156
rect 353088 265128 353342 265156
rect 353506 265142 353534 274027
rect 353698 267653 353726 277870
rect 354454 277859 354506 277865
rect 354454 277801 354506 277807
rect 353686 267647 353738 267653
rect 353686 267589 353738 267595
rect 354262 267647 354314 267653
rect 354262 267589 354314 267595
rect 354274 267209 354302 267589
rect 354262 267203 354314 267209
rect 354262 267145 354314 267151
rect 353974 266981 354026 266987
rect 353974 266923 354026 266929
rect 353986 265142 354014 266923
rect 354466 265142 354494 277801
rect 354850 271131 354878 277870
rect 355798 277785 355850 277791
rect 355798 277727 355850 277733
rect 355702 274159 355754 274165
rect 355702 274101 355754 274107
rect 355222 271199 355274 271205
rect 355222 271141 355274 271147
rect 354838 271125 354890 271131
rect 354838 271067 354890 271073
rect 355234 270803 355262 271141
rect 355220 270794 355276 270803
rect 355220 270729 355276 270738
rect 355414 270163 355466 270169
rect 355414 270105 355466 270111
rect 355426 268911 355454 270105
rect 355606 270089 355658 270095
rect 355606 270031 355658 270037
rect 355414 268905 355466 268911
rect 355414 268847 355466 268853
rect 355510 268905 355562 268911
rect 355510 268847 355562 268853
rect 355414 268313 355466 268319
rect 355414 268255 355466 268261
rect 355426 267949 355454 268255
rect 355414 267943 355466 267949
rect 355414 267885 355466 267891
rect 355030 267203 355082 267209
rect 355030 267145 355082 267151
rect 355042 265156 355070 267145
rect 355522 265156 355550 268847
rect 355618 268245 355646 270031
rect 355606 268239 355658 268245
rect 355606 268181 355658 268187
rect 354816 265128 355070 265156
rect 355296 265128 355550 265156
rect 355714 265142 355742 274101
rect 355810 265156 355838 277727
rect 356098 276015 356126 277870
rect 357250 277569 357278 277870
rect 357238 277563 357290 277569
rect 357238 277505 357290 277511
rect 357718 276897 357770 276903
rect 357718 276839 357770 276845
rect 356086 276009 356138 276015
rect 356086 275951 356138 275957
rect 356948 270942 357004 270951
rect 356948 270877 357004 270886
rect 355894 268239 355946 268245
rect 355894 268181 355946 268187
rect 355906 268097 355934 268181
rect 356962 268139 356990 270877
rect 357046 268461 357098 268467
rect 357046 268403 357098 268409
rect 356948 268130 357004 268139
rect 355894 268091 355946 268097
rect 356948 268065 357004 268074
rect 355894 268033 355946 268039
rect 356854 267721 356906 267727
rect 356854 267663 356906 267669
rect 356950 267721 357002 267727
rect 356950 267663 357002 267669
rect 356866 267505 356894 267663
rect 356962 267579 356990 267663
rect 356950 267573 357002 267579
rect 356950 267515 357002 267521
rect 356854 267499 356906 267505
rect 356854 267441 356906 267447
rect 357058 265156 357086 268403
rect 357622 268387 357674 268393
rect 357622 268329 357674 268335
rect 357430 268165 357482 268171
rect 357430 268107 357482 268113
rect 357334 267869 357386 267875
rect 357442 267857 357470 268107
rect 357386 267829 357470 267857
rect 357334 267811 357386 267817
rect 357634 266784 357662 268329
rect 357538 266756 357662 266784
rect 357538 266543 357566 266756
rect 357526 266537 357578 266543
rect 357526 266479 357578 266485
rect 357730 265156 357758 276839
rect 358102 274011 358154 274017
rect 358102 273953 358154 273959
rect 357812 267834 357868 267843
rect 357812 267769 357868 267778
rect 357826 266321 357854 267769
rect 357814 266315 357866 266321
rect 357814 266257 357866 266263
rect 358114 265156 358142 273953
rect 358402 271131 358430 277870
rect 358774 277711 358826 277717
rect 358774 277653 358826 277659
rect 358486 271791 358538 271797
rect 358486 271733 358538 271739
rect 358582 271791 358634 271797
rect 358582 271733 358634 271739
rect 358498 271131 358526 271733
rect 358594 271501 358622 271733
rect 358582 271495 358634 271501
rect 358582 271437 358634 271443
rect 358390 271125 358442 271131
rect 358390 271067 358442 271073
rect 358486 271125 358538 271131
rect 358486 271067 358538 271073
rect 358486 270977 358538 270983
rect 358486 270919 358538 270925
rect 358498 270761 358526 270919
rect 358486 270755 358538 270761
rect 358486 270697 358538 270703
rect 358678 268017 358730 268023
rect 358678 267959 358730 267965
rect 358690 267357 358718 267959
rect 358678 267351 358730 267357
rect 358678 267293 358730 267299
rect 358294 266537 358346 266543
rect 358294 266479 358346 266485
rect 355810 265128 356208 265156
rect 357024 265128 357086 265156
rect 357504 265128 357758 265156
rect 357840 265128 358142 265156
rect 358306 265142 358334 266479
rect 358786 265142 358814 277653
rect 359650 273869 359678 277870
rect 360226 277856 360816 277884
rect 359734 274233 359786 274239
rect 359734 274175 359786 274181
rect 359638 273863 359690 273869
rect 359638 273805 359690 273811
rect 359446 270311 359498 270317
rect 359446 270253 359498 270259
rect 359062 267869 359114 267875
rect 359062 267811 359114 267817
rect 359074 267283 359102 267811
rect 359062 267277 359114 267283
rect 359062 267219 359114 267225
rect 359158 267277 359210 267283
rect 359158 267219 359210 267225
rect 359170 266173 359198 267219
rect 359158 266167 359210 266173
rect 359158 266109 359210 266115
rect 359458 265156 359486 270253
rect 359746 265156 359774 274175
rect 360118 268313 360170 268319
rect 360118 268255 360170 268261
rect 360130 268153 360158 268255
rect 360226 268245 360254 277856
rect 360502 277045 360554 277051
rect 360502 276987 360554 276993
rect 360406 268313 360458 268319
rect 360322 268273 360406 268301
rect 360214 268239 360266 268245
rect 360214 268181 360266 268187
rect 360322 268153 360350 268273
rect 360406 268255 360458 268261
rect 360130 268125 360350 268153
rect 360022 266167 360074 266173
rect 360022 266109 360074 266115
rect 359232 265128 359486 265156
rect 359616 265128 359774 265156
rect 360034 265142 360062 266109
rect 360514 265142 360542 276987
rect 361942 273863 361994 273869
rect 361942 273805 361994 273811
rect 360982 269497 361034 269503
rect 360982 269439 361034 269445
rect 360886 268905 360938 268911
rect 360886 268847 360938 268853
rect 360898 268393 360926 268847
rect 360886 268387 360938 268393
rect 360886 268329 360938 268335
rect 360994 265142 361022 269439
rect 361558 267573 361610 267579
rect 361558 267515 361610 267521
rect 361570 265156 361598 267515
rect 361954 265156 361982 273805
rect 362050 273499 362078 277870
rect 362134 276823 362186 276829
rect 362134 276765 362186 276771
rect 362038 273493 362090 273499
rect 362038 273435 362090 273441
rect 361344 265128 361598 265156
rect 361824 265128 361982 265156
rect 362146 265156 362174 276765
rect 363202 275719 363230 277870
rect 364450 276681 364478 277870
rect 365410 277856 365616 277884
rect 364438 276675 364490 276681
rect 364438 276617 364490 276623
rect 365014 276453 365066 276459
rect 365014 276395 365066 276401
rect 363190 275713 363242 275719
rect 363190 275655 363242 275661
rect 364246 275713 364298 275719
rect 364246 275655 364298 275661
rect 362710 274825 362762 274831
rect 362710 274767 362762 274773
rect 362722 270539 362750 274767
rect 363010 273129 363422 273148
rect 362998 273123 363434 273129
rect 363050 273120 363382 273123
rect 362998 273065 363050 273071
rect 363382 273065 363434 273071
rect 362902 273049 362954 273055
rect 362954 273009 363230 273037
rect 362902 272991 362954 272997
rect 363202 272981 363230 273009
rect 363190 272975 363242 272981
rect 363190 272917 363242 272923
rect 362998 271495 363050 271501
rect 362998 271437 363050 271443
rect 363010 271057 363038 271437
rect 363764 271386 363820 271395
rect 363764 271321 363820 271330
rect 362998 271051 363050 271057
rect 362998 270993 363050 270999
rect 363094 271051 363146 271057
rect 363094 270993 363146 270999
rect 362710 270533 362762 270539
rect 362710 270475 362762 270481
rect 362710 268905 362762 268911
rect 362710 268847 362762 268853
rect 362146 265128 362256 265156
rect 362722 265142 362750 268847
rect 363106 265142 363134 270993
rect 363778 265156 363806 271321
rect 364150 270755 364202 270761
rect 364150 270697 364202 270703
rect 364162 270169 364190 270697
rect 364150 270163 364202 270169
rect 364150 270105 364202 270111
rect 364258 265156 364286 275655
rect 365026 271131 365054 276395
rect 365410 271501 365438 277856
rect 365878 276971 365930 276977
rect 365878 276913 365930 276919
rect 365398 271495 365450 271501
rect 365398 271437 365450 271443
rect 365014 271125 365066 271131
rect 365014 271067 365066 271073
rect 365206 270533 365258 270539
rect 365206 270475 365258 270481
rect 364342 270163 364394 270169
rect 364342 270105 364394 270111
rect 363552 265128 363806 265156
rect 364032 265128 364286 265156
rect 364354 265142 364382 270105
rect 365218 269725 365246 270475
rect 365206 269719 365258 269725
rect 365206 269661 365258 269667
rect 365302 269719 365354 269725
rect 365302 269661 365354 269667
rect 365314 265142 365342 269661
rect 365890 265156 365918 276913
rect 366166 267203 366218 267209
rect 366166 267145 366218 267151
rect 366178 266821 366206 267145
rect 366370 267135 366398 278393
rect 371362 278013 371568 278032
rect 371350 278007 371568 278013
rect 371402 278004 371568 278007
rect 371926 278007 371978 278013
rect 371350 277949 371402 277955
rect 371926 277949 371978 277955
rect 366754 269133 366782 277870
rect 366850 277856 367920 277884
rect 366742 269127 366794 269133
rect 366742 269069 366794 269075
rect 366850 269004 366878 277856
rect 368278 277563 368330 277569
rect 368278 277505 368330 277511
rect 367510 276157 367562 276163
rect 367510 276099 367562 276105
rect 367030 271125 367082 271131
rect 367030 271067 367082 271073
rect 366466 268976 366878 269004
rect 366466 267431 366494 268976
rect 366742 267721 366794 267727
rect 366742 267663 366794 267669
rect 366838 267721 366890 267727
rect 366838 267663 366890 267669
rect 366646 267647 366698 267653
rect 366646 267589 366698 267595
rect 366658 267505 366686 267589
rect 366646 267499 366698 267505
rect 366646 267441 366698 267447
rect 366454 267425 366506 267431
rect 366454 267367 366506 267373
rect 366754 267357 366782 267663
rect 366742 267351 366794 267357
rect 366742 267293 366794 267299
rect 366850 267228 366878 267663
rect 366934 267647 366986 267653
rect 366934 267589 366986 267595
rect 366466 267200 366878 267228
rect 366358 267129 366410 267135
rect 366358 267071 366410 267077
rect 366262 267055 366314 267061
rect 366262 266997 366314 267003
rect 366274 266932 366302 266997
rect 366466 266932 366494 267200
rect 366274 266904 366494 266932
rect 366550 266981 366602 266987
rect 366550 266923 366602 266929
rect 366562 266821 366590 266923
rect 366178 266793 366590 266821
rect 366454 266315 366506 266321
rect 366454 266257 366506 266263
rect 366466 265156 366494 266257
rect 366946 265156 366974 267589
rect 365760 265128 365918 265156
rect 366144 265128 366494 265156
rect 366576 265128 366974 265156
rect 367042 265142 367070 271067
rect 367318 269127 367370 269133
rect 367318 269069 367370 269075
rect 367330 266321 367358 269069
rect 367414 267425 367466 267431
rect 367414 267367 367466 267373
rect 367426 266691 367454 267367
rect 367414 266685 367466 266691
rect 367414 266627 367466 266633
rect 367414 266537 367466 266543
rect 367414 266479 367466 266485
rect 367426 266321 367454 266479
rect 367318 266315 367370 266321
rect 367318 266257 367370 266263
rect 367414 266315 367466 266321
rect 367414 266257 367466 266263
rect 367522 265142 367550 276099
rect 368086 276009 368138 276015
rect 368086 275951 368138 275957
rect 367894 267499 367946 267505
rect 367894 267441 367946 267447
rect 367906 267135 367934 267441
rect 367990 267277 368042 267283
rect 367990 267219 368042 267225
rect 367894 267129 367946 267135
rect 367894 267071 367946 267077
rect 368002 267061 368030 267219
rect 367990 267055 368042 267061
rect 367990 266997 368042 267003
rect 367606 266981 367658 266987
rect 367606 266923 367658 266929
rect 367618 266691 367646 266923
rect 367606 266685 367658 266691
rect 367606 266627 367658 266633
rect 367606 266537 367658 266543
rect 367606 266479 367658 266485
rect 349846 265073 349898 265079
rect 367618 265063 367646 266479
rect 368098 265156 368126 275951
rect 368180 271090 368236 271099
rect 368180 271025 368236 271034
rect 368194 268139 368222 271025
rect 368180 268130 368236 268139
rect 368180 268065 368236 268074
rect 368182 267499 368234 267505
rect 368182 267441 368234 267447
rect 368194 267357 368222 267441
rect 368182 267351 368234 267357
rect 368182 267293 368234 267299
rect 368290 265304 368318 277505
rect 369154 276459 369182 277870
rect 369142 276453 369194 276459
rect 369142 276395 369194 276401
rect 370306 275645 370334 277870
rect 371350 276453 371402 276459
rect 371350 276395 371402 276401
rect 370294 275639 370346 275645
rect 370294 275581 370346 275587
rect 370004 274938 370060 274947
rect 370004 274873 370060 274882
rect 368468 274790 368524 274799
rect 368468 274725 368524 274734
rect 368482 274313 368510 274725
rect 368470 274307 368522 274313
rect 368470 274249 368522 274255
rect 368854 274307 368906 274313
rect 368854 274249 368906 274255
rect 369622 274307 369674 274313
rect 369622 274249 369674 274255
rect 368662 273493 368714 273499
rect 368662 273435 368714 273441
rect 368674 272727 368702 273435
rect 368866 272727 368894 274249
rect 369142 273493 369194 273499
rect 369140 273458 369142 273467
rect 369194 273458 369196 273467
rect 369140 273393 369196 273402
rect 368660 272718 368716 272727
rect 368660 272653 368716 272662
rect 368852 272718 368908 272727
rect 368852 272653 368908 272662
rect 368482 270937 368990 270965
rect 368372 270794 368428 270803
rect 368372 270729 368428 270738
rect 368386 268287 368414 270729
rect 368482 270539 368510 270937
rect 368578 270863 368894 270891
rect 368470 270533 368522 270539
rect 368470 270475 368522 270481
rect 368578 270465 368606 270863
rect 368756 270794 368812 270803
rect 368756 270729 368812 270738
rect 368566 270459 368618 270465
rect 368566 270401 368618 270407
rect 368770 269767 368798 270729
rect 368866 270465 368894 270863
rect 368962 270803 368990 270937
rect 368948 270794 369004 270803
rect 368948 270729 369004 270738
rect 369046 270755 369098 270761
rect 369046 270697 369098 270703
rect 369058 270669 369086 270697
rect 369238 270681 369290 270687
rect 369058 270641 369238 270669
rect 369238 270623 369290 270629
rect 368854 270459 368906 270465
rect 368854 270401 368906 270407
rect 369046 270311 369098 270317
rect 368866 270271 369046 270299
rect 368564 269758 368620 269767
rect 368564 269693 368620 269702
rect 368756 269758 368812 269767
rect 368756 269693 368812 269702
rect 368578 269596 368606 269693
rect 368866 269596 368894 270271
rect 369046 270253 369098 270259
rect 368578 269568 368894 269596
rect 368662 268609 368714 268615
rect 368714 268569 368990 268597
rect 368662 268551 368714 268557
rect 368854 268535 368906 268541
rect 368854 268477 368906 268483
rect 368372 268278 368428 268287
rect 368372 268213 368428 268222
rect 368756 268130 368812 268139
rect 368756 268065 368812 268074
rect 368770 267949 368798 268065
rect 368866 268023 368894 268477
rect 368962 268023 368990 268569
rect 369236 268278 369292 268287
rect 369236 268213 369292 268222
rect 369250 268171 369278 268213
rect 369238 268165 369290 268171
rect 369238 268107 369290 268113
rect 368854 268017 368906 268023
rect 368854 267959 368906 267965
rect 368950 268017 369002 268023
rect 368950 267959 369002 267965
rect 368758 267943 368810 267949
rect 368758 267885 368810 267891
rect 369334 267721 369386 267727
rect 369334 267663 369386 267669
rect 368470 267351 368522 267357
rect 368470 267293 368522 267299
rect 368374 267277 368426 267283
rect 368374 267219 368426 267225
rect 368386 266659 368414 267219
rect 368482 266955 368510 267293
rect 368758 267277 368810 267283
rect 368758 267219 368810 267225
rect 369046 267277 369098 267283
rect 369046 267219 369098 267225
rect 368770 267103 368798 267219
rect 368756 267094 368812 267103
rect 368756 267029 368812 267038
rect 368468 266946 368524 266955
rect 368660 266946 368716 266955
rect 368468 266881 368524 266890
rect 368578 266904 368660 266932
rect 368372 266650 368428 266659
rect 368372 266585 368428 266594
rect 367872 265128 368126 265156
rect 368194 265276 368318 265304
rect 356854 265057 356906 265063
rect 356592 265005 356854 265008
rect 367606 265057 367658 265063
rect 356592 264999 356906 265005
rect 347734 264983 347786 264989
rect 356592 264980 356894 264999
rect 364848 264994 365054 265008
rect 367606 264999 367658 265005
rect 364848 264985 365068 264994
rect 364848 264980 365012 264985
rect 347734 264925 347786 264931
rect 365012 264920 365068 264929
rect 343702 264909 343754 264915
rect 328354 264832 328704 264860
rect 343702 264851 343754 264857
rect 368194 264860 368222 265276
rect 368578 265063 368606 266904
rect 368660 266881 368716 266890
rect 369058 265156 369086 267219
rect 369346 266839 369374 267663
rect 369142 266833 369194 266839
rect 369142 266775 369194 266781
rect 369334 266833 369386 266839
rect 369334 266775 369386 266781
rect 368784 265128 369086 265156
rect 369154 265063 369182 266775
rect 369634 265142 369662 274249
rect 370018 273499 370046 274873
rect 370388 274790 370444 274799
rect 370388 274725 370444 274734
rect 370402 273795 370430 274725
rect 370966 273937 371018 273943
rect 370966 273879 371018 273885
rect 370390 273789 370442 273795
rect 370390 273731 370442 273737
rect 370006 273493 370058 273499
rect 370006 273435 370058 273441
rect 370390 272827 370442 272833
rect 370390 272769 370442 272775
rect 370402 272315 370430 272769
rect 370390 272309 370442 272315
rect 370390 272251 370442 272257
rect 370198 272235 370250 272241
rect 370198 272177 370250 272183
rect 370006 271495 370058 271501
rect 370006 271437 370058 271443
rect 370018 271205 370046 271437
rect 370210 271279 370238 272177
rect 370978 271543 371006 273879
rect 370964 271534 371020 271543
rect 370964 271469 371020 271478
rect 370580 271386 370636 271395
rect 370580 271321 370636 271330
rect 370198 271273 370250 271279
rect 370198 271215 370250 271221
rect 370006 271199 370058 271205
rect 370006 271141 370058 271147
rect 369812 271090 369868 271099
rect 369812 271025 369868 271034
rect 369826 270507 369854 271025
rect 369812 270498 369868 270507
rect 369812 270433 369868 270442
rect 370004 270498 370060 270507
rect 370004 270433 370060 270442
rect 370018 270095 370046 270433
rect 370006 270089 370058 270095
rect 370006 270031 370058 270037
rect 370198 270089 370250 270095
rect 370198 270031 370250 270037
rect 370210 268615 370238 270031
rect 370198 268609 370250 268615
rect 370198 268551 370250 268557
rect 370294 268609 370346 268615
rect 370594 268583 370622 271321
rect 370294 268551 370346 268557
rect 370580 268574 370636 268583
rect 370306 265156 370334 268551
rect 370580 268509 370636 268518
rect 370772 268574 370828 268583
rect 370772 268509 370828 268518
rect 370786 265156 370814 268509
rect 370966 267943 371018 267949
rect 370966 267885 371018 267891
rect 370080 265128 370334 265156
rect 370560 265128 370814 265156
rect 370978 265142 371006 267885
rect 371362 265142 371390 276395
rect 371444 271534 371500 271543
rect 371444 271469 371500 271478
rect 371458 270951 371486 271469
rect 371938 271131 371966 277949
rect 372514 276385 372542 278467
rect 372502 276379 372554 276385
rect 372502 276321 372554 276327
rect 372404 274642 372460 274651
rect 372404 274577 372460 274586
rect 372418 273721 372446 274577
rect 372406 273715 372458 273721
rect 372406 273657 372458 273663
rect 372502 273715 372554 273721
rect 372502 273657 372554 273663
rect 371926 271125 371978 271131
rect 371926 271067 371978 271073
rect 371444 270942 371500 270951
rect 371444 270877 371500 270886
rect 371444 268574 371500 268583
rect 371444 268509 371500 268518
rect 371458 268097 371486 268509
rect 371830 268165 371882 268171
rect 371830 268107 371882 268113
rect 371446 268091 371498 268097
rect 371446 268033 371498 268039
rect 371842 265142 371870 268107
rect 372514 265156 372542 273657
rect 372706 273277 372734 277870
rect 373474 277856 373872 277884
rect 372982 276675 373034 276681
rect 372982 276617 373034 276623
rect 372994 275719 373022 276617
rect 372982 275713 373034 275719
rect 372982 275655 373034 275661
rect 373366 273789 373418 273795
rect 373366 273731 373418 273737
rect 372694 273271 372746 273277
rect 372694 273213 372746 273219
rect 373078 272827 373130 272833
rect 373078 272769 373130 272775
rect 373090 272463 373118 272769
rect 373078 272457 373130 272463
rect 373078 272399 373130 272405
rect 373174 272457 373226 272463
rect 373174 272399 373226 272405
rect 372886 271125 372938 271131
rect 372886 271067 372938 271073
rect 372898 270835 372926 271067
rect 372886 270829 372938 270835
rect 372886 270771 372938 270777
rect 372982 270829 373034 270835
rect 373186 270803 373214 272399
rect 372982 270771 373034 270777
rect 373172 270794 373228 270803
rect 372694 268091 372746 268097
rect 372694 268033 372746 268039
rect 372706 267843 372734 268033
rect 372692 267834 372748 267843
rect 372692 267769 372748 267778
rect 372886 267647 372938 267653
rect 372886 267589 372938 267595
rect 372898 265156 372926 267589
rect 372288 265128 372542 265156
rect 372672 265128 372926 265156
rect 372994 265137 373022 270771
rect 373172 270729 373228 270738
rect 373378 265156 373406 273731
rect 373474 270761 373502 277856
rect 374146 276459 374174 278596
rect 395060 278638 395116 278647
rect 374324 278573 374380 278582
rect 380194 278596 380414 278624
rect 393826 278605 394128 278624
rect 374614 278525 374666 278531
rect 374614 278467 374666 278473
rect 374710 278525 374762 278531
rect 374710 278467 374762 278473
rect 374326 276527 374378 276533
rect 374326 276469 374378 276475
rect 374134 276453 374186 276459
rect 374134 276395 374186 276401
rect 374230 276453 374282 276459
rect 374230 276395 374282 276401
rect 374038 275713 374090 275719
rect 374038 275655 374090 275661
rect 373556 270794 373612 270803
rect 373462 270755 373514 270761
rect 373556 270729 373612 270738
rect 373462 270697 373514 270703
rect 372982 265131 373034 265137
rect 373152 265128 373406 265156
rect 373570 265142 373598 270729
rect 374050 265142 374078 275655
rect 374242 268023 374270 276395
rect 374338 275867 374366 276469
rect 374626 275867 374654 278467
rect 374722 276385 374750 278467
rect 378370 278457 378672 278476
rect 380194 278457 380222 278596
rect 378358 278451 378672 278457
rect 378410 278448 378672 278451
rect 380182 278451 380234 278457
rect 378358 278393 378410 278399
rect 380182 278393 380234 278399
rect 380278 278451 380330 278457
rect 380278 278393 380330 278399
rect 374806 278377 374858 278383
rect 375286 278377 375338 278383
rect 374858 278325 375120 278328
rect 374806 278319 375120 278325
rect 375286 278319 375338 278325
rect 378550 278377 378602 278383
rect 378550 278319 378602 278325
rect 374818 278300 375120 278319
rect 375298 277736 375326 278319
rect 375202 277708 375326 277736
rect 375202 277569 375230 277708
rect 375190 277563 375242 277569
rect 375190 277505 375242 277511
rect 375286 277563 375338 277569
rect 375286 277505 375338 277511
rect 375188 276862 375244 276871
rect 375188 276797 375244 276806
rect 375202 276755 375230 276797
rect 375190 276749 375242 276755
rect 375298 276723 375326 277505
rect 375380 276862 375436 276871
rect 375380 276797 375436 276806
rect 375190 276691 375242 276697
rect 375284 276714 375340 276723
rect 375284 276649 375340 276658
rect 374710 276379 374762 276385
rect 374710 276321 374762 276327
rect 375394 276163 375422 276797
rect 375476 276714 375532 276723
rect 375476 276649 375532 276658
rect 375490 276459 375518 276649
rect 375478 276453 375530 276459
rect 375478 276395 375530 276401
rect 375670 276453 375722 276459
rect 375670 276395 375722 276401
rect 375574 276379 375626 276385
rect 375574 276321 375626 276327
rect 375382 276157 375434 276163
rect 375382 276099 375434 276105
rect 374326 275861 374378 275867
rect 374326 275803 374378 275809
rect 374614 275861 374666 275867
rect 374614 275803 374666 275809
rect 375586 274461 375614 276321
rect 375682 276015 375710 276395
rect 375670 276009 375722 276015
rect 375670 275951 375722 275957
rect 375766 276009 375818 276015
rect 375766 275951 375818 275957
rect 375778 274831 375806 275951
rect 375766 274825 375818 274831
rect 375766 274767 375818 274773
rect 375574 274455 375626 274461
rect 375574 274397 375626 274403
rect 375766 274455 375818 274461
rect 375766 274397 375818 274403
rect 374422 273271 374474 273277
rect 374422 273213 374474 273219
rect 374434 271797 374462 273213
rect 374996 272274 375052 272283
rect 374530 272232 374996 272260
rect 374530 271987 374558 272232
rect 374996 272209 375052 272218
rect 374516 271978 374572 271987
rect 374516 271913 374572 271922
rect 374422 271791 374474 271797
rect 374422 271733 374474 271739
rect 375574 271791 375626 271797
rect 375574 271733 375626 271739
rect 374998 270755 375050 270761
rect 374998 270697 375050 270703
rect 375010 270095 375038 270697
rect 374998 270089 375050 270095
rect 374998 270031 375050 270037
rect 375094 270089 375146 270095
rect 375094 270031 375146 270037
rect 374230 268017 374282 268023
rect 374230 267959 374282 267965
rect 374710 268017 374762 268023
rect 374710 267959 374762 267965
rect 374146 267311 374558 267339
rect 374146 267251 374174 267311
rect 374422 267277 374474 267283
rect 374132 267242 374188 267251
rect 374420 267242 374422 267251
rect 374474 267242 374476 267251
rect 374132 267177 374188 267186
rect 374230 267203 374282 267209
rect 374530 267228 374558 267311
rect 374612 267242 374668 267251
rect 374530 267200 374612 267228
rect 374420 267177 374476 267186
rect 374612 267177 374668 267186
rect 374230 267145 374282 267151
rect 374242 267117 374270 267145
rect 374422 267129 374474 267135
rect 374242 267089 374422 267117
rect 374422 267071 374474 267077
rect 374722 265156 374750 267959
rect 374806 267277 374858 267283
rect 374806 267219 374858 267225
rect 374818 267135 374846 267219
rect 374806 267129 374858 267135
rect 374806 267071 374858 267077
rect 375106 265156 375134 270031
rect 375586 265156 375614 271733
rect 374448 265128 374750 265156
rect 374880 265128 375134 265156
rect 375360 265128 375614 265156
rect 375778 265142 375806 274397
rect 376258 273277 376286 277870
rect 376342 276157 376394 276163
rect 376342 276099 376394 276105
rect 376354 274387 376382 276099
rect 377506 275349 377534 277870
rect 378562 276108 378590 278319
rect 377698 276080 378590 276108
rect 377494 275343 377546 275349
rect 377494 275285 377546 275291
rect 377590 275343 377642 275349
rect 377590 275285 377642 275291
rect 377602 274461 377630 275285
rect 377590 274455 377642 274461
rect 377590 274397 377642 274403
rect 376342 274381 376394 274387
rect 376342 274323 376394 274329
rect 377302 274381 377354 274387
rect 377302 274323 377354 274329
rect 376246 273271 376298 273277
rect 376246 273213 376298 273219
rect 376342 273271 376394 273277
rect 376342 273213 376394 273219
rect 376354 273171 376382 273213
rect 376340 273162 376396 273171
rect 376340 273097 376396 273106
rect 376532 273162 376588 273171
rect 376532 273097 376588 273106
rect 376546 265156 376574 273097
rect 376628 270942 376684 270951
rect 376628 270877 376684 270886
rect 376642 267949 376670 270877
rect 377110 268239 377162 268245
rect 377110 268181 377162 268187
rect 377122 267991 377150 268181
rect 377108 267982 377164 267991
rect 376630 267943 376682 267949
rect 377108 267917 377164 267926
rect 377206 267943 377258 267949
rect 376630 267885 376682 267891
rect 377206 267885 377258 267891
rect 376820 267834 376876 267843
rect 376820 267769 376876 267778
rect 376834 267547 376862 267769
rect 377218 267653 377246 267885
rect 377206 267647 377258 267653
rect 377206 267589 377258 267595
rect 377110 267573 377162 267579
rect 376820 267538 376876 267547
rect 377110 267515 377162 267521
rect 376820 267473 376876 267482
rect 377122 267283 377150 267515
rect 377110 267277 377162 267283
rect 377110 267219 377162 267225
rect 377314 265156 377342 274323
rect 377698 273721 377726 276080
rect 379906 276015 379934 277870
rect 380290 277347 380318 278393
rect 380386 277347 380414 278596
rect 384406 278599 384458 278605
rect 384406 278541 384458 278547
rect 393814 278599 394128 278605
rect 393866 278596 394128 278599
rect 432240 278605 432446 278624
rect 395060 278573 395116 278582
rect 407542 278599 407594 278605
rect 393814 278541 393866 278547
rect 384418 278235 384446 278541
rect 384694 278377 384746 278383
rect 384694 278319 384746 278325
rect 382006 278229 382058 278235
rect 382390 278229 382442 278235
rect 382058 278177 382320 278180
rect 382006 278171 382320 278177
rect 382390 278171 382442 278177
rect 384022 278229 384074 278235
rect 384022 278171 384074 278177
rect 384406 278229 384458 278235
rect 384406 278171 384458 278177
rect 382018 278152 382320 278171
rect 380482 277856 381072 277884
rect 380278 277341 380330 277347
rect 380278 277283 380330 277289
rect 380374 277341 380426 277347
rect 380374 277283 380426 277289
rect 379990 276749 380042 276755
rect 379990 276691 380042 276697
rect 380086 276749 380138 276755
rect 380086 276691 380138 276697
rect 380002 276015 380030 276691
rect 379894 276009 379946 276015
rect 377986 275932 378206 275960
rect 379894 275951 379946 275957
rect 379990 276009 380042 276015
rect 379990 275951 380042 275957
rect 377986 275867 378014 275932
rect 377974 275861 378026 275867
rect 377974 275803 378026 275809
rect 378070 275861 378122 275867
rect 378070 275803 378122 275809
rect 377782 275639 377834 275645
rect 377782 275581 377834 275587
rect 377686 273715 377738 273721
rect 377686 273657 377738 273663
rect 377794 270835 377822 275581
rect 377878 274825 377930 274831
rect 377878 274767 377930 274773
rect 377890 274313 377918 274767
rect 377878 274307 377930 274313
rect 377878 274249 377930 274255
rect 377974 274307 378026 274313
rect 377974 274249 378026 274255
rect 377986 273615 378014 274249
rect 378082 273795 378110 275803
rect 378178 275368 378206 275932
rect 378178 275340 379262 275368
rect 378836 274938 378892 274947
rect 378836 274873 378892 274882
rect 378550 274381 378602 274387
rect 378550 274323 378602 274329
rect 378070 273789 378122 273795
rect 378070 273731 378122 273737
rect 378166 273789 378218 273795
rect 378166 273731 378218 273737
rect 378178 273615 378206 273731
rect 377972 273606 378028 273615
rect 377972 273541 378028 273550
rect 378164 273606 378220 273615
rect 378164 273541 378220 273550
rect 377986 273425 378398 273444
rect 377974 273419 378410 273425
rect 378026 273416 378358 273419
rect 377974 273361 378026 273367
rect 378562 273407 378590 274323
rect 378850 273721 378878 274873
rect 379234 274461 379262 275340
rect 379126 274455 379178 274461
rect 379126 274397 379178 274403
rect 379222 274455 379274 274461
rect 379222 274397 379274 274403
rect 378838 273715 378890 273721
rect 378838 273657 378890 273663
rect 378934 273715 378986 273721
rect 378934 273657 378986 273663
rect 378646 273641 378698 273647
rect 378646 273583 378698 273589
rect 378658 273499 378686 273583
rect 378646 273493 378698 273499
rect 378646 273435 378698 273441
rect 378358 273361 378410 273367
rect 378466 273379 378590 273407
rect 378466 273296 378494 273379
rect 378370 273268 378494 273296
rect 378370 273259 378398 273268
rect 378274 273231 378398 273259
rect 378274 272963 378302 273231
rect 378358 273197 378410 273203
rect 378742 273197 378794 273203
rect 378358 273139 378410 273145
rect 378562 273157 378742 273185
rect 377890 272935 378302 272963
rect 377782 270829 377834 270835
rect 377782 270771 377834 270777
rect 377590 268905 377642 268911
rect 377590 268847 377642 268853
rect 377396 267982 377452 267991
rect 377396 267917 377452 267926
rect 377410 267357 377438 267917
rect 377494 267721 377546 267727
rect 377494 267663 377546 267669
rect 377398 267351 377450 267357
rect 377398 267293 377450 267299
rect 377506 267135 377534 267663
rect 377602 267431 377630 268847
rect 377590 267425 377642 267431
rect 377590 267367 377642 267373
rect 377494 267129 377546 267135
rect 377494 267071 377546 267077
rect 377686 267129 377738 267135
rect 377686 267071 377738 267077
rect 377698 266617 377726 267071
rect 377890 266969 377918 272935
rect 378166 272901 378218 272907
rect 378218 272861 378302 272889
rect 378166 272843 378218 272849
rect 377974 272679 378026 272685
rect 377974 272621 378026 272627
rect 377986 272445 378014 272621
rect 378274 272593 378302 272861
rect 378370 272685 378398 273139
rect 378562 272759 378590 273157
rect 378742 273139 378794 273145
rect 378946 273023 378974 273657
rect 379138 273647 379166 274397
rect 380098 274036 380126 276691
rect 380482 275701 380510 277856
rect 382402 276848 382430 278171
rect 381154 276820 382430 276848
rect 382978 277856 383376 277884
rect 381154 276755 381182 276820
rect 381142 276749 381194 276755
rect 381142 276691 381194 276697
rect 381238 276749 381290 276755
rect 381238 276691 381290 276697
rect 380002 274008 380126 274036
rect 380290 275673 380510 275701
rect 379702 273715 379754 273721
rect 379702 273657 379754 273663
rect 379030 273641 379082 273647
rect 379030 273583 379082 273589
rect 379126 273641 379178 273647
rect 379714 273615 379742 273657
rect 379126 273583 379178 273589
rect 379700 273606 379756 273615
rect 379042 273319 379070 273583
rect 379700 273541 379756 273550
rect 379126 273493 379178 273499
rect 379126 273435 379178 273441
rect 379220 273458 379276 273467
rect 379028 273310 379084 273319
rect 379028 273245 379084 273254
rect 378932 273014 378988 273023
rect 378742 272975 378794 272981
rect 378932 272949 378988 272958
rect 378742 272917 378794 272923
rect 378754 272889 378782 272917
rect 378658 272861 378782 272889
rect 378934 272901 378986 272907
rect 378550 272753 378602 272759
rect 378550 272695 378602 272701
rect 378358 272679 378410 272685
rect 378358 272621 378410 272627
rect 378658 272611 378686 272861
rect 378934 272843 378986 272849
rect 378838 272679 378890 272685
rect 378838 272621 378890 272627
rect 378646 272605 378698 272611
rect 378274 272565 378494 272593
rect 378358 272457 378410 272463
rect 377986 272417 378206 272445
rect 378178 271797 378206 272417
rect 378358 272399 378410 272405
rect 378370 271964 378398 272399
rect 378466 272149 378494 272565
rect 378646 272547 378698 272553
rect 378850 272519 378878 272621
rect 378562 272491 378878 272519
rect 378562 272241 378590 272491
rect 378946 272241 378974 272843
rect 379138 272593 379166 273435
rect 379412 273458 379468 273467
rect 379220 273393 379276 273402
rect 379330 273416 379412 273444
rect 379234 273023 379262 273393
rect 379330 273277 379358 273416
rect 379412 273393 379468 273402
rect 379318 273271 379370 273277
rect 379318 273213 379370 273219
rect 379414 273271 379466 273277
rect 379414 273213 379466 273219
rect 379316 273162 379372 273171
rect 379316 273097 379372 273106
rect 379220 273014 379276 273023
rect 379220 272949 379276 272958
rect 379330 272907 379358 273097
rect 379318 272901 379370 272907
rect 379318 272843 379370 272849
rect 379042 272565 379166 272593
rect 379042 272537 379070 272565
rect 379030 272531 379082 272537
rect 379318 272531 379370 272537
rect 379030 272473 379082 272479
rect 379138 272491 379318 272519
rect 378550 272235 378602 272241
rect 378550 272177 378602 272183
rect 378646 272235 378698 272241
rect 378646 272177 378698 272183
rect 378934 272235 378986 272241
rect 378934 272177 378986 272183
rect 378658 272149 378686 272177
rect 379138 272167 379166 272491
rect 379318 272473 379370 272479
rect 379316 272274 379372 272283
rect 379316 272209 379372 272218
rect 378466 272121 378686 272149
rect 379126 272161 379178 272167
rect 379126 272103 379178 272109
rect 378370 271936 379070 271964
rect 378070 271791 378122 271797
rect 378070 271733 378122 271739
rect 378166 271791 378218 271797
rect 378166 271733 378218 271739
rect 378082 271057 378110 271733
rect 377974 271051 378026 271057
rect 377974 270993 378026 270999
rect 378070 271051 378122 271057
rect 378934 271051 378986 271057
rect 378070 270993 378122 270999
rect 378754 271011 378934 271039
rect 377794 266941 377918 266969
rect 377686 266611 377738 266617
rect 377686 266553 377738 266559
rect 377794 265156 377822 266941
rect 377986 266913 378014 270993
rect 378178 270604 378686 270632
rect 378178 270169 378206 270604
rect 378658 270539 378686 270604
rect 378550 270533 378602 270539
rect 378550 270475 378602 270481
rect 378646 270533 378698 270539
rect 378646 270475 378698 270481
rect 378166 270163 378218 270169
rect 378166 270105 378218 270111
rect 378562 270095 378590 270475
rect 378550 270089 378602 270095
rect 378550 270031 378602 270037
rect 378754 269596 378782 271011
rect 378934 270993 378986 270999
rect 379042 270965 379070 271936
rect 379330 271691 379358 272209
rect 379316 271682 379372 271691
rect 379316 271617 379372 271626
rect 379426 271057 379454 273213
rect 379510 273049 379562 273055
rect 379510 272991 379562 272997
rect 379606 273049 379658 273055
rect 379606 272991 379658 272997
rect 379522 272315 379550 272991
rect 379510 272309 379562 272315
rect 379510 272251 379562 272257
rect 379414 271051 379466 271057
rect 379414 270993 379466 270999
rect 379510 271051 379562 271057
rect 379510 270993 379562 270999
rect 379522 270965 379550 270993
rect 379042 270937 379550 270965
rect 378178 269568 378782 269596
rect 378178 267635 378206 269568
rect 378550 269497 378602 269503
rect 378550 269439 378602 269445
rect 378646 269497 378698 269503
rect 378646 269439 378698 269445
rect 378358 268905 378410 268911
rect 378358 268847 378410 268853
rect 378082 267607 378206 267635
rect 377878 266907 377930 266913
rect 377878 266849 377930 266855
rect 377974 266907 378026 266913
rect 377974 266849 378026 266855
rect 377890 266617 377918 266849
rect 377878 266611 377930 266617
rect 377878 266553 377930 266559
rect 378082 265156 378110 267607
rect 376176 265128 376574 265156
rect 376656 265137 376958 265156
rect 376656 265131 376970 265137
rect 376656 265128 376918 265131
rect 372982 265073 373034 265079
rect 377088 265128 377342 265156
rect 377568 265128 377822 265156
rect 377904 265128 378110 265156
rect 378370 265142 378398 268847
rect 378562 268227 378590 269439
rect 378658 269133 378686 269439
rect 378646 269127 378698 269133
rect 378646 269069 378698 269075
rect 378742 269127 378794 269133
rect 378742 269069 378794 269075
rect 378754 268615 378782 269069
rect 378742 268609 378794 268615
rect 378742 268551 378794 268557
rect 378838 268609 378890 268615
rect 378838 268551 378890 268557
rect 378646 268239 378698 268245
rect 378562 268199 378646 268227
rect 378646 268181 378698 268187
rect 378850 268023 378878 268551
rect 378838 268017 378890 268023
rect 378838 267959 378890 267965
rect 379222 268017 379274 268023
rect 379222 267959 379274 267965
rect 378742 267647 378794 267653
rect 378742 267589 378794 267595
rect 378754 267547 378782 267589
rect 378740 267538 378796 267547
rect 378740 267473 378796 267482
rect 378934 267425 378986 267431
rect 378934 267367 378986 267373
rect 378550 267351 378602 267357
rect 378550 267293 378602 267299
rect 378562 266617 378590 267293
rect 378946 267080 378974 267367
rect 378754 267052 378974 267080
rect 378754 266765 378782 267052
rect 379234 266932 379262 267959
rect 378850 266904 379262 266932
rect 378742 266759 378794 266765
rect 378742 266701 378794 266707
rect 378454 266611 378506 266617
rect 378454 266553 378506 266559
rect 378550 266611 378602 266617
rect 378550 266553 378602 266559
rect 378466 266525 378494 266553
rect 378850 266525 378878 266904
rect 379030 266833 379082 266839
rect 379030 266775 379082 266781
rect 378466 266497 378878 266525
rect 379042 265600 379070 266775
rect 378658 265572 379070 265600
rect 376918 265073 376970 265079
rect 378658 265063 378686 265572
rect 379618 265304 379646 272991
rect 379798 272457 379850 272463
rect 379798 272399 379850 272405
rect 379810 272283 379838 272399
rect 379796 272274 379852 272283
rect 379796 272209 379852 272218
rect 379714 271085 379934 271113
rect 379714 269725 379742 271085
rect 379906 271057 379934 271085
rect 379798 271051 379850 271057
rect 379798 270993 379850 270999
rect 379894 271051 379946 271057
rect 379894 270993 379946 270999
rect 379810 269725 379838 270993
rect 379702 269719 379754 269725
rect 379702 269661 379754 269667
rect 379798 269719 379850 269725
rect 379798 269661 379850 269667
rect 380002 268745 380030 274008
rect 380290 273740 380318 275673
rect 381250 274184 381278 276691
rect 380674 274156 381278 274184
rect 380086 273715 380138 273721
rect 380290 273712 380414 273740
rect 380086 273657 380138 273663
rect 380098 271057 380126 273657
rect 380180 272274 380236 272283
rect 380180 272209 380236 272218
rect 380086 271051 380138 271057
rect 380086 270993 380138 270999
rect 380086 270089 380138 270095
rect 380086 270031 380138 270037
rect 379138 265276 379646 265304
rect 379810 268717 380030 268745
rect 379138 265156 379166 265276
rect 379810 265156 379838 268717
rect 379894 268683 379946 268689
rect 379894 268625 379946 268631
rect 379906 268153 379934 268625
rect 380098 268227 380126 270031
rect 380194 269767 380222 272209
rect 380278 271051 380330 271057
rect 380278 270993 380330 270999
rect 380290 270169 380318 270993
rect 380386 270687 380414 273712
rect 380374 270681 380426 270687
rect 380374 270623 380426 270629
rect 380278 270163 380330 270169
rect 380278 270105 380330 270111
rect 380374 270163 380426 270169
rect 380374 270105 380426 270111
rect 380180 269758 380236 269767
rect 380180 269693 380236 269702
rect 380182 269275 380234 269281
rect 380386 269263 380414 270105
rect 380470 270089 380522 270095
rect 380470 270031 380522 270037
rect 380234 269235 380414 269263
rect 380182 269217 380234 269223
rect 380182 268831 380234 268837
rect 380482 268819 380510 270031
rect 380564 269758 380620 269767
rect 380564 269693 380620 269702
rect 380182 268773 380234 268779
rect 380290 268791 380510 268819
rect 380194 268689 380222 268773
rect 380182 268683 380234 268689
rect 380182 268625 380234 268631
rect 380290 268615 380318 268791
rect 380578 268745 380606 269693
rect 380386 268717 380606 268745
rect 380278 268609 380330 268615
rect 380278 268551 380330 268557
rect 380386 268319 380414 268717
rect 380566 268609 380618 268615
rect 380566 268551 380618 268557
rect 380374 268313 380426 268319
rect 380374 268255 380426 268261
rect 380470 268313 380522 268319
rect 380470 268255 380522 268261
rect 380482 268227 380510 268255
rect 380098 268199 380510 268227
rect 379906 268125 380126 268153
rect 380098 267727 380126 268125
rect 380578 268005 380606 268551
rect 380290 267977 380606 268005
rect 380290 267949 380318 267977
rect 380278 267943 380330 267949
rect 380278 267885 380330 267891
rect 380374 267943 380426 267949
rect 380374 267885 380426 267891
rect 379990 267721 380042 267727
rect 379990 267663 380042 267669
rect 380086 267721 380138 267727
rect 380086 267663 380138 267669
rect 380002 267635 380030 267663
rect 380386 267635 380414 267885
rect 380002 267607 380414 267635
rect 380674 265452 380702 274156
rect 381236 273754 381292 273763
rect 381236 273689 381292 273698
rect 380950 271051 381002 271057
rect 380950 270993 381002 270999
rect 380962 270095 380990 270993
rect 381250 270983 381278 273689
rect 381812 273458 381868 273467
rect 381812 273393 381868 273402
rect 381826 272431 381854 273393
rect 381620 272422 381676 272431
rect 381620 272357 381676 272366
rect 381812 272422 381868 272431
rect 381812 272357 381868 272366
rect 381634 272297 381662 272357
rect 381634 272269 381950 272297
rect 381812 272126 381868 272135
rect 381812 272061 381868 272070
rect 381346 271085 381662 271113
rect 381142 270977 381194 270983
rect 381142 270919 381194 270925
rect 381238 270977 381290 270983
rect 381238 270919 381290 270925
rect 381154 270743 381182 270919
rect 381238 270755 381290 270761
rect 381154 270715 381238 270743
rect 381238 270697 381290 270703
rect 381346 270447 381374 271085
rect 381430 271051 381482 271057
rect 381430 270993 381482 270999
rect 381058 270419 381374 270447
rect 381058 270169 381086 270419
rect 381046 270163 381098 270169
rect 381046 270105 381098 270111
rect 381142 270163 381194 270169
rect 381142 270105 381194 270111
rect 380854 270089 380906 270095
rect 380854 270031 380906 270037
rect 380950 270089 381002 270095
rect 380950 270031 381002 270037
rect 380866 269892 380894 270031
rect 381154 269892 381182 270105
rect 380866 269864 381182 269892
rect 381442 269448 381470 270993
rect 381250 269420 381470 269448
rect 380854 268831 380906 268837
rect 380854 268773 380906 268779
rect 380866 268689 380894 268773
rect 381250 268745 381278 269420
rect 381634 269281 381662 271085
rect 381622 269275 381674 269281
rect 381622 269217 381674 269223
rect 381826 269152 381854 272061
rect 381634 269124 381854 269152
rect 381250 268717 381374 268745
rect 380854 268683 380906 268689
rect 381238 268683 381290 268689
rect 380854 268625 380906 268631
rect 380962 268643 381238 268671
rect 380962 265748 380990 268643
rect 381238 268625 381290 268631
rect 380482 265424 380702 265452
rect 380770 265720 380990 265748
rect 380482 265156 380510 265424
rect 380770 265304 380798 265720
rect 381346 265304 381374 268717
rect 380674 265276 380798 265304
rect 381250 265276 381374 265304
rect 380674 265156 380702 265276
rect 381250 265156 381278 265276
rect 381634 265156 381662 269124
rect 381922 265452 381950 272269
rect 382006 270903 382058 270909
rect 382006 270845 382058 270851
rect 378864 265128 379166 265156
rect 379680 265128 379838 265156
rect 380112 265128 380510 265156
rect 380592 265128 380702 265156
rect 380976 265128 381278 265156
rect 381408 265128 381662 265156
rect 381874 265424 381950 265452
rect 381874 265142 381902 265424
rect 382018 265156 382046 270845
rect 382978 267949 383006 277856
rect 383830 277563 383882 277569
rect 383830 277505 383882 277511
rect 383926 277563 383978 277569
rect 383926 277505 383978 277511
rect 383542 276009 383594 276015
rect 383542 275951 383594 275957
rect 383554 273763 383582 275951
rect 383842 274387 383870 277505
rect 383938 276163 383966 277505
rect 384034 276552 384062 278171
rect 384322 277856 384624 277884
rect 384322 277569 384350 277856
rect 384406 277711 384458 277717
rect 384406 277653 384458 277659
rect 384502 277711 384554 277717
rect 384502 277653 384554 277659
rect 384418 277569 384446 277653
rect 384310 277563 384362 277569
rect 384310 277505 384362 277511
rect 384406 277563 384458 277569
rect 384406 277505 384458 277511
rect 384118 277341 384170 277347
rect 384118 277283 384170 277289
rect 384214 277341 384266 277347
rect 384214 277283 384266 277289
rect 384130 276700 384158 277283
rect 384226 277051 384254 277283
rect 384514 277144 384542 277653
rect 384322 277116 384542 277144
rect 384214 277045 384266 277051
rect 384214 276987 384266 276993
rect 384322 276903 384350 277116
rect 384406 277045 384458 277051
rect 384406 276987 384458 276993
rect 384310 276897 384362 276903
rect 384310 276839 384362 276845
rect 384418 276700 384446 276987
rect 384502 276971 384554 276977
rect 384502 276913 384554 276919
rect 384130 276672 384446 276700
rect 384514 276681 384542 276913
rect 384502 276675 384554 276681
rect 384502 276617 384554 276623
rect 384034 276524 384254 276552
rect 384226 276459 384254 276524
rect 384118 276453 384170 276459
rect 384118 276395 384170 276401
rect 384214 276453 384266 276459
rect 384214 276395 384266 276401
rect 383926 276157 383978 276163
rect 383926 276099 383978 276105
rect 384130 275516 384158 276395
rect 384706 276163 384734 278319
rect 385378 277856 385776 277884
rect 384898 276487 385310 276515
rect 384898 276459 384926 276487
rect 384886 276453 384938 276459
rect 384886 276395 384938 276401
rect 385078 276453 385130 276459
rect 385078 276395 385130 276401
rect 384694 276157 384746 276163
rect 384694 276099 384746 276105
rect 384310 276009 384362 276015
rect 384310 275951 384362 275957
rect 384322 275867 384350 275951
rect 384310 275861 384362 275867
rect 384310 275803 384362 275809
rect 384406 275861 384458 275867
rect 384406 275803 384458 275809
rect 384418 275719 384446 275803
rect 385090 275719 385118 276395
rect 384406 275713 384458 275719
rect 384406 275655 384458 275661
rect 384790 275713 384842 275719
rect 384790 275655 384842 275661
rect 385078 275713 385130 275719
rect 385078 275655 385130 275661
rect 385174 275713 385226 275719
rect 385174 275655 385226 275661
rect 384130 275488 384542 275516
rect 384514 274387 384542 275488
rect 383734 274381 383786 274387
rect 383734 274323 383786 274329
rect 383830 274381 383882 274387
rect 383830 274323 383882 274329
rect 384406 274381 384458 274387
rect 384406 274323 384458 274329
rect 384502 274381 384554 274387
rect 384502 274323 384554 274329
rect 383746 273795 383774 274323
rect 383926 274307 383978 274313
rect 383926 274249 383978 274255
rect 383638 273789 383690 273795
rect 383348 273754 383404 273763
rect 383348 273689 383404 273698
rect 383540 273754 383596 273763
rect 383638 273731 383690 273737
rect 383734 273789 383786 273795
rect 383734 273731 383786 273737
rect 383540 273689 383596 273698
rect 383252 273606 383308 273615
rect 383252 273541 383308 273550
rect 383156 273458 383212 273467
rect 383156 273393 383212 273402
rect 383170 271205 383198 273393
rect 383266 271501 383294 273541
rect 383362 272135 383390 273689
rect 383540 272570 383596 272579
rect 383540 272505 383596 272514
rect 383348 272126 383404 272135
rect 383348 272061 383404 272070
rect 383444 271978 383500 271987
rect 383444 271913 383500 271922
rect 383254 271495 383306 271501
rect 383254 271437 383306 271443
rect 383350 271495 383402 271501
rect 383350 271437 383402 271443
rect 383158 271199 383210 271205
rect 383158 271141 383210 271147
rect 383158 270903 383210 270909
rect 383158 270845 383210 270851
rect 383170 269915 383198 270845
rect 383362 270761 383390 271437
rect 383350 270755 383402 270761
rect 383350 270697 383402 270703
rect 383156 269906 383212 269915
rect 383156 269841 383212 269850
rect 382966 267943 383018 267949
rect 382966 267885 383018 267891
rect 383062 267943 383114 267949
rect 383062 267885 383114 267891
rect 383074 267727 383102 267885
rect 383062 267721 383114 267727
rect 383062 267663 383114 267669
rect 383458 265156 383486 271913
rect 383554 265452 383582 272505
rect 383650 271987 383678 273731
rect 383938 272579 383966 274249
rect 384418 273888 384446 274323
rect 384502 274233 384554 274239
rect 384502 274175 384554 274181
rect 384514 274017 384542 274175
rect 384502 274011 384554 274017
rect 384502 273953 384554 273959
rect 384598 274011 384650 274017
rect 384598 273953 384650 273959
rect 384610 273888 384638 273953
rect 384418 273860 384638 273888
rect 384802 273171 384830 275655
rect 385186 275349 385214 275655
rect 385282 275349 385310 276487
rect 385174 275343 385226 275349
rect 385174 275285 385226 275291
rect 385270 275343 385322 275349
rect 385270 275285 385322 275291
rect 385078 274455 385130 274461
rect 385078 274397 385130 274403
rect 384404 273162 384460 273171
rect 384404 273097 384460 273106
rect 384788 273162 384844 273171
rect 384788 273097 384844 273106
rect 383924 272570 383980 272579
rect 383924 272505 383980 272514
rect 383636 271978 383692 271987
rect 383636 271913 383692 271922
rect 383638 270903 383690 270909
rect 383638 270845 383690 270851
rect 383650 270761 383678 270845
rect 383924 270794 383980 270803
rect 383638 270755 383690 270761
rect 383924 270729 383980 270738
rect 383638 270697 383690 270703
rect 383938 270317 383966 270729
rect 383638 270311 383690 270317
rect 383638 270253 383690 270259
rect 383926 270311 383978 270317
rect 383926 270253 383978 270259
rect 383650 265600 383678 270253
rect 384214 267573 384266 267579
rect 384214 267515 384266 267521
rect 384226 266913 384254 267515
rect 384214 266907 384266 266913
rect 384214 266849 384266 266855
rect 383650 265572 383774 265600
rect 383554 265424 383630 265452
rect 382018 265128 382320 265156
rect 383184 265128 383486 265156
rect 383602 265142 383630 265424
rect 383746 265156 383774 265572
rect 383746 265128 384096 265156
rect 384418 265142 384446 273097
rect 384884 272126 384940 272135
rect 384884 272061 384940 272070
rect 384898 265142 384926 272061
rect 385090 265156 385118 274397
rect 385378 268023 385406 277856
rect 386230 276749 386282 276755
rect 386230 276691 386282 276697
rect 386132 272422 386188 272431
rect 386132 272357 386188 272366
rect 385556 271978 385612 271987
rect 385556 271913 385612 271922
rect 385462 271199 385514 271205
rect 385462 271141 385514 271147
rect 385366 268017 385418 268023
rect 385366 267959 385418 267965
rect 385474 266839 385502 271141
rect 385462 266833 385514 266839
rect 385462 266775 385514 266781
rect 385570 265156 385598 271913
rect 386036 270942 386092 270951
rect 385942 270903 385994 270909
rect 386036 270877 386092 270886
rect 385942 270845 385994 270851
rect 385954 270687 385982 270845
rect 386050 270687 386078 270877
rect 385942 270681 385994 270687
rect 385942 270623 385994 270629
rect 386038 270681 386090 270687
rect 386038 270623 386090 270629
rect 386146 265156 386174 272357
rect 386242 267135 386270 276691
rect 387010 276607 387038 277870
rect 387190 276675 387242 276681
rect 387190 276617 387242 276623
rect 386998 276601 387050 276607
rect 386998 276543 387050 276549
rect 387202 273647 387230 276617
rect 387190 273641 387242 273647
rect 387190 273583 387242 273589
rect 387092 272570 387148 272579
rect 387092 272505 387148 272514
rect 386612 272422 386668 272431
rect 386612 272357 386668 272366
rect 386230 267129 386282 267135
rect 386230 267071 386282 267077
rect 385090 265128 385392 265156
rect 385570 265128 385824 265156
rect 386146 265128 386208 265156
rect 386626 265142 386654 272357
rect 387106 265142 387134 272505
rect 388052 271682 388108 271691
rect 388052 271617 388108 271626
rect 387572 270794 387628 270803
rect 387572 270729 387628 270738
rect 387764 270794 387820 270803
rect 387764 270729 387766 270738
rect 387586 265142 387614 270729
rect 387818 270729 387820 270738
rect 387766 270697 387818 270703
rect 387670 268535 387722 268541
rect 387670 268477 387722 268483
rect 387766 268535 387818 268541
rect 387766 268477 387818 268483
rect 387682 265156 387710 268477
rect 387778 267357 387806 268477
rect 387766 267351 387818 267357
rect 387766 267293 387818 267299
rect 388066 265156 388094 271617
rect 388162 267949 388190 277870
rect 388724 276714 388780 276723
rect 388724 276649 388780 276658
rect 388630 273641 388682 273647
rect 388630 273583 388682 273589
rect 388642 273277 388670 273583
rect 388738 273277 388766 276649
rect 389014 273419 389066 273425
rect 389014 273361 389066 273367
rect 388630 273271 388682 273277
rect 388630 273213 388682 273219
rect 388726 273271 388778 273277
rect 388726 273213 388778 273219
rect 388726 272901 388778 272907
rect 388726 272843 388778 272849
rect 388822 272901 388874 272907
rect 388822 272843 388874 272849
rect 388738 271797 388766 272843
rect 388834 271945 388862 272843
rect 389026 272579 389054 273361
rect 389012 272570 389068 272579
rect 389012 272505 389068 272514
rect 388822 271939 388874 271945
rect 388822 271881 388874 271887
rect 388918 271939 388970 271945
rect 388918 271881 388970 271887
rect 388930 271816 388958 271881
rect 388630 271791 388682 271797
rect 388630 271733 388682 271739
rect 388726 271791 388778 271797
rect 388726 271733 388778 271739
rect 388834 271788 388958 271816
rect 389204 271830 389260 271839
rect 388642 271691 388670 271733
rect 388834 271723 388862 271788
rect 389204 271765 389260 271774
rect 388822 271717 388874 271723
rect 388628 271682 388684 271691
rect 388918 271717 388970 271723
rect 388822 271659 388874 271665
rect 388916 271682 388918 271691
rect 388970 271682 388972 271691
rect 388628 271617 388684 271626
rect 388916 271617 388972 271626
rect 388918 271051 388970 271057
rect 388918 270993 388970 270999
rect 388930 270507 388958 270993
rect 389014 270755 389066 270761
rect 389014 270697 389066 270703
rect 388724 270498 388780 270507
rect 388916 270498 388972 270507
rect 388780 270456 388862 270484
rect 388724 270433 388780 270442
rect 388438 270385 388490 270391
rect 388438 270327 388490 270333
rect 388534 270385 388586 270391
rect 388534 270327 388586 270333
rect 388450 268245 388478 270327
rect 388546 268615 388574 270327
rect 388834 268615 388862 270456
rect 388916 270433 388972 270442
rect 388534 268609 388586 268615
rect 388534 268551 388586 268557
rect 388822 268609 388874 268615
rect 388822 268551 388874 268557
rect 389026 268264 389054 270697
rect 388438 268239 388490 268245
rect 388438 268181 388490 268187
rect 388834 268236 389054 268264
rect 388246 268165 388298 268171
rect 388246 268107 388298 268113
rect 388150 267943 388202 267949
rect 388150 267885 388202 267891
rect 388258 267709 388286 268107
rect 388834 267875 388862 268236
rect 389012 268130 389068 268139
rect 388918 268091 388970 268097
rect 389012 268065 389068 268074
rect 388918 268033 388970 268039
rect 388822 267869 388874 267875
rect 388822 267811 388874 267817
rect 388930 267709 388958 268033
rect 389026 268023 389054 268065
rect 389014 268017 389066 268023
rect 389014 267959 389066 267965
rect 389110 267869 389162 267875
rect 389110 267811 389162 267817
rect 388258 267681 388958 267709
rect 388916 267538 388972 267547
rect 388972 267496 389054 267524
rect 388916 267473 388972 267482
rect 388822 267351 388874 267357
rect 388822 267293 388874 267299
rect 388834 266955 388862 267293
rect 389026 267209 389054 267496
rect 389014 267203 389066 267209
rect 389014 267145 389066 267151
rect 388820 266946 388876 266955
rect 388820 266881 388876 266890
rect 388628 266650 388684 266659
rect 388628 266585 388684 266594
rect 387682 265128 387936 265156
rect 388066 265128 388416 265156
rect 368566 265057 368618 265063
rect 368566 264999 368618 265005
rect 369142 265057 369194 265063
rect 378646 265057 378698 265063
rect 369142 264999 369194 265005
rect 369264 264989 369566 265008
rect 379510 265057 379562 265063
rect 378646 264999 378698 265005
rect 379296 265005 379510 265008
rect 379296 264999 379562 265005
rect 369264 264983 369578 264989
rect 369264 264980 369526 264983
rect 379296 264980 379550 264999
rect 382402 264980 382704 265008
rect 388642 264989 388670 266585
rect 389122 265156 389150 267811
rect 388848 265128 389150 265156
rect 389218 265142 389246 271765
rect 389314 271205 389342 277870
rect 390562 275645 390590 277870
rect 391606 277045 391658 277051
rect 391606 276987 391658 276993
rect 390550 275639 390602 275645
rect 390550 275581 390602 275587
rect 389684 273754 389740 273763
rect 389684 273689 389740 273698
rect 389698 273171 389726 273689
rect 391222 273641 391274 273647
rect 391222 273583 391274 273589
rect 391234 273499 391262 273583
rect 391222 273493 391274 273499
rect 391222 273435 391274 273441
rect 389684 273162 389740 273171
rect 389684 273097 389740 273106
rect 391618 272852 391646 276987
rect 391714 276385 391742 277870
rect 391702 276379 391754 276385
rect 391702 276321 391754 276327
rect 392854 274011 392906 274017
rect 392854 273953 392906 273959
rect 391618 272824 391838 272852
rect 391810 272759 391838 272824
rect 392470 272827 392522 272833
rect 392470 272769 392522 272775
rect 391702 272753 391754 272759
rect 391702 272695 391754 272701
rect 391798 272753 391850 272759
rect 391798 272695 391850 272701
rect 390934 272605 390986 272611
rect 389972 272570 390028 272579
rect 389878 272531 389930 272537
rect 390934 272547 390986 272553
rect 389972 272505 389974 272514
rect 389878 272473 389930 272479
rect 390026 272505 390028 272514
rect 389974 272473 390026 272479
rect 389398 271273 389450 271279
rect 389398 271215 389450 271221
rect 389302 271199 389354 271205
rect 389302 271141 389354 271147
rect 389410 268671 389438 271215
rect 389314 268643 389438 268671
rect 389314 265156 389342 268643
rect 389398 268609 389450 268615
rect 389398 268551 389450 268557
rect 389494 268609 389546 268615
rect 389494 268551 389546 268557
rect 389410 268435 389438 268551
rect 389396 268426 389452 268435
rect 389396 268361 389452 268370
rect 389506 266599 389534 268551
rect 389590 266759 389642 266765
rect 389642 266719 389822 266747
rect 389590 266701 389642 266707
rect 389794 266691 389822 266719
rect 389782 266685 389834 266691
rect 389782 266627 389834 266633
rect 389410 266571 389534 266599
rect 389410 266469 389438 266571
rect 389398 266463 389450 266469
rect 389398 266405 389450 266411
rect 389890 265156 389918 272473
rect 390550 272087 390602 272093
rect 390550 272029 390602 272035
rect 390454 271273 390506 271279
rect 390454 271215 390506 271221
rect 390466 270909 390494 271215
rect 390562 270909 390590 272029
rect 390836 271682 390892 271691
rect 390836 271617 390892 271626
rect 390646 271125 390698 271131
rect 390646 271067 390698 271073
rect 390454 270903 390506 270909
rect 390454 270845 390506 270851
rect 390550 270903 390602 270909
rect 390550 270845 390602 270851
rect 390658 268763 390686 271067
rect 390646 268757 390698 268763
rect 390646 268699 390698 268705
rect 390850 265156 390878 271617
rect 389314 265128 389712 265156
rect 389890 265128 390144 265156
rect 390624 265128 390878 265156
rect 390946 265142 390974 272547
rect 391412 271830 391468 271839
rect 391412 271765 391468 271774
rect 391028 267834 391084 267843
rect 391028 267769 391084 267778
rect 391042 266913 391070 267769
rect 391030 266907 391082 266913
rect 391030 266849 391082 266855
rect 391426 265142 391454 271765
rect 391714 265156 391742 272695
rect 391990 272383 392042 272389
rect 391990 272325 392042 272331
rect 392002 267653 392030 272325
rect 392086 270829 392138 270835
rect 392086 270771 392138 270777
rect 391990 267647 392042 267653
rect 391990 267589 392042 267595
rect 392098 265156 392126 270771
rect 392482 265156 392510 272769
rect 392866 265156 392894 273953
rect 392962 267431 392990 277870
rect 393716 276862 393772 276871
rect 393716 276797 393772 276806
rect 393730 273425 393758 276797
rect 395074 276385 395102 278573
rect 432240 278599 432458 278605
rect 432240 278596 432406 278599
rect 407542 278541 407594 278547
rect 432406 278541 432458 278547
rect 400930 278457 401232 278476
rect 400918 278451 401232 278457
rect 400970 278448 401232 278451
rect 400918 278393 400970 278399
rect 407554 278235 407582 278541
rect 474740 278490 474796 278499
rect 408130 278457 408432 278476
rect 408118 278451 408432 278457
rect 408170 278448 408432 278451
rect 474796 278448 475056 278476
rect 474740 278425 474796 278434
rect 408118 278393 408170 278399
rect 481844 278342 481900 278351
rect 460450 278309 460752 278328
rect 460438 278303 460752 278309
rect 460490 278300 460752 278303
rect 481900 278300 482160 278328
rect 481844 278277 481900 278286
rect 460438 278245 460490 278251
rect 407542 278229 407594 278235
rect 485396 278194 485452 278203
rect 407542 278171 407594 278177
rect 446338 278161 446544 278180
rect 446326 278155 446544 278161
rect 446378 278152 446544 278155
rect 485452 278152 485712 278180
rect 485396 278129 485452 278138
rect 446326 278097 446378 278103
rect 453238 278081 453290 278087
rect 488948 278046 489004 278055
rect 453290 278029 453552 278032
rect 453238 278023 453552 278029
rect 397366 278007 397418 278013
rect 453250 278004 453552 278023
rect 489004 278004 489264 278032
rect 488948 277981 489004 277990
rect 397366 277949 397418 277955
rect 395062 276379 395114 276385
rect 395062 276321 395114 276327
rect 394486 275343 394538 275349
rect 394486 275285 394538 275291
rect 394498 274387 394526 275285
rect 394390 274381 394442 274387
rect 394390 274323 394442 274329
rect 394486 274381 394538 274387
rect 394486 274323 394538 274329
rect 393622 273419 393674 273425
rect 393622 273361 393674 273367
rect 393718 273419 393770 273425
rect 393718 273361 393770 273367
rect 393142 272531 393194 272537
rect 393142 272473 393194 272479
rect 393154 269503 393182 272473
rect 393142 269497 393194 269503
rect 393142 269439 393194 269445
rect 392950 267425 393002 267431
rect 392950 267367 393002 267373
rect 393046 267129 393098 267135
rect 393046 267071 393098 267077
rect 393058 266913 393086 267071
rect 393046 266907 393098 266913
rect 393046 266849 393098 266855
rect 393046 266759 393098 266765
rect 393046 266701 393098 266707
rect 393058 266617 393086 266701
rect 393046 266611 393098 266617
rect 393046 266553 393098 266559
rect 391714 265128 391920 265156
rect 392098 265128 392352 265156
rect 392482 265128 392736 265156
rect 392866 265128 393168 265156
rect 393634 265142 393662 273361
rect 394402 272981 394430 274323
rect 394486 273715 394538 273721
rect 394486 273657 394538 273663
rect 394198 272975 394250 272981
rect 394198 272917 394250 272923
rect 394390 272975 394442 272981
rect 394390 272917 394442 272923
rect 393730 268680 394046 268708
rect 393730 268139 393758 268680
rect 393908 268574 393964 268583
rect 394018 268560 394046 268680
rect 394100 268574 394156 268583
rect 394018 268532 394100 268560
rect 393908 268509 393964 268518
rect 394100 268509 394156 268518
rect 393922 268139 393950 268509
rect 393716 268130 393772 268139
rect 393716 268065 393772 268074
rect 393908 268130 393964 268139
rect 393908 268065 393964 268074
rect 393814 267943 393866 267949
rect 393814 267885 393866 267891
rect 393910 267943 393962 267949
rect 393910 267885 393962 267891
rect 393826 265156 393854 267885
rect 393922 266321 393950 267885
rect 393910 266315 393962 266321
rect 393910 266257 393962 266263
rect 394210 265156 394238 272917
rect 394498 272907 394526 273657
rect 395362 273277 395390 277870
rect 396514 277643 396542 277870
rect 396502 277637 396554 277643
rect 396502 277579 396554 277585
rect 396118 273937 396170 273943
rect 396118 273879 396170 273885
rect 395350 273271 395402 273277
rect 395350 273213 395402 273219
rect 396022 273271 396074 273277
rect 396022 273213 396074 273219
rect 394676 273162 394732 273171
rect 394676 273097 394732 273106
rect 394486 272901 394538 272907
rect 394486 272843 394538 272849
rect 394390 271273 394442 271279
rect 394390 271215 394442 271221
rect 394486 271273 394538 271279
rect 394486 271215 394538 271221
rect 394402 270835 394430 271215
rect 394390 270829 394442 270835
rect 394390 270771 394442 270777
rect 394498 270539 394526 271215
rect 394580 270794 394636 270803
rect 394580 270729 394636 270738
rect 394594 270539 394622 270729
rect 394486 270533 394538 270539
rect 394486 270475 394538 270481
rect 394582 270533 394634 270539
rect 394582 270475 394634 270481
rect 394690 265156 394718 273097
rect 395348 273014 395404 273023
rect 395348 272949 395404 272958
rect 393826 265128 394128 265156
rect 394210 265128 394464 265156
rect 394690 265128 394944 265156
rect 395362 265142 395390 272949
rect 396034 272759 396062 273213
rect 396130 272759 396158 273879
rect 397378 273203 397406 277949
rect 415318 277933 415370 277939
rect 397078 273197 397130 273203
rect 397078 273139 397130 273145
rect 397366 273197 397418 273203
rect 397366 273139 397418 273145
rect 396022 272753 396074 272759
rect 396022 272695 396074 272701
rect 396118 272753 396170 272759
rect 396118 272695 396170 272701
rect 396214 271717 396266 271723
rect 396214 271659 396266 271665
rect 395828 270794 395884 270803
rect 395828 270729 395884 270738
rect 395842 265142 395870 270729
rect 396226 265142 396254 271659
rect 396884 267982 396940 267991
rect 396884 267917 396940 267926
rect 396598 267647 396650 267653
rect 396598 267589 396650 267595
rect 396610 267399 396638 267589
rect 396596 267390 396652 267399
rect 396596 267325 396652 267334
rect 396788 267390 396844 267399
rect 396788 267325 396790 267334
rect 396842 267325 396844 267334
rect 396790 267293 396842 267299
rect 396898 265156 396926 267917
rect 396672 265128 396926 265156
rect 397090 265156 397118 273139
rect 397366 271717 397418 271723
rect 397366 271659 397418 271665
rect 397378 268541 397406 271659
rect 397366 268535 397418 268541
rect 397366 268477 397418 268483
rect 397558 268017 397610 268023
rect 397558 267959 397610 267965
rect 397174 267647 397226 267653
rect 397174 267589 397226 267595
rect 397270 267647 397322 267653
rect 397270 267589 397322 267595
rect 397186 267399 397214 267589
rect 397172 267390 397228 267399
rect 397172 267325 397228 267334
rect 397282 267061 397310 267589
rect 397570 267376 397598 267959
rect 397762 267505 397790 277870
rect 398626 277856 398928 277884
rect 398626 274535 398654 277856
rect 398998 276897 399050 276903
rect 398998 276839 399050 276845
rect 398902 275639 398954 275645
rect 398902 275581 398954 275587
rect 398806 275343 398858 275349
rect 398806 275285 398858 275291
rect 398614 274529 398666 274535
rect 398614 274471 398666 274477
rect 398818 274387 398846 275285
rect 398806 274381 398858 274387
rect 398806 274323 398858 274329
rect 398914 273795 398942 275581
rect 398902 273789 398954 273795
rect 398902 273731 398954 273737
rect 398626 273277 398942 273296
rect 398626 273271 398954 273277
rect 398626 273268 398902 273271
rect 398626 273055 398654 273268
rect 398902 273213 398954 273219
rect 398710 273197 398762 273203
rect 398710 273139 398762 273145
rect 398614 273049 398666 273055
rect 398614 272991 398666 272997
rect 398722 272556 398750 273139
rect 399010 272981 399038 276839
rect 400066 276755 400094 277870
rect 400054 276749 400106 276755
rect 400054 276691 400106 276697
rect 400342 273863 400394 273869
rect 400342 273805 400394 273811
rect 400354 273203 400382 273805
rect 399862 273197 399914 273203
rect 399862 273139 399914 273145
rect 400342 273197 400394 273203
rect 400342 273139 400394 273145
rect 398998 272975 399050 272981
rect 398998 272917 399050 272923
rect 398722 272528 399038 272556
rect 398806 272457 398858 272463
rect 398806 272399 398858 272405
rect 398038 271199 398090 271205
rect 398038 271141 398090 271147
rect 398230 271199 398282 271205
rect 398230 271141 398282 271147
rect 397942 267573 397994 267579
rect 397942 267515 397994 267521
rect 397750 267499 397802 267505
rect 397750 267441 397802 267447
rect 397954 267376 397982 267515
rect 397570 267348 397982 267376
rect 397270 267055 397322 267061
rect 397270 266997 397322 267003
rect 397750 266833 397802 266839
rect 397750 266775 397802 266781
rect 397762 265156 397790 266775
rect 398050 265156 398078 271141
rect 398242 268171 398270 271141
rect 398818 271057 398846 272399
rect 399010 272389 399038 272528
rect 398998 272383 399050 272389
rect 398998 272325 399050 272331
rect 399874 272315 399902 273139
rect 402358 272679 402410 272685
rect 402358 272621 402410 272627
rect 401590 272383 401642 272389
rect 401590 272325 401642 272331
rect 399190 272309 399242 272315
rect 399190 272251 399242 272257
rect 399862 272309 399914 272315
rect 399862 272251 399914 272257
rect 398806 271051 398858 271057
rect 398806 270993 398858 270999
rect 398900 269758 398956 269767
rect 398900 269693 398956 269702
rect 398806 269497 398858 269503
rect 398806 269439 398858 269445
rect 398818 268911 398846 269439
rect 398806 268905 398858 268911
rect 398806 268847 398858 268853
rect 398914 268583 398942 269693
rect 398900 268574 398956 268583
rect 398900 268509 398956 268518
rect 398230 268165 398282 268171
rect 398230 268107 398282 268113
rect 398326 267129 398378 267135
rect 398326 267071 398378 267077
rect 398338 266247 398366 267071
rect 399094 266463 399146 266469
rect 399094 266405 399146 266411
rect 398326 266241 398378 266247
rect 399106 266192 399134 266405
rect 398326 266183 398378 266189
rect 398626 266164 399134 266192
rect 398626 265156 398654 266164
rect 399202 265304 399230 272251
rect 399670 272235 399722 272241
rect 399670 272177 399722 272183
rect 399382 267943 399434 267949
rect 399382 267885 399434 267891
rect 399286 267055 399338 267061
rect 399286 266997 399338 267003
rect 399298 266659 399326 266997
rect 399284 266650 399340 266659
rect 399284 266585 399340 266594
rect 399394 266321 399422 267885
rect 399574 267425 399626 267431
rect 399574 267367 399626 267373
rect 399476 266650 399532 266659
rect 399476 266585 399532 266594
rect 399382 266315 399434 266321
rect 399382 266257 399434 266263
rect 399106 265276 399230 265304
rect 399106 265156 399134 265276
rect 399490 265156 399518 266585
rect 399586 266395 399614 267367
rect 399574 266389 399626 266395
rect 399574 266331 399626 266337
rect 397090 265128 397152 265156
rect 397488 265128 397790 265156
rect 397968 265128 398078 265156
rect 398448 265128 398654 265156
rect 398880 265128 399134 265156
rect 399264 265128 399518 265156
rect 399682 265142 399710 272177
rect 400630 272161 400682 272167
rect 400630 272103 400682 272109
rect 400532 268426 400588 268435
rect 400532 268361 400588 268370
rect 400546 267991 400574 268361
rect 400532 267982 400588 267991
rect 400532 267917 400588 267926
rect 400148 266650 400204 266659
rect 400436 266650 400492 266659
rect 400148 266585 400204 266594
rect 400258 266608 400436 266636
rect 400162 265142 400190 266585
rect 400258 266469 400286 266608
rect 400436 266585 400492 266594
rect 400246 266463 400298 266469
rect 400246 266405 400298 266411
rect 400642 265142 400670 272103
rect 401302 272087 401354 272093
rect 401302 272029 401354 272035
rect 400726 268609 400778 268615
rect 400726 268551 400778 268557
rect 400738 266469 400766 268551
rect 401108 268426 401164 268435
rect 401108 268361 401164 268370
rect 401122 267875 401150 268361
rect 401110 267869 401162 267875
rect 401110 267811 401162 267817
rect 401204 266650 401260 266659
rect 401204 266585 401260 266594
rect 400726 266463 400778 266469
rect 400726 266405 400778 266411
rect 401218 265156 401246 266585
rect 400992 265128 401246 265156
rect 401314 265156 401342 272029
rect 401602 270951 401630 272325
rect 401588 270942 401644 270951
rect 401588 270877 401644 270886
rect 401314 265128 401472 265156
rect 402370 265142 402398 272621
rect 402466 270835 402494 277870
rect 403618 277495 403646 277870
rect 404482 277856 404784 277884
rect 403606 277489 403658 277495
rect 403606 277431 403658 277437
rect 403222 276823 403274 276829
rect 403222 276765 403274 276771
rect 403234 273425 403262 276765
rect 402550 273419 402602 273425
rect 402550 273361 402602 273367
rect 403222 273419 403274 273425
rect 403222 273361 403274 273367
rect 402562 270835 402590 273361
rect 404086 273345 404138 273351
rect 404086 273287 404138 273293
rect 403318 273123 403370 273129
rect 403318 273065 403370 273071
rect 402454 270829 402506 270835
rect 402454 270771 402506 270777
rect 402550 270829 402602 270835
rect 402550 270771 402602 270777
rect 403126 270533 403178 270539
rect 403126 270475 403178 270481
rect 403138 269915 403166 270475
rect 403124 269906 403180 269915
rect 403124 269841 403180 269850
rect 403222 266833 403274 266839
rect 403222 266775 403274 266781
rect 403234 266659 403262 266775
rect 402452 266650 402508 266659
rect 402452 266585 402508 266594
rect 403220 266650 403276 266659
rect 403220 266585 403276 266594
rect 402466 265156 402494 266585
rect 403330 265156 403358 273065
rect 403892 266650 403948 266659
rect 403892 266585 403948 266594
rect 403906 265156 403934 266585
rect 402466 265128 402768 265156
rect 403200 265128 403358 265156
rect 403680 265128 403934 265156
rect 404098 265142 404126 273287
rect 404482 266913 404510 277856
rect 406018 274609 406046 277870
rect 406006 274603 406058 274609
rect 406006 274545 406058 274551
rect 404950 272605 405002 272611
rect 404950 272547 405002 272553
rect 405046 272605 405098 272611
rect 405046 272547 405098 272553
rect 404470 266907 404522 266913
rect 404470 266849 404522 266855
rect 404756 266650 404812 266659
rect 404756 266585 404812 266594
rect 404770 265156 404798 266585
rect 404496 265128 404798 265156
rect 404962 265142 404990 272547
rect 405058 271723 405086 272547
rect 406006 272309 406058 272315
rect 406006 272251 406058 272257
rect 405526 272013 405578 272019
rect 405526 271955 405578 271961
rect 405046 271717 405098 271723
rect 405046 271659 405098 271665
rect 405236 266650 405292 266659
rect 405236 266585 405292 266594
rect 405250 265156 405278 266585
rect 405538 265156 405566 271955
rect 406018 267505 406046 272251
rect 406102 272161 406154 272167
rect 406102 272103 406154 272109
rect 406114 269767 406142 272103
rect 406774 272087 406826 272093
rect 406774 272029 406826 272035
rect 406786 270909 406814 272029
rect 406678 270903 406730 270909
rect 406678 270845 406730 270851
rect 406774 270903 406826 270909
rect 406774 270845 406826 270851
rect 406100 269758 406156 269767
rect 406100 269693 406156 269702
rect 406006 267499 406058 267505
rect 406006 267441 406058 267447
rect 406102 266907 406154 266913
rect 406102 266849 406154 266855
rect 406114 266469 406142 266849
rect 406196 266650 406252 266659
rect 406196 266585 406252 266594
rect 406580 266650 406636 266659
rect 406580 266585 406636 266594
rect 406102 266463 406154 266469
rect 406102 266405 406154 266411
rect 406210 265156 406238 266585
rect 406594 266469 406622 266585
rect 406582 266463 406634 266469
rect 406582 266405 406634 266411
rect 405250 265128 405408 265156
rect 405538 265128 405792 265156
rect 406210 265128 406272 265156
rect 406690 265142 406718 270845
rect 407170 266913 407198 277870
rect 409172 274642 409228 274651
rect 409172 274577 409228 274586
rect 409186 273763 409214 274577
rect 409172 273754 409228 273763
rect 409172 273689 409228 273698
rect 407638 272975 407690 272981
rect 407638 272917 407690 272923
rect 407734 272975 407786 272981
rect 407734 272917 407786 272923
rect 407650 272833 407678 272917
rect 407542 272827 407594 272833
rect 407542 272769 407594 272775
rect 407638 272827 407690 272833
rect 407638 272769 407690 272775
rect 407158 266907 407210 266913
rect 407158 266849 407210 266855
rect 407350 266759 407402 266765
rect 407350 266701 407402 266707
rect 407362 266659 407390 266701
rect 406868 266650 406924 266659
rect 406868 266585 406870 266594
rect 406922 266585 406924 266594
rect 407156 266650 407212 266659
rect 407156 266585 407212 266594
rect 407348 266650 407404 266659
rect 407348 266585 407404 266594
rect 406870 266553 406922 266559
rect 407170 265142 407198 266585
rect 407554 265142 407582 272769
rect 407746 272241 407774 272917
rect 407734 272235 407786 272241
rect 407734 272177 407786 272183
rect 409078 272087 409130 272093
rect 409078 272029 409130 272035
rect 408214 271939 408266 271945
rect 408214 271881 408266 271887
rect 407734 266611 407786 266617
rect 407734 266553 407786 266559
rect 407746 265156 407774 266553
rect 408226 265156 408254 271881
rect 408596 267834 408652 267843
rect 408596 267769 408652 267778
rect 408788 267834 408844 267843
rect 408788 267769 408844 267778
rect 408500 266946 408556 266955
rect 408500 266881 408502 266890
rect 408554 266881 408556 266890
rect 408502 266849 408554 266855
rect 408610 266839 408638 267769
rect 408802 267579 408830 267769
rect 408790 267573 408842 267579
rect 408692 267538 408748 267547
rect 408790 267515 408842 267521
rect 408884 267538 408940 267547
rect 408692 267473 408748 267482
rect 408884 267473 408940 267482
rect 408598 266833 408650 266839
rect 408598 266775 408650 266781
rect 408706 266765 408734 267473
rect 408898 267061 408926 267473
rect 408982 267425 409034 267431
rect 408982 267367 409034 267373
rect 408886 267055 408938 267061
rect 408886 266997 408938 267003
rect 408994 266987 409022 267367
rect 409090 267283 409118 272029
rect 409270 271643 409322 271649
rect 409270 271585 409322 271591
rect 409078 267277 409130 267283
rect 409078 267219 409130 267225
rect 408982 266981 409034 266987
rect 408788 266946 408844 266955
rect 408982 266923 409034 266929
rect 408788 266881 408844 266890
rect 408694 266759 408746 266765
rect 408694 266701 408746 266707
rect 408802 266659 408830 266881
rect 408788 266650 408844 266659
rect 408788 266585 408844 266594
rect 409076 266650 409132 266659
rect 409076 266585 409078 266594
rect 409130 266585 409132 266594
rect 409078 266553 409130 266559
rect 408598 266463 408650 266469
rect 408598 266405 408650 266411
rect 408610 265156 408638 266405
rect 407746 265128 408000 265156
rect 408226 265128 408480 265156
rect 408610 265128 408912 265156
rect 409282 265142 409310 271585
rect 409570 271131 409598 277870
rect 410818 277421 410846 277870
rect 411874 277856 411984 277884
rect 569878 277933 569930 277939
rect 496148 277898 496204 277907
rect 415370 277881 415632 277884
rect 415318 277875 415632 277881
rect 410806 277415 410858 277421
rect 410806 277357 410858 277363
rect 411286 272013 411338 272019
rect 411286 271955 411338 271961
rect 409942 271569 409994 271575
rect 409942 271511 409994 271517
rect 409558 271125 409610 271131
rect 409558 271067 409610 271073
rect 409654 266759 409706 266765
rect 409654 266701 409706 266707
rect 409666 266659 409694 266701
rect 409460 266650 409516 266659
rect 409460 266585 409516 266594
rect 409652 266650 409708 266659
rect 409652 266585 409708 266594
rect 409474 265156 409502 266585
rect 409954 265156 409982 271511
rect 410998 271347 411050 271353
rect 410998 271289 411050 271295
rect 410422 271125 410474 271131
rect 410422 271067 410474 271073
rect 410434 268837 410462 271067
rect 410422 268831 410474 268837
rect 410422 268773 410474 268779
rect 410326 266611 410378 266617
rect 410326 266553 410378 266559
rect 410338 265156 410366 266553
rect 409474 265128 409776 265156
rect 409954 265128 410208 265156
rect 410338 265128 410688 265156
rect 411010 265142 411038 271289
rect 411298 268245 411326 271955
rect 411478 270755 411530 270761
rect 411478 270697 411530 270703
rect 411286 268239 411338 268245
rect 411286 268181 411338 268187
rect 411490 265142 411518 270697
rect 411874 267653 411902 277856
rect 413218 274683 413246 277870
rect 413206 274677 413258 274683
rect 413206 274619 413258 274625
rect 411958 271421 412010 271427
rect 411958 271363 412010 271369
rect 411862 267647 411914 267653
rect 411862 267589 411914 267595
rect 411970 265142 411998 271363
rect 413782 267351 413834 267357
rect 413782 267293 413834 267299
rect 412534 267203 412586 267209
rect 412534 267145 412586 267151
rect 412546 265031 412574 267145
rect 413398 266981 413450 266987
rect 413398 266923 413450 266929
rect 413206 266389 413258 266395
rect 413206 266331 413258 266337
rect 413218 265771 413246 266331
rect 413410 265919 413438 266923
rect 413686 266833 413738 266839
rect 413686 266775 413738 266781
rect 413698 266215 413726 266775
rect 413794 266363 413822 267293
rect 413780 266354 413836 266363
rect 413780 266289 413836 266298
rect 414370 266247 414398 277870
rect 415330 277856 415632 277875
rect 416674 271131 416702 277870
rect 417922 277273 417950 277870
rect 417910 277267 417962 277273
rect 417910 277209 417962 277215
rect 418966 272679 419018 272685
rect 418966 272621 419018 272627
rect 418978 272315 419006 272621
rect 418966 272309 419018 272315
rect 418966 272251 419018 272257
rect 416662 271125 416714 271131
rect 416662 271067 416714 271073
rect 414838 270755 414890 270761
rect 414838 270697 414890 270703
rect 414740 269906 414796 269915
rect 414740 269841 414796 269850
rect 414754 269744 414782 269841
rect 414850 269744 414878 270697
rect 414754 269716 414878 269744
rect 417718 269571 417770 269577
rect 417718 269513 417770 269519
rect 417730 268911 417758 269513
rect 417718 268905 417770 268911
rect 417718 268847 417770 268853
rect 419074 268319 419102 277870
rect 420226 274757 420254 277870
rect 420214 274751 420266 274757
rect 420214 274693 420266 274699
rect 419062 268313 419114 268319
rect 419062 268255 419114 268261
rect 421474 267135 421502 277870
rect 422626 274091 422654 277870
rect 422614 274085 422666 274091
rect 422614 274027 422666 274033
rect 423874 268985 423902 277870
rect 425026 277125 425054 277870
rect 425014 277119 425066 277125
rect 425014 277061 425066 277067
rect 423862 268979 423914 268985
rect 423862 268921 423914 268927
rect 426274 267431 426302 277870
rect 427426 274905 427454 277870
rect 427414 274899 427466 274905
rect 427414 274841 427466 274847
rect 427606 270533 427658 270539
rect 427606 270475 427658 270481
rect 427618 270095 427646 270475
rect 427606 270089 427658 270095
rect 427606 270031 427658 270037
rect 427606 269941 427658 269947
rect 427604 269906 427606 269915
rect 427658 269906 427660 269915
rect 427604 269841 427660 269850
rect 426262 267425 426314 267431
rect 426262 267367 426314 267373
rect 421462 267129 421514 267135
rect 421462 267071 421514 267077
rect 419156 266946 419212 266955
rect 419156 266881 419212 266890
rect 419348 266946 419404 266955
rect 419348 266881 419404 266890
rect 419170 266659 419198 266881
rect 419156 266650 419212 266659
rect 419156 266585 419212 266594
rect 419362 266363 419390 266881
rect 419348 266354 419404 266363
rect 419348 266289 419404 266298
rect 414358 266241 414410 266247
rect 413684 266206 413740 266215
rect 414358 266183 414410 266189
rect 413684 266141 413740 266150
rect 428674 266099 428702 277870
rect 429538 277865 429840 277884
rect 429526 277859 429840 277865
rect 429578 277856 429840 277859
rect 429526 277801 429578 277807
rect 429140 276122 429196 276131
rect 429140 276057 429196 276066
rect 429044 274642 429100 274651
rect 429044 274577 429100 274586
rect 428948 273754 429004 273763
rect 429058 273740 429086 274577
rect 429154 273763 429182 276057
rect 429238 274677 429290 274683
rect 429236 274642 429238 274651
rect 429290 274642 429292 274651
rect 429236 274577 429292 274586
rect 429004 273712 429086 273740
rect 429140 273754 429196 273763
rect 428948 273689 429004 273698
rect 429140 273689 429196 273698
rect 429140 270498 429196 270507
rect 429140 270433 429196 270442
rect 429154 268435 429182 270433
rect 431074 269059 431102 277870
rect 431062 269053 431114 269059
rect 431062 268995 431114 269001
rect 429140 268426 429196 268435
rect 429140 268361 429196 268370
rect 433378 266691 433406 277870
rect 434530 274979 434558 277870
rect 434518 274973 434570 274979
rect 434518 274915 434570 274921
rect 434806 270755 434858 270761
rect 434806 270697 434858 270703
rect 434818 269767 434846 270697
rect 434804 269758 434860 269767
rect 434804 269693 434860 269702
rect 433366 266685 433418 266691
rect 433366 266627 433418 266633
rect 428662 266093 428714 266099
rect 428662 266035 428714 266041
rect 435682 266025 435710 277870
rect 436930 268393 436958 277870
rect 437686 270533 437738 270539
rect 437686 270475 437738 270481
rect 437698 270095 437726 270475
rect 437686 270089 437738 270095
rect 437686 270031 437738 270037
rect 437590 269941 437642 269947
rect 437588 269906 437590 269915
rect 437642 269906 437644 269915
rect 437110 269867 437162 269873
rect 437110 269809 437162 269815
rect 437494 269867 437546 269873
rect 438082 269892 438110 277870
rect 439330 277199 439358 277870
rect 439318 277193 439370 277199
rect 439318 277135 439370 277141
rect 440482 274165 440510 277870
rect 441730 276311 441758 277870
rect 441718 276305 441770 276311
rect 441718 276247 441770 276253
rect 440470 274159 440522 274165
rect 440470 274101 440522 274107
rect 438082 269864 438398 269892
rect 437588 269841 437644 269850
rect 437494 269809 437546 269815
rect 437122 269744 437150 269809
rect 437506 269744 437534 269809
rect 437122 269716 437534 269744
rect 437986 269725 438206 269744
rect 437974 269719 438218 269725
rect 438026 269716 438166 269719
rect 437974 269661 438026 269667
rect 438166 269661 438218 269667
rect 437398 269645 437450 269651
rect 437590 269645 437642 269651
rect 437450 269605 437590 269633
rect 437398 269587 437450 269593
rect 437590 269587 437642 269593
rect 437782 269645 437834 269651
rect 437878 269645 437930 269651
rect 437834 269593 437878 269596
rect 437782 269587 437930 269593
rect 437686 269571 437738 269577
rect 437794 269568 437918 269587
rect 437686 269513 437738 269519
rect 437494 269497 437546 269503
rect 437590 269497 437642 269503
rect 437546 269445 437590 269448
rect 437494 269439 437642 269445
rect 437302 269423 437354 269429
rect 437398 269423 437450 269429
rect 437354 269383 437398 269411
rect 437302 269365 437354 269371
rect 437506 269420 437630 269439
rect 437398 269365 437450 269371
rect 437698 268911 437726 269513
rect 437794 269429 437918 269448
rect 437782 269423 437918 269429
rect 437834 269420 437918 269423
rect 437782 269365 437834 269371
rect 437890 269300 437918 269420
rect 438262 269423 438314 269429
rect 438262 269365 438314 269371
rect 438274 269300 438302 269365
rect 437890 269272 438302 269300
rect 438370 269207 438398 269864
rect 438358 269201 438410 269207
rect 438358 269143 438410 269149
rect 437686 268905 437738 268911
rect 437686 268847 437738 268853
rect 436918 268387 436970 268393
rect 436918 268329 436970 268335
rect 439124 266798 439180 266807
rect 439124 266733 439180 266742
rect 439028 266354 439084 266363
rect 439028 266289 439084 266298
rect 435670 266019 435722 266025
rect 435670 265961 435722 265967
rect 413396 265910 413452 265919
rect 413396 265845 413452 265854
rect 413204 265762 413260 265771
rect 413204 265697 413260 265706
rect 439042 265623 439070 266289
rect 439138 266067 439166 266733
rect 439220 266650 439276 266659
rect 439220 266585 439276 266594
rect 439124 266058 439180 266067
rect 439124 265993 439180 266002
rect 439234 265919 439262 266585
rect 439316 266206 439372 266215
rect 439316 266141 439372 266150
rect 439220 265910 439276 265919
rect 439220 265845 439276 265854
rect 439028 265614 439084 265623
rect 439028 265549 439084 265558
rect 439330 265475 439358 266141
rect 442882 265951 442910 277870
rect 443842 277856 444144 277884
rect 443842 277791 443870 277856
rect 443830 277785 443882 277791
rect 443830 277727 443882 277733
rect 445282 270613 445310 277870
rect 445270 270607 445322 270613
rect 445270 270549 445322 270555
rect 447682 266543 447710 277870
rect 448834 276237 448862 277870
rect 448822 276231 448874 276237
rect 448822 276173 448874 276179
rect 449204 276122 449260 276131
rect 449204 276057 449260 276066
rect 449110 274677 449162 274683
rect 449108 274642 449110 274651
rect 449162 274642 449164 274651
rect 449108 274577 449164 274586
rect 449218 273763 449246 276057
rect 449204 273754 449260 273763
rect 449204 273689 449260 273698
rect 449204 270498 449260 270507
rect 449204 270433 449260 270442
rect 449218 268435 449246 270433
rect 449204 268426 449260 268435
rect 449204 268361 449260 268370
rect 447670 266537 447722 266543
rect 447670 266479 447722 266485
rect 442870 265945 442922 265951
rect 442870 265887 442922 265893
rect 449986 265877 450014 277870
rect 451138 268467 451166 277870
rect 452386 270465 452414 277870
rect 454786 277717 454814 277870
rect 454774 277711 454826 277717
rect 454774 277653 454826 277659
rect 455938 276089 455966 277870
rect 455926 276083 455978 276089
rect 455926 276025 455978 276031
rect 452374 270459 452426 270465
rect 452374 270401 452426 270407
rect 451126 268461 451178 268467
rect 451126 268403 451178 268409
rect 449974 265871 450026 265877
rect 449974 265813 450026 265819
rect 457186 265803 457214 277870
rect 458338 274239 458366 277870
rect 458326 274233 458378 274239
rect 458326 274175 458378 274181
rect 459586 270243 459614 277870
rect 459574 270237 459626 270243
rect 459574 270179 459626 270185
rect 457940 269758 457996 269767
rect 457940 269693 457996 269702
rect 458612 269758 458668 269767
rect 458612 269693 458668 269702
rect 457954 269503 457982 269693
rect 458230 269571 458282 269577
rect 458230 269513 458282 269519
rect 457942 269497 457994 269503
rect 457942 269439 457994 269445
rect 458242 269448 458270 269513
rect 458626 269503 458654 269693
rect 458614 269497 458666 269503
rect 458242 269420 458558 269448
rect 458614 269439 458666 269445
rect 457942 269201 457994 269207
rect 457942 269143 457994 269149
rect 457954 269004 457982 269143
rect 458038 269053 458090 269059
rect 457954 269001 458038 269004
rect 457954 268995 458090 269001
rect 457954 268976 458078 268995
rect 458530 268985 458558 269420
rect 458518 268979 458570 268985
rect 458518 268921 458570 268927
rect 459284 266798 459340 266807
rect 459284 266733 459340 266742
rect 458132 266354 458188 266363
rect 458132 266289 458188 266298
rect 457174 265797 457226 265803
rect 457174 265739 457226 265745
rect 458146 265623 458174 266289
rect 459298 266067 459326 266733
rect 459380 266650 459436 266659
rect 459380 266585 459436 266594
rect 459284 266058 459340 266067
rect 459284 265993 459340 266002
rect 459394 265919 459422 266585
rect 461986 266321 462014 277870
rect 463138 275941 463166 277870
rect 463126 275935 463178 275941
rect 463126 275877 463178 275883
rect 461974 266315 462026 266321
rect 461974 266257 462026 266263
rect 459380 265910 459436 265919
rect 459380 265845 459436 265854
rect 459572 265910 459628 265919
rect 459572 265845 459628 265854
rect 458132 265614 458188 265623
rect 458132 265549 458188 265558
rect 459586 265475 459614 265845
rect 464290 265729 464318 277870
rect 465538 277569 465566 277870
rect 465526 277563 465578 277569
rect 465526 277505 465578 277511
rect 466594 270021 466622 277870
rect 467842 276575 467870 277870
rect 467828 276566 467884 276575
rect 467828 276501 467884 276510
rect 468994 272019 469022 277870
rect 469460 276122 469516 276131
rect 469460 276057 469516 276066
rect 469474 273763 469502 276057
rect 470242 275793 470270 277870
rect 470230 275787 470282 275793
rect 470230 275729 470282 275735
rect 469556 274642 469612 274651
rect 469556 274577 469612 274586
rect 469570 274239 469598 274577
rect 469558 274233 469610 274239
rect 469558 274175 469610 274181
rect 469460 273754 469516 273763
rect 469460 273689 469516 273698
rect 468982 272013 469034 272019
rect 468982 271955 469034 271961
rect 469460 270498 469516 270507
rect 469516 270456 469598 270484
rect 469460 270433 469516 270442
rect 466582 270015 466634 270021
rect 466582 269957 466634 269963
rect 469570 269915 469598 270456
rect 469364 269906 469420 269915
rect 469556 269906 469612 269915
rect 469420 269864 469502 269892
rect 469364 269841 469420 269850
rect 469474 269767 469502 269864
rect 469556 269841 469612 269850
rect 469460 269758 469516 269767
rect 469460 269693 469516 269702
rect 467926 269275 467978 269281
rect 467926 269217 467978 269223
rect 467938 269059 467966 269217
rect 467926 269053 467978 269059
rect 467926 268995 467978 269001
rect 464278 265723 464330 265729
rect 464278 265665 464330 265671
rect 471394 265655 471422 277870
rect 472642 274313 472670 277870
rect 472630 274307 472682 274313
rect 472630 274249 472682 274255
rect 473794 269947 473822 277870
rect 473782 269941 473834 269947
rect 473782 269883 473834 269889
rect 476194 266173 476222 277870
rect 477442 273911 477470 277870
rect 477622 274233 477674 274239
rect 477622 274175 477674 274181
rect 477634 273911 477662 274175
rect 477428 273902 477484 273911
rect 477428 273837 477484 273846
rect 477620 273902 477676 273911
rect 477620 273837 477676 273846
rect 478006 269571 478058 269577
rect 478006 269513 478058 269519
rect 478018 268985 478046 269513
rect 478006 268979 478058 268985
rect 478006 268921 478058 268927
rect 476182 266167 476234 266173
rect 476182 266109 476234 266115
rect 471382 265649 471434 265655
rect 471382 265591 471434 265597
rect 478594 265581 478622 277870
rect 479746 277347 479774 277870
rect 479734 277341 479786 277347
rect 479734 277283 479786 277289
rect 480994 272408 481022 277870
rect 480994 272380 481118 272408
rect 480982 272235 481034 272241
rect 480982 272177 481034 272183
rect 480994 267991 481022 272177
rect 481090 269799 481118 272380
rect 483298 271205 483326 277870
rect 484450 274059 484478 277870
rect 484436 274050 484492 274059
rect 484436 273985 484492 273994
rect 486742 272309 486794 272315
rect 486742 272251 486794 272257
rect 483286 271199 483338 271205
rect 483286 271141 483338 271147
rect 481078 269793 481130 269799
rect 483958 269793 484010 269799
rect 481078 269735 481130 269741
rect 483860 269758 483916 269767
rect 483916 269741 483958 269744
rect 483916 269735 484010 269741
rect 483916 269716 483998 269735
rect 483860 269693 483916 269702
rect 483874 269619 484190 269633
rect 483860 269610 484204 269619
rect 483916 269605 484148 269610
rect 483860 269545 483916 269554
rect 484148 269545 484204 269554
rect 483958 268905 484010 268911
rect 483958 268847 484010 268853
rect 483862 268831 483914 268837
rect 483862 268773 483914 268779
rect 483874 268708 483902 268773
rect 483970 268708 483998 268847
rect 483874 268680 483998 268708
rect 486754 268139 486782 272251
rect 486850 272093 486878 277870
rect 486838 272087 486890 272093
rect 486838 272029 486890 272035
rect 488098 269725 488126 277870
rect 489524 276122 489580 276131
rect 489524 276057 489580 276066
rect 489428 274642 489484 274651
rect 489428 274577 489484 274586
rect 489442 273911 489470 274577
rect 489428 273902 489484 273911
rect 489428 273837 489484 273846
rect 489538 273763 489566 276057
rect 489524 273754 489580 273763
rect 489524 273689 489580 273698
rect 490498 273203 490526 277870
rect 491650 274207 491678 277870
rect 491636 274198 491692 274207
rect 491636 274133 491692 274142
rect 490486 273197 490538 273203
rect 490486 273139 490538 273145
rect 489524 270498 489580 270507
rect 489524 270433 489580 270442
rect 489428 269906 489484 269915
rect 489538 269892 489566 270433
rect 489484 269864 489566 269892
rect 489428 269841 489484 269850
rect 488086 269719 488138 269725
rect 488086 269661 488138 269667
rect 486740 268130 486796 268139
rect 486740 268065 486796 268074
rect 480980 267982 481036 267991
rect 480980 267917 481036 267926
rect 479348 266798 479404 266807
rect 479348 266733 479404 266742
rect 479540 266798 479596 266807
rect 479540 266733 479596 266742
rect 479362 266067 479390 266733
rect 479444 266650 479500 266659
rect 479444 266585 479500 266594
rect 479458 266215 479486 266585
rect 479554 266363 479582 266733
rect 479636 266650 479692 266659
rect 479636 266585 479692 266594
rect 479540 266354 479596 266363
rect 479540 266289 479596 266298
rect 479444 266206 479500 266215
rect 479444 266141 479500 266150
rect 479348 266058 479404 266067
rect 479348 265993 479404 266002
rect 479650 265919 479678 266585
rect 479636 265910 479692 265919
rect 479636 265845 479692 265854
rect 478582 265575 478634 265581
rect 478582 265517 478634 265523
rect 492898 265507 492926 277870
rect 494050 273425 494078 277870
rect 494038 273419 494090 273425
rect 494038 273361 494090 273367
rect 495202 269651 495230 277870
rect 496204 277856 496464 277884
rect 496148 277833 496204 277842
rect 497602 272611 497630 277870
rect 498850 274207 498878 277870
rect 498836 274198 498892 274207
rect 498836 274133 498892 274142
rect 497590 272605 497642 272611
rect 497590 272547 497642 272553
rect 497686 272605 497738 272611
rect 497686 272547 497738 272553
rect 495190 269645 495242 269651
rect 495190 269587 495242 269593
rect 497698 265919 497726 272547
rect 497684 265910 497740 265919
rect 497684 265845 497740 265854
rect 492886 265501 492938 265507
rect 439316 265466 439372 265475
rect 459572 265466 459628 265475
rect 439316 265401 439372 265410
rect 455074 265424 455198 265452
rect 455074 265327 455102 265424
rect 413204 265318 413260 265327
rect 413204 265253 413260 265262
rect 455060 265318 455116 265327
rect 455060 265253 455116 265262
rect 412532 265022 412588 265031
rect 401602 264994 401904 265008
rect 388630 264983 388682 264989
rect 369526 264925 369578 264931
rect 382402 264915 382430 264980
rect 388630 264925 388682 264931
rect 401588 264985 401904 264994
rect 401644 264980 401904 264985
rect 413218 264989 413246 265253
rect 455170 264989 455198 265424
rect 492886 265443 492938 265449
rect 499906 265433 499934 277870
rect 501154 272685 501182 277870
rect 501238 273123 501290 273129
rect 501238 273065 501290 273071
rect 501142 272679 501194 272685
rect 501142 272621 501194 272627
rect 501058 269577 501182 269596
rect 501046 269571 501194 269577
rect 501098 269568 501142 269571
rect 501046 269513 501098 269519
rect 501142 269513 501194 269519
rect 501250 266215 501278 273065
rect 502306 268879 502334 277870
rect 503266 277856 503568 277884
rect 569878 277875 569930 277881
rect 503266 277759 503294 277856
rect 503252 277750 503308 277759
rect 503252 277685 503308 277694
rect 504404 274642 504460 274651
rect 504404 274577 504460 274586
rect 504418 274207 504446 274577
rect 504404 274198 504460 274207
rect 504404 274133 504460 274142
rect 504706 272759 504734 277870
rect 505954 274503 505982 277870
rect 505940 274494 505996 274503
rect 505940 274429 505996 274438
rect 504694 272753 504746 272759
rect 504694 272695 504746 272701
rect 505270 272679 505322 272685
rect 505270 272621 505322 272627
rect 502292 268870 502348 268879
rect 502292 268805 502348 268814
rect 505282 266511 505310 272621
rect 505268 266502 505324 266511
rect 505268 266437 505324 266446
rect 501622 266389 501674 266395
rect 501622 266331 501674 266337
rect 501236 266206 501292 266215
rect 501236 266141 501292 266150
rect 459572 265401 459628 265410
rect 499894 265427 499946 265433
rect 499894 265369 499946 265375
rect 475124 265170 475180 265179
rect 475124 265105 475180 265114
rect 483860 265170 483916 265179
rect 483860 265105 483916 265114
rect 475138 264989 475166 265105
rect 483874 264989 483902 265105
rect 412532 264957 412588 264966
rect 413206 264983 413258 264989
rect 401588 264920 401644 264929
rect 413206 264925 413258 264931
rect 455158 264983 455210 264989
rect 455158 264925 455210 264931
rect 475126 264983 475178 264989
rect 475126 264925 475178 264931
rect 483862 264983 483914 264989
rect 483862 264925 483914 264931
rect 382390 264909 382442 264915
rect 368194 264832 368352 264860
rect 382390 264851 382442 264857
rect 501634 251669 501662 266331
rect 507106 265359 507134 277870
rect 508354 276977 508382 277870
rect 508342 276971 508394 276977
rect 508342 276913 508394 276919
rect 509506 269027 509534 277870
rect 509780 276122 509836 276131
rect 509780 276057 509836 276066
rect 509794 274503 509822 276057
rect 509780 274494 509836 274503
rect 509780 274429 509836 274438
rect 509780 270498 509836 270507
rect 509780 270433 509836 270442
rect 509794 269027 509822 270433
rect 509878 269645 509930 269651
rect 509878 269587 509930 269593
rect 509890 269207 509918 269587
rect 509878 269201 509930 269207
rect 509878 269143 509930 269149
rect 509492 269018 509548 269027
rect 509492 268953 509548 268962
rect 509780 269018 509836 269027
rect 509780 268953 509836 268962
rect 507094 265353 507146 265359
rect 507094 265295 507146 265301
rect 510658 265285 510686 277870
rect 511906 271279 511934 277870
rect 511894 271273 511946 271279
rect 511894 271215 511946 271221
rect 513058 269175 513086 277870
rect 513044 269166 513100 269175
rect 513044 269101 513100 269110
rect 510646 265279 510698 265285
rect 510646 265221 510698 265227
rect 514306 265211 514334 277870
rect 515458 267727 515486 277870
rect 516610 271057 516638 277870
rect 517762 277611 517790 277870
rect 517748 277602 517804 277611
rect 517748 277537 517804 277546
rect 519010 272907 519038 277870
rect 518998 272901 519050 272907
rect 518998 272843 519050 272849
rect 516598 271051 516650 271057
rect 516598 270993 516650 270999
rect 518326 269793 518378 269799
rect 518324 269758 518326 269767
rect 518378 269758 518380 269767
rect 518324 269693 518380 269702
rect 520162 269281 520190 277870
rect 520150 269275 520202 269281
rect 520150 269217 520202 269223
rect 515446 267721 515498 267727
rect 515446 267663 515498 267669
rect 514294 265205 514346 265211
rect 511124 265170 511180 265179
rect 514294 265147 514346 265153
rect 511124 265105 511180 265114
rect 511138 264989 511166 265105
rect 521410 265031 521438 277870
rect 522562 272833 522590 277870
rect 522550 272827 522602 272833
rect 522550 272769 522602 272775
rect 523810 270359 523838 277870
rect 524962 277463 524990 277870
rect 524948 277454 525004 277463
rect 524948 277389 525004 277398
rect 526114 272537 526142 277870
rect 526102 272531 526154 272537
rect 526102 272473 526154 272479
rect 527362 270983 527390 277870
rect 527350 270977 527402 270983
rect 527350 270919 527402 270925
rect 524372 270498 524428 270507
rect 524372 270433 524428 270442
rect 523796 270350 523852 270359
rect 523796 270285 523852 270294
rect 524386 269027 524414 270433
rect 524372 269018 524428 269027
rect 524372 268953 524428 268962
rect 528514 267843 528542 277870
rect 529762 272463 529790 277870
rect 529844 276122 529900 276131
rect 529844 276057 529900 276066
rect 529858 274503 529886 276057
rect 529844 274494 529900 274503
rect 529844 274429 529900 274438
rect 529750 272457 529802 272463
rect 529750 272399 529802 272405
rect 529940 269906 529996 269915
rect 529940 269841 529996 269850
rect 529844 269758 529900 269767
rect 529954 269744 529982 269841
rect 529900 269716 529982 269744
rect 529844 269693 529900 269702
rect 529846 269571 529898 269577
rect 529846 269513 529898 269519
rect 529858 269207 529886 269513
rect 529846 269201 529898 269207
rect 529846 269143 529898 269149
rect 528500 267834 528556 267843
rect 528500 267769 528556 267778
rect 530914 267695 530942 277870
rect 532162 277315 532190 277870
rect 532148 277306 532204 277315
rect 532148 277241 532204 277250
rect 533218 272981 533246 277870
rect 533206 272975 533258 272981
rect 533206 272917 533258 272923
rect 532822 269497 532874 269503
rect 532822 269439 532874 269445
rect 533110 269497 533162 269503
rect 533110 269439 533162 269445
rect 532834 269300 532862 269439
rect 533122 269300 533150 269439
rect 532834 269272 533150 269300
rect 530900 267686 530956 267695
rect 530900 267621 530956 267630
rect 534466 267399 534494 277870
rect 535618 277167 535646 277870
rect 535604 277158 535660 277167
rect 535604 277093 535660 277102
rect 536866 270835 536894 277870
rect 536854 270829 536906 270835
rect 536854 270771 536906 270777
rect 538018 267547 538046 277870
rect 539266 269873 539294 277870
rect 540418 273055 540446 277870
rect 540406 273049 540458 273055
rect 540406 272991 540458 272997
rect 539254 269867 539306 269873
rect 539254 269809 539306 269815
rect 538004 267538 538060 267547
rect 538004 267473 538060 267482
rect 534452 267390 534508 267399
rect 534452 267325 534508 267334
rect 541570 267251 541598 277870
rect 541556 267242 541612 267251
rect 541556 267177 541612 267186
rect 542818 266955 542846 277870
rect 543970 270909 543998 277870
rect 543958 270903 544010 270909
rect 543958 270845 544010 270851
rect 545218 267103 545246 277870
rect 546370 277019 546398 277870
rect 546356 277010 546412 277019
rect 546356 276945 546412 276954
rect 545684 276122 545740 276131
rect 545684 276057 545740 276066
rect 545698 274503 545726 276057
rect 545684 274494 545740 274503
rect 545684 274429 545740 274438
rect 547618 272389 547646 277870
rect 547606 272383 547658 272389
rect 547606 272325 547658 272331
rect 548770 271099 548798 277870
rect 549922 271871 549950 277870
rect 549910 271865 549962 271871
rect 549910 271807 549962 271813
rect 548756 271090 548812 271099
rect 548756 271025 548812 271034
rect 545204 267094 545260 267103
rect 545204 267029 545260 267038
rect 542804 266946 542860 266955
rect 542804 266881 542860 266890
rect 521396 265022 521452 265031
rect 511126 264983 511178 264989
rect 521396 264957 521452 264966
rect 511126 264925 511178 264931
rect 551074 264915 551102 277870
rect 552322 271247 552350 277870
rect 552982 274233 553034 274239
rect 552980 274198 552982 274207
rect 553034 274198 553036 274207
rect 552980 274133 553036 274142
rect 553474 273573 553502 277870
rect 554722 274831 554750 277870
rect 554710 274825 554762 274831
rect 554710 274767 554762 274773
rect 553462 273567 553514 273573
rect 553462 273509 553514 273515
rect 555874 271395 555902 277870
rect 557026 275571 557054 277870
rect 557014 275565 557066 275571
rect 557014 275507 557066 275513
rect 555860 271386 555916 271395
rect 555860 271321 555916 271330
rect 552308 271238 552364 271247
rect 552308 271173 552364 271182
rect 552980 270498 553036 270507
rect 552980 270433 552982 270442
rect 553034 270433 553036 270442
rect 552982 270401 553034 270407
rect 552980 269906 553036 269915
rect 552980 269841 553036 269850
rect 552994 269744 553022 269841
rect 553076 269758 553132 269767
rect 552994 269716 553076 269744
rect 553076 269693 553132 269702
rect 558274 269133 558302 277870
rect 559426 271543 559454 277870
rect 560086 272383 560138 272389
rect 560086 272325 560138 272331
rect 559412 271534 559468 271543
rect 559412 271469 559468 271478
rect 558262 269127 558314 269133
rect 558262 269069 558314 269075
rect 560098 268837 560126 272325
rect 560674 269577 560702 277870
rect 561826 276459 561854 277870
rect 561814 276453 561866 276459
rect 561814 276395 561866 276401
rect 563074 272727 563102 277870
rect 564226 275497 564254 277870
rect 564214 275491 564266 275497
rect 564214 275433 564266 275439
rect 563060 272718 563116 272727
rect 563060 272653 563116 272662
rect 565474 270687 565502 277870
rect 566530 272875 566558 277870
rect 566516 272866 566572 272875
rect 566516 272801 566572 272810
rect 565462 270681 565514 270687
rect 565462 270623 565514 270629
rect 560662 269571 560714 269577
rect 560662 269513 560714 269519
rect 567778 269429 567806 277870
rect 568930 276385 568958 277870
rect 568918 276379 568970 276385
rect 568918 276321 568970 276327
rect 567766 269423 567818 269429
rect 567766 269365 567818 269371
rect 560086 268831 560138 268837
rect 560086 268773 560138 268779
rect 569890 266395 569918 277875
rect 570068 276122 570124 276131
rect 570068 276057 570124 276066
rect 570082 274503 570110 276057
rect 570068 274494 570124 274503
rect 570068 274429 570124 274438
rect 570178 269619 570206 277870
rect 571330 275423 571358 277870
rect 571318 275417 571370 275423
rect 571318 275359 571370 275365
rect 570164 269610 570220 269619
rect 570164 269545 570220 269554
rect 572482 268097 572510 277870
rect 573044 274346 573100 274355
rect 573044 274281 573100 274290
rect 573058 274239 573086 274281
rect 573046 274233 573098 274239
rect 573046 274175 573098 274181
rect 573730 272283 573758 277870
rect 573716 272274 573772 272283
rect 573716 272209 573772 272218
rect 573046 270459 573098 270465
rect 573046 270401 573098 270407
rect 573058 270359 573086 270401
rect 573044 270350 573100 270359
rect 573044 270285 573100 270294
rect 573140 270202 573196 270211
rect 573140 270137 573196 270146
rect 573154 270021 573182 270137
rect 573142 270015 573194 270021
rect 573142 269957 573194 269963
rect 573140 269610 573196 269619
rect 573140 269545 573142 269554
rect 573194 269545 573196 269554
rect 573142 269513 573194 269519
rect 574882 269355 574910 277870
rect 576130 276163 576158 277870
rect 576118 276157 576170 276163
rect 576118 276099 576170 276105
rect 574870 269349 574922 269355
rect 574870 269291 574922 269297
rect 577282 268731 577310 277870
rect 578530 275275 578558 277870
rect 578518 275269 578570 275275
rect 578518 275211 578570 275217
rect 579682 270391 579710 277870
rect 579670 270385 579722 270391
rect 579670 270327 579722 270333
rect 580930 269323 580958 277870
rect 582082 270655 582110 277870
rect 583234 276015 583262 277870
rect 583222 276009 583274 276015
rect 583222 275951 583274 275957
rect 584386 273319 584414 277870
rect 585634 275201 585662 277870
rect 585622 275195 585674 275201
rect 585622 275137 585674 275143
rect 584756 274494 584812 274503
rect 584756 274429 584812 274438
rect 584564 274346 584620 274355
rect 584770 274332 584798 274429
rect 584620 274304 584798 274332
rect 584564 274281 584620 274290
rect 584372 273310 584428 273319
rect 584372 273245 584428 273254
rect 582068 270646 582124 270655
rect 582068 270581 582124 270590
rect 586786 270317 586814 277870
rect 587938 276131 587966 277870
rect 587924 276122 587980 276131
rect 587924 276057 587980 276066
rect 586774 270311 586826 270317
rect 586774 270253 586826 270259
rect 589186 270021 589214 277870
rect 590338 275867 590366 277870
rect 591586 275983 591614 277870
rect 591572 275974 591628 275983
rect 591572 275909 591628 275918
rect 590326 275861 590378 275867
rect 590326 275803 590378 275809
rect 592738 275127 592766 277870
rect 592726 275121 592778 275127
rect 592726 275063 592778 275069
rect 593300 274494 593356 274503
rect 593300 274429 593302 274438
rect 593354 274429 593356 274438
rect 593302 274397 593354 274403
rect 590420 270498 590476 270507
rect 590420 270433 590422 270442
rect 590474 270433 590476 270442
rect 590422 270401 590474 270407
rect 593986 270169 594014 277870
rect 595138 275835 595166 277870
rect 595124 275826 595180 275835
rect 595124 275761 595180 275770
rect 593974 270163 594026 270169
rect 593974 270105 594026 270111
rect 596386 270063 596414 277870
rect 597538 270095 597566 277870
rect 598786 275687 598814 277870
rect 598772 275678 598828 275687
rect 598772 275613 598828 275622
rect 599842 275053 599870 277870
rect 599830 275047 599882 275053
rect 599830 274989 599882 274995
rect 601090 271501 601118 277870
rect 602242 275539 602270 277870
rect 603394 276427 603422 277870
rect 603380 276418 603436 276427
rect 603380 276353 603436 276362
rect 604642 275719 604670 277870
rect 604630 275713 604682 275719
rect 604630 275655 604682 275661
rect 602228 275530 602284 275539
rect 602228 275465 602284 275474
rect 605794 273467 605822 277870
rect 605780 273458 605836 273467
rect 605780 273393 605836 273402
rect 601078 271495 601130 271501
rect 601078 271437 601130 271443
rect 600500 270498 600556 270507
rect 600500 270433 600502 270442
rect 600554 270433 600556 270442
rect 600502 270401 600554 270407
rect 597526 270089 597578 270095
rect 596372 270054 596428 270063
rect 589174 270015 589226 270021
rect 597526 270031 597578 270037
rect 596372 269989 596428 269998
rect 589174 269957 589226 269963
rect 593204 269758 593260 269767
rect 593204 269693 593260 269702
rect 593218 269577 593246 269693
rect 593206 269571 593258 269577
rect 593206 269513 593258 269519
rect 580916 269314 580972 269323
rect 580916 269249 580972 269258
rect 577268 268722 577324 268731
rect 577268 268657 577324 268666
rect 572470 268091 572522 268097
rect 572470 268033 572522 268039
rect 569878 266389 569930 266395
rect 569878 266331 569930 266337
rect 607042 265179 607070 277870
rect 608194 271797 608222 277870
rect 609442 272167 609470 277870
rect 609430 272161 609482 272167
rect 609430 272103 609482 272109
rect 608182 271791 608234 271797
rect 608182 271733 608234 271739
rect 610594 269767 610622 277870
rect 610580 269758 610636 269767
rect 610580 269693 610636 269702
rect 607028 265170 607084 265179
rect 611842 265137 611870 277870
rect 612994 275391 613022 277870
rect 612980 275382 613036 275391
rect 612980 275317 613036 275326
rect 613364 274494 613420 274503
rect 613364 274429 613366 274438
rect 613418 274429 613420 274438
rect 613366 274397 613418 274403
rect 614242 272611 614270 277870
rect 615394 276681 615422 277870
rect 615382 276675 615434 276681
rect 615382 276617 615434 276623
rect 616546 275243 616574 277870
rect 616532 275234 616588 275243
rect 616532 275169 616588 275178
rect 617698 273129 617726 277870
rect 618850 275645 618878 277870
rect 618838 275639 618890 275645
rect 618838 275581 618890 275587
rect 619126 274603 619178 274609
rect 619126 274545 619178 274551
rect 619138 274355 619166 274545
rect 619124 274346 619180 274355
rect 619124 274281 619180 274290
rect 617686 273123 617738 273129
rect 617686 273065 617738 273071
rect 614230 272605 614282 272611
rect 614230 272547 614282 272553
rect 620098 268583 620126 277870
rect 620564 275234 620620 275243
rect 620564 275169 620620 275178
rect 620578 274799 620606 275169
rect 620564 274790 620620 274799
rect 620564 274725 620620 274734
rect 621250 272685 621278 277870
rect 622498 273499 622526 277870
rect 623650 275095 623678 277870
rect 624898 276279 624926 277870
rect 624884 276270 624940 276279
rect 624884 276205 624940 276214
rect 623636 275086 623692 275095
rect 623636 275021 623692 275030
rect 622486 273493 622538 273499
rect 622486 273435 622538 273441
rect 621238 272679 621290 272685
rect 621238 272621 621290 272627
rect 626050 269503 626078 277870
rect 627298 274609 627326 277870
rect 627286 274603 627338 274609
rect 627286 274545 627338 274551
rect 626038 269497 626090 269503
rect 626038 269439 626090 269445
rect 620084 268574 620140 268583
rect 620084 268509 620140 268518
rect 628450 267801 628478 277870
rect 629698 273277 629726 277870
rect 629686 273271 629738 273277
rect 629686 273213 629738 273219
rect 630850 268287 630878 277870
rect 632098 269471 632126 277870
rect 632084 269462 632140 269471
rect 632084 269397 632140 269406
rect 632086 269275 632138 269281
rect 632086 269217 632138 269223
rect 630836 268278 630892 268287
rect 630836 268213 630892 268222
rect 628438 267795 628490 267801
rect 628438 267737 628490 267743
rect 607028 265105 607084 265114
rect 611830 265131 611882 265137
rect 611830 265073 611882 265079
rect 551062 264909 551114 264915
rect 551062 264851 551114 264857
rect 632098 253519 632126 269217
rect 633154 265063 633182 277870
rect 634306 272241 634334 277870
rect 634294 272235 634346 272241
rect 634294 272177 634346 272183
rect 635554 265771 635582 277870
rect 636706 275349 636734 277870
rect 636694 275343 636746 275349
rect 636694 275285 636746 275291
rect 637954 275243 637982 277870
rect 639106 276533 639134 277870
rect 640354 276607 640382 277870
rect 640342 276601 640394 276607
rect 640342 276543 640394 276549
rect 639094 276527 639146 276533
rect 639094 276469 639146 276475
rect 637940 275234 637996 275243
rect 637940 275169 637996 275178
rect 641506 272315 641534 277870
rect 641494 272309 641546 272315
rect 641494 272251 641546 272257
rect 642754 266807 642782 277870
rect 643906 272389 643934 277870
rect 645154 274947 645182 277870
rect 645140 274938 645196 274947
rect 645140 274873 645196 274882
rect 643894 272383 643946 272389
rect 643894 272325 643946 272331
rect 642740 266798 642796 266807
rect 642740 266733 642796 266742
rect 646306 266659 646334 277870
rect 647554 270803 647582 277870
rect 648706 273615 648734 277870
rect 648692 273606 648748 273615
rect 648692 273541 648748 273550
rect 647540 270794 647596 270803
rect 647540 270729 647596 270738
rect 649378 269281 649406 983465
rect 649474 277939 649502 993455
rect 649558 987815 649610 987821
rect 649558 987757 649610 987763
rect 649570 941835 649598 987757
rect 649654 987667 649706 987673
rect 649654 987609 649706 987615
rect 649556 941826 649612 941835
rect 649556 941761 649612 941770
rect 649558 927431 649610 927437
rect 649558 927373 649610 927379
rect 649462 277933 649514 277939
rect 649462 277875 649514 277881
rect 649366 269275 649418 269281
rect 649366 269217 649418 269223
rect 646292 266650 646348 266659
rect 646292 266585 646348 266594
rect 635540 265762 635596 265771
rect 635540 265697 635596 265706
rect 633142 265057 633194 265063
rect 633142 264999 633194 265005
rect 639286 256399 639338 256405
rect 639286 256341 639338 256347
rect 632086 253513 632138 253519
rect 632086 253455 632138 253461
rect 625174 253439 625226 253445
rect 625174 253381 625226 253387
rect 497494 251663 497546 251669
rect 497494 251605 497546 251611
rect 501622 251663 501674 251669
rect 501622 251605 501674 251611
rect 212182 247223 212234 247229
rect 212182 247165 212234 247171
rect 216884 246818 216940 246827
rect 212662 246779 212714 246785
rect 227924 246818 227980 246827
rect 216884 246753 216940 246762
rect 221590 246779 221642 246785
rect 212662 246721 212714 246727
rect 212278 246557 212330 246563
rect 212278 246499 212330 246505
rect 212084 244598 212140 244607
rect 212084 244533 212140 244542
rect 211892 233794 211948 233803
rect 211892 233729 211948 233738
rect 211028 233646 211084 233655
rect 211028 233581 211084 233590
rect 211316 233646 211372 233655
rect 211316 233581 211372 233590
rect 211700 233646 211756 233655
rect 211700 233581 211756 233590
rect 211714 233521 211742 233581
rect 211412 233498 211468 233507
rect 210946 233456 211412 233484
rect 211570 233493 211742 233521
rect 211570 233470 211598 233493
rect 211906 233470 211934 233729
rect 212180 233646 212236 233655
rect 212180 233581 212236 233590
rect 212194 233484 212222 233581
rect 212290 233484 212318 246499
rect 212386 243719 212414 246494
rect 212372 243710 212428 243719
rect 212372 243645 212428 243654
rect 212374 233681 212426 233687
rect 212374 233623 212426 233629
rect 212194 233470 212318 233484
rect 212386 233484 212414 233623
rect 212674 233484 212702 246721
rect 212770 240865 212798 246494
rect 213142 245743 213194 245749
rect 213142 245685 213194 245691
rect 212758 240859 212810 240865
rect 212758 240801 212810 240807
rect 213046 236197 213098 236203
rect 213046 236139 213098 236145
rect 212386 233470 212702 233484
rect 213058 233470 213086 236139
rect 213154 233539 213182 245685
rect 213250 235135 213278 246494
rect 213696 246480 213950 246508
rect 214080 246480 214334 246508
rect 213526 244855 213578 244861
rect 213526 244797 213578 244803
rect 213236 235126 213292 235135
rect 213236 235061 213292 235070
rect 213538 233613 213566 244797
rect 213922 241457 213950 246480
rect 214198 245003 214250 245009
rect 214198 244945 214250 244951
rect 214102 244929 214154 244935
rect 214102 244871 214154 244877
rect 213910 241451 213962 241457
rect 213910 241393 213962 241399
rect 213526 233607 213578 233613
rect 213526 233549 213578 233555
rect 213142 233533 213194 233539
rect 213538 233484 213566 233549
rect 213910 233533 213962 233539
rect 213194 233481 213408 233484
rect 213142 233475 213408 233481
rect 212194 233456 212304 233470
rect 212386 233456 212688 233470
rect 213154 233456 213408 233475
rect 213538 233456 213792 233484
rect 214114 233484 214142 244871
rect 213962 233481 214142 233484
rect 213910 233475 214142 233481
rect 213922 233470 214142 233475
rect 214210 233484 214238 244945
rect 214306 243571 214334 246480
rect 214292 243562 214348 243571
rect 214292 243497 214348 243506
rect 214498 239681 214526 246494
rect 214486 239675 214538 239681
rect 214486 239617 214538 239623
rect 214868 237790 214924 237799
rect 214868 237725 214924 237734
rect 214292 233498 214348 233507
rect 213922 233456 214128 233470
rect 214210 233456 214292 233484
rect 211412 233433 211468 233442
rect 214348 233456 214512 233484
rect 214882 233470 214910 237725
rect 214978 234987 215006 246494
rect 215458 241679 215486 246494
rect 215808 246480 215966 246508
rect 216288 246480 216542 246508
rect 215446 241673 215498 241679
rect 215446 241615 215498 241621
rect 215938 239311 215966 246480
rect 216514 245009 216542 246480
rect 216502 245003 216554 245009
rect 216502 244945 216554 244951
rect 216706 241013 216734 246494
rect 216898 245749 216926 246753
rect 246452 246818 246508 246827
rect 227924 246753 227980 246762
rect 228214 246779 228266 246785
rect 221590 246721 221642 246727
rect 221602 246563 221630 246721
rect 226390 246705 226442 246711
rect 226390 246647 226442 246653
rect 226006 246631 226058 246637
rect 226006 246573 226058 246579
rect 221590 246557 221642 246563
rect 216886 245743 216938 245749
rect 216886 245685 216938 245691
rect 216694 241007 216746 241013
rect 216694 240949 216746 240955
rect 215926 239305 215978 239311
rect 215926 239247 215978 239253
rect 216694 239009 216746 239015
rect 216694 238951 216746 238957
rect 216310 238417 216362 238423
rect 216310 238359 216362 238365
rect 215828 238086 215884 238095
rect 215828 238021 215884 238030
rect 215252 237938 215308 237947
rect 215252 237873 215308 237882
rect 214964 234978 215020 234987
rect 214964 234913 215020 234922
rect 215266 233470 215294 237873
rect 215842 233484 215870 238021
rect 215924 237642 215980 237651
rect 215924 237577 215980 237586
rect 215616 233456 215870 233484
rect 215938 233484 215966 237577
rect 215938 233456 216000 233484
rect 216322 233470 216350 238359
rect 216706 233470 216734 238951
rect 217078 238639 217130 238645
rect 217078 238581 217130 238587
rect 217090 233470 217118 238581
rect 217186 235875 217214 246494
rect 217570 241827 217598 246494
rect 218016 246480 218270 246508
rect 218496 246480 218750 246508
rect 218928 246480 219230 246508
rect 218242 243867 218270 246480
rect 218228 243858 218284 243867
rect 218228 243793 218284 243802
rect 217558 241821 217610 241827
rect 217558 241763 217610 241769
rect 218518 240415 218570 240421
rect 218518 240357 218570 240363
rect 218422 240193 218474 240199
rect 218422 240135 218474 240141
rect 218038 238491 218090 238497
rect 218038 238433 218090 238439
rect 217462 236863 217514 236869
rect 217462 236805 217514 236811
rect 217172 235866 217228 235875
rect 217172 235801 217228 235810
rect 217474 233470 217502 236805
rect 218050 233484 218078 238433
rect 218434 233484 218462 240135
rect 217824 233456 218078 233484
rect 218208 233456 218462 233484
rect 218530 233470 218558 240357
rect 218722 239829 218750 246480
rect 218710 239823 218762 239829
rect 218710 239765 218762 239771
rect 218902 239305 218954 239311
rect 218902 239247 218954 239253
rect 218914 233470 218942 239247
rect 219202 235283 219230 246480
rect 219298 241753 219326 246494
rect 219778 244015 219806 246494
rect 220224 246480 220478 246508
rect 220608 246480 220862 246508
rect 221590 246499 221642 246505
rect 219764 244006 219820 244015
rect 219764 243941 219820 243950
rect 219286 241747 219338 241753
rect 219286 241689 219338 241695
rect 220450 241605 220478 246480
rect 220438 241599 220490 241605
rect 220438 241541 220490 241547
rect 219286 240785 219338 240791
rect 219286 240727 219338 240733
rect 219188 235274 219244 235283
rect 219188 235209 219244 235218
rect 219298 233470 219326 240727
rect 219670 240637 219722 240643
rect 219670 240579 219722 240585
rect 219682 233470 219710 240579
rect 220630 240563 220682 240569
rect 220630 240505 220682 240511
rect 220246 240489 220298 240495
rect 220246 240431 220298 240437
rect 220258 233484 220286 240431
rect 220642 233484 220670 240505
rect 220726 236937 220778 236943
rect 220726 236879 220778 236885
rect 220032 233456 220286 233484
rect 220416 233456 220670 233484
rect 220738 233470 220766 236879
rect 220834 235579 220862 246480
rect 221026 244459 221054 246494
rect 221012 244450 221068 244459
rect 221012 244385 221068 244394
rect 221506 239977 221534 246494
rect 222000 246480 222206 246508
rect 222336 246480 222590 246508
rect 222816 246480 223070 246508
rect 221494 239971 221546 239977
rect 221494 239913 221546 239919
rect 221878 237825 221930 237831
rect 221878 237767 221930 237773
rect 221494 237751 221546 237757
rect 221494 237693 221546 237699
rect 221110 237085 221162 237091
rect 221110 237027 221162 237033
rect 220820 235570 220876 235579
rect 220820 235505 220876 235514
rect 221122 233470 221150 237027
rect 221506 233470 221534 237693
rect 221890 233470 221918 237767
rect 221974 237603 222026 237609
rect 221974 237545 222026 237551
rect 221986 233484 222014 237545
rect 222178 235431 222206 246480
rect 222454 246261 222506 246267
rect 222454 246203 222506 246209
rect 222466 245453 222494 246203
rect 222454 245447 222506 245453
rect 222454 245389 222506 245395
rect 222562 241087 222590 246480
rect 223042 242979 223070 246480
rect 223028 242970 223084 242979
rect 223028 242905 223084 242914
rect 223234 241531 223262 246494
rect 223728 246480 224030 246508
rect 223222 241525 223274 241531
rect 223222 241467 223274 241473
rect 222550 241081 222602 241087
rect 222550 241023 222602 241029
rect 222838 238047 222890 238053
rect 222838 237989 222890 237995
rect 222164 235422 222220 235431
rect 222164 235357 222220 235366
rect 222850 233484 222878 237989
rect 223318 237973 223370 237979
rect 223318 237915 223370 237921
rect 222934 237899 222986 237905
rect 222934 237841 222986 237847
rect 221986 233456 222240 233484
rect 222624 233456 222878 233484
rect 222946 233470 222974 237841
rect 223330 233470 223358 237915
rect 223702 237603 223754 237609
rect 223702 237545 223754 237551
rect 223714 233470 223742 237545
rect 224002 235727 224030 246480
rect 224098 241235 224126 246494
rect 224544 246480 224606 246508
rect 225024 246480 225278 246508
rect 224578 243127 224606 246480
rect 224564 243118 224620 243127
rect 224564 243053 224620 243062
rect 224086 241229 224138 241235
rect 224086 241171 224138 241177
rect 225250 241161 225278 246480
rect 225238 241155 225290 241161
rect 225238 241097 225290 241103
rect 225442 240273 225470 246494
rect 225826 244163 225854 246494
rect 226018 246193 226046 246573
rect 226006 246187 226058 246193
rect 226006 246129 226058 246135
rect 225812 244154 225868 244163
rect 225812 244089 225868 244098
rect 225430 240267 225482 240273
rect 225430 240209 225482 240215
rect 226306 240125 226334 246494
rect 226402 244755 226430 246647
rect 226752 246480 227006 246508
rect 227232 246480 227390 246508
rect 227568 246480 227870 246508
rect 226388 244746 226444 244755
rect 226388 244681 226444 244690
rect 226294 240119 226346 240125
rect 226294 240061 226346 240067
rect 225142 239675 225194 239681
rect 225142 239617 225194 239623
rect 224566 238787 224618 238793
rect 224566 238729 224618 238735
rect 224086 237677 224138 237683
rect 224086 237619 224138 237625
rect 223988 235718 224044 235727
rect 223988 235653 224044 235662
rect 224098 233470 224126 237619
rect 224578 233484 224606 238729
rect 225046 236493 225098 236499
rect 225046 236435 225098 236441
rect 225058 233484 225086 236435
rect 224448 233456 224606 233484
rect 224832 233456 225086 233484
rect 225154 233470 225182 239617
rect 226294 239601 226346 239607
rect 226294 239543 226346 239549
rect 225526 237307 225578 237313
rect 225526 237249 225578 237255
rect 225538 233470 225566 237249
rect 225910 236197 225962 236203
rect 225910 236139 225962 236145
rect 225922 233470 225950 236139
rect 226306 233470 226334 239543
rect 226870 238861 226922 238867
rect 226870 238803 226922 238809
rect 226882 233484 226910 238803
rect 226978 234723 227006 246480
rect 227062 245077 227114 245083
rect 227060 245042 227062 245051
rect 227114 245042 227116 245051
rect 227060 244977 227116 244986
rect 227362 240939 227390 246480
rect 227542 245595 227594 245601
rect 227542 245537 227594 245543
rect 227446 245151 227498 245157
rect 227446 245093 227498 245099
rect 227458 244755 227486 245093
rect 227444 244746 227500 244755
rect 227444 244681 227500 244690
rect 227554 244607 227582 245537
rect 227638 244781 227690 244787
rect 227636 244746 227638 244755
rect 227690 244746 227692 244755
rect 227636 244681 227692 244690
rect 227540 244598 227596 244607
rect 227540 244533 227596 244542
rect 227842 243381 227870 246480
rect 227938 245083 227966 246753
rect 228214 246721 228266 246727
rect 229654 246779 229706 246785
rect 229654 246721 229706 246727
rect 243094 246779 243146 246785
rect 243094 246721 243146 246727
rect 246166 246779 246218 246785
rect 246452 246753 246508 246762
rect 247796 246818 247852 246827
rect 247796 246753 247852 246762
rect 248372 246818 248428 246827
rect 259220 246818 259276 246827
rect 248372 246753 248428 246762
rect 254038 246779 254090 246785
rect 246166 246721 246218 246727
rect 227926 245077 227978 245083
rect 227926 245019 227978 245025
rect 227830 243375 227882 243381
rect 227830 243317 227882 243323
rect 227350 240933 227402 240939
rect 227350 240875 227402 240881
rect 228034 239755 228062 246494
rect 228226 246341 228254 246721
rect 229666 246563 229694 246721
rect 229654 246557 229706 246563
rect 228310 246483 228362 246489
rect 228528 246480 228638 246508
rect 228310 246425 228362 246431
rect 228322 246341 228350 246425
rect 228214 246335 228266 246341
rect 228214 246277 228266 246283
rect 228310 246335 228362 246341
rect 228310 246277 228362 246283
rect 228214 245743 228266 245749
rect 228214 245685 228266 245691
rect 228116 245042 228172 245051
rect 228116 244977 228172 244986
rect 228130 244787 228158 244977
rect 228118 244781 228170 244787
rect 228226 244755 228254 245685
rect 228118 244723 228170 244729
rect 228212 244746 228268 244755
rect 228212 244681 228268 244690
rect 228022 239749 228074 239755
rect 228022 239691 228074 239697
rect 228118 239009 228170 239015
rect 228118 238951 228170 238957
rect 227350 237233 227402 237239
rect 227350 237175 227402 237181
rect 227254 237011 227306 237017
rect 227254 236953 227306 236959
rect 226966 234717 227018 234723
rect 226966 234659 227018 234665
rect 227266 233484 227294 236953
rect 226656 233456 226910 233484
rect 227040 233456 227294 233484
rect 227362 233470 227390 237175
rect 227734 236271 227786 236277
rect 227734 236213 227786 236219
rect 227746 233470 227774 236213
rect 228130 233470 228158 238951
rect 228214 238121 228266 238127
rect 228214 238063 228266 238069
rect 228226 237757 228254 238063
rect 228502 237899 228554 237905
rect 228502 237841 228554 237847
rect 228214 237751 228266 237757
rect 228214 237693 228266 237699
rect 228514 233470 228542 237841
rect 228610 236171 228638 246480
rect 228694 246483 228746 246489
rect 228864 246480 229214 246508
rect 229344 246480 229598 246508
rect 229654 246499 229706 246505
rect 229942 246557 229994 246563
rect 229942 246499 229994 246505
rect 228694 246425 228746 246431
rect 228706 246193 228734 246425
rect 228694 246187 228746 246193
rect 228694 246129 228746 246135
rect 229186 241624 229214 246480
rect 229570 244607 229598 246480
rect 229556 244598 229612 244607
rect 229556 244533 229612 244542
rect 229186 241596 229406 241624
rect 229174 241451 229226 241457
rect 229174 241393 229226 241399
rect 229078 239675 229130 239681
rect 229078 239617 229130 239623
rect 228596 236162 228652 236171
rect 228596 236097 228652 236106
rect 229090 233484 229118 239617
rect 228864 233456 229118 233484
rect 229186 233484 229214 241393
rect 229378 233484 229406 241596
rect 229762 236023 229790 246494
rect 229954 246341 229982 246499
rect 229942 246335 229994 246341
rect 229942 246277 229994 246283
rect 229942 239749 229994 239755
rect 229942 239691 229994 239697
rect 229748 236014 229804 236023
rect 229748 235949 229804 235958
rect 229186 233456 229248 233484
rect 229378 233456 229584 233484
rect 229954 233470 229982 239691
rect 230242 239681 230270 246494
rect 230626 243455 230654 246494
rect 230818 246480 231072 246508
rect 231552 246480 231710 246508
rect 230614 243449 230666 243455
rect 230614 243391 230666 243397
rect 230326 240933 230378 240939
rect 230326 240875 230378 240881
rect 230230 239675 230282 239681
rect 230230 239617 230282 239623
rect 230338 233470 230366 240875
rect 230710 240119 230762 240125
rect 230710 240061 230762 240067
rect 230722 233470 230750 240061
rect 230818 237905 230846 246480
rect 231190 241155 231242 241161
rect 231190 241097 231242 241103
rect 230902 240267 230954 240273
rect 230902 240209 230954 240215
rect 230806 237899 230858 237905
rect 230806 237841 230858 237847
rect 230914 233484 230942 240209
rect 231202 233484 231230 241097
rect 231682 234797 231710 246480
rect 231766 241229 231818 241235
rect 231766 241171 231818 241177
rect 231670 234791 231722 234797
rect 231670 234733 231722 234739
rect 230914 233456 231072 233484
rect 231202 233456 231456 233484
rect 231778 233470 231806 241171
rect 231970 239015 231998 246494
rect 232354 243275 232382 246494
rect 232340 243266 232396 243275
rect 232340 243201 232396 243210
rect 232150 241525 232202 241531
rect 232150 241467 232202 241473
rect 231958 239009 232010 239015
rect 231958 238951 232010 238957
rect 232162 233470 232190 241467
rect 232534 241081 232586 241087
rect 232534 241023 232586 241029
rect 232546 233470 232574 241023
rect 232834 236277 232862 246494
rect 233280 246480 233342 246508
rect 233314 241235 233342 246480
rect 233506 246480 233760 246508
rect 233398 241599 233450 241605
rect 233398 241541 233450 241547
rect 233302 241229 233354 241235
rect 233302 241171 233354 241177
rect 233206 240859 233258 240865
rect 233206 240801 233258 240807
rect 232918 239971 232970 239977
rect 232918 239913 232970 239919
rect 232822 236271 232874 236277
rect 232822 236213 232874 236219
rect 232930 233470 232958 239913
rect 233218 233780 233246 240801
rect 233218 233752 233294 233780
rect 233266 233470 233294 233752
rect 233410 233484 233438 241541
rect 233506 237239 233534 246480
rect 233974 241747 234026 241753
rect 233974 241689 234026 241695
rect 233494 237233 233546 237239
rect 233494 237175 233546 237181
rect 233410 233456 233664 233484
rect 233986 233470 234014 241689
rect 234082 237017 234110 246494
rect 234562 239903 234590 246494
rect 234742 241821 234794 241827
rect 234742 241763 234794 241769
rect 234550 239897 234602 239903
rect 234550 239839 234602 239845
rect 234358 239823 234410 239829
rect 234358 239765 234410 239771
rect 234070 237011 234122 237017
rect 234070 236953 234122 236959
rect 234370 233470 234398 239765
rect 234754 233470 234782 241763
rect 235042 238867 235070 246494
rect 235488 246480 235742 246508
rect 235126 244633 235178 244639
rect 235126 244575 235178 244581
rect 235030 238861 235082 238867
rect 235030 238803 235082 238809
rect 235138 233470 235166 244575
rect 235606 243301 235658 243307
rect 235606 243243 235658 243249
rect 235618 233484 235646 243243
rect 235714 242091 235742 246480
rect 235858 246212 235886 246494
rect 235810 246184 235886 246212
rect 235700 242082 235756 242091
rect 235700 242017 235756 242026
rect 235810 239607 235838 246184
rect 236182 241007 236234 241013
rect 236182 240949 236234 240955
rect 235798 239601 235850 239607
rect 235798 239543 235850 239549
rect 236194 239089 236222 240949
rect 236290 240051 236318 246494
rect 236470 240119 236522 240125
rect 236470 240061 236522 240067
rect 236278 240045 236330 240051
rect 236278 239987 236330 239993
rect 236182 239083 236234 239089
rect 236182 239025 236234 239031
rect 236086 235457 236138 235463
rect 236086 235399 236138 235405
rect 236098 233484 236126 235399
rect 236482 233484 236510 240061
rect 236566 236271 236618 236277
rect 236566 236213 236618 236219
rect 235488 233456 235646 233484
rect 235872 233456 236126 233484
rect 236208 233456 236510 233484
rect 236578 233470 236606 236213
rect 236770 236203 236798 246494
rect 237154 243603 237182 246494
rect 237442 246480 237600 246508
rect 238080 246480 238238 246508
rect 237142 243597 237194 243603
rect 237142 243539 237194 243545
rect 236950 241525 237002 241531
rect 236950 241467 237002 241473
rect 236758 236197 236810 236203
rect 236758 236139 236810 236145
rect 236962 233470 236990 241467
rect 237334 240341 237386 240347
rect 237334 240283 237386 240289
rect 237346 233470 237374 240283
rect 237442 237313 237470 246480
rect 237718 241599 237770 241605
rect 237718 241541 237770 241547
rect 237526 239009 237578 239015
rect 237526 238951 237578 238957
rect 237538 238423 237566 238951
rect 237526 238417 237578 238423
rect 237526 238359 237578 238365
rect 237430 237307 237482 237313
rect 237430 237249 237482 237255
rect 237730 233780 237758 241541
rect 237910 240933 237962 240939
rect 237910 240875 237962 240881
rect 237814 240859 237866 240865
rect 237814 240801 237866 240807
rect 237826 240421 237854 240801
rect 237814 240415 237866 240421
rect 237814 240357 237866 240363
rect 237922 240199 237950 240875
rect 237910 240193 237962 240199
rect 237910 240135 237962 240141
rect 238210 239681 238238 246480
rect 238498 241901 238526 246494
rect 238486 241895 238538 241901
rect 238486 241837 238538 241843
rect 238678 241229 238730 241235
rect 238678 241171 238730 241177
rect 238294 239971 238346 239977
rect 238294 239913 238346 239919
rect 238198 239675 238250 239681
rect 238198 239617 238250 239623
rect 237682 233752 237758 233780
rect 237682 233470 237710 233752
rect 238306 233484 238334 239913
rect 238582 239897 238634 239903
rect 238582 239839 238634 239845
rect 238390 239083 238442 239089
rect 238390 239025 238442 239031
rect 238080 233456 238334 233484
rect 238402 233470 238430 239025
rect 238594 234871 238622 239839
rect 238690 235093 238718 241171
rect 238774 240267 238826 240273
rect 238774 240209 238826 240215
rect 238678 235087 238730 235093
rect 238678 235029 238730 235035
rect 238582 234865 238634 234871
rect 238582 234807 238634 234813
rect 238786 233470 238814 240209
rect 238882 236499 238910 246494
rect 238966 240415 239018 240421
rect 238966 240357 239018 240363
rect 238870 236493 238922 236499
rect 238870 236435 238922 236441
rect 238978 236277 239006 240357
rect 239158 238861 239210 238867
rect 239158 238803 239210 238809
rect 238966 236271 239018 236277
rect 238966 236213 239018 236219
rect 239170 233470 239198 238803
rect 239362 235315 239390 246494
rect 239554 246480 239808 246508
rect 240288 246480 240542 246508
rect 239554 238793 239582 246480
rect 240514 243529 240542 246480
rect 240658 246212 240686 246494
rect 240658 246184 240734 246212
rect 240502 243523 240554 243529
rect 240502 243465 240554 243471
rect 240502 239231 240554 239237
rect 240502 239173 240554 239179
rect 240118 238935 240170 238941
rect 240118 238877 240170 238883
rect 239542 238787 239594 238793
rect 239542 238729 239594 238735
rect 239542 237381 239594 237387
rect 239542 237323 239594 237329
rect 239350 235309 239402 235315
rect 239350 235251 239402 235257
rect 239554 233470 239582 237323
rect 240130 233484 240158 238877
rect 240514 233484 240542 239173
rect 240598 238417 240650 238423
rect 240598 238359 240650 238365
rect 239904 233456 240158 233484
rect 240288 233456 240542 233484
rect 240610 233470 240638 238359
rect 240706 237683 240734 246184
rect 240980 240602 241036 240611
rect 240980 240537 241036 240546
rect 240694 237677 240746 237683
rect 240694 237619 240746 237625
rect 240994 233470 241022 240537
rect 241090 239755 241118 246494
rect 241078 239749 241130 239755
rect 241078 239691 241130 239697
rect 241364 238234 241420 238243
rect 241364 238169 241420 238178
rect 241378 233470 241406 238169
rect 241570 237609 241598 246494
rect 242016 246480 242270 246508
rect 242242 244565 242270 246480
rect 242386 246212 242414 246494
rect 242626 246480 242880 246508
rect 242386 246184 242462 246212
rect 242230 244559 242282 244565
rect 242230 244501 242282 244507
rect 241748 240750 241804 240759
rect 241748 240685 241804 240694
rect 241654 240045 241706 240051
rect 241654 239987 241706 239993
rect 241558 237603 241610 237609
rect 241558 237545 241610 237551
rect 241666 235019 241694 239987
rect 241654 235013 241706 235019
rect 241654 234955 241706 234961
rect 241762 233470 241790 240685
rect 241846 239675 241898 239681
rect 241846 239617 241898 239623
rect 241858 235167 241886 239617
rect 242324 238382 242380 238391
rect 242324 238317 242380 238326
rect 241846 235161 241898 235167
rect 241846 235103 241898 235109
rect 242338 233484 242366 238317
rect 242434 237979 242462 246184
rect 242422 237973 242474 237979
rect 242422 237915 242474 237921
rect 242626 237831 242654 246480
rect 243106 246193 243134 246721
rect 243382 246705 243434 246711
rect 243382 246647 243434 246653
rect 243190 246557 243242 246563
rect 243190 246499 243242 246505
rect 243094 246187 243146 246193
rect 243094 246129 243146 246135
rect 243202 245971 243230 246499
rect 243190 245965 243242 245971
rect 243190 245907 243242 245913
rect 243298 243899 243326 246494
rect 243394 245749 243422 246647
rect 243382 245743 243434 245749
rect 243382 245685 243434 245691
rect 243286 243893 243338 243899
rect 243286 243835 243338 243841
rect 243188 241194 243244 241203
rect 243188 241129 243244 241138
rect 242708 241046 242764 241055
rect 242708 240981 242764 240990
rect 242614 237825 242666 237831
rect 242614 237767 242666 237773
rect 242722 233484 242750 240981
rect 242804 238678 242860 238687
rect 242804 238613 242860 238622
rect 242112 233456 242366 233484
rect 242496 233456 242750 233484
rect 242818 233470 242846 238613
rect 243202 233470 243230 241129
rect 243572 238826 243628 238835
rect 243572 238761 243628 238770
rect 243586 233470 243614 238761
rect 243778 238053 243806 246494
rect 243956 241342 244012 241351
rect 243956 241277 244012 241286
rect 243766 238047 243818 238053
rect 243766 237989 243818 237995
rect 243970 233470 243998 241277
rect 244162 240199 244190 246494
rect 244608 246480 244766 246508
rect 244738 243825 244766 246480
rect 244834 246480 245088 246508
rect 245424 246480 245726 246508
rect 244726 243819 244778 243825
rect 244726 243761 244778 243767
rect 244438 241007 244490 241013
rect 244438 240949 244490 240955
rect 244150 240193 244202 240199
rect 244150 240135 244202 240141
rect 244340 238974 244396 238983
rect 244340 238909 244396 238918
rect 244354 233780 244382 238909
rect 244306 233752 244382 233780
rect 244306 233470 244334 233752
rect 244450 233484 244478 240949
rect 244630 239749 244682 239755
rect 244630 239691 244682 239697
rect 244642 234945 244670 239691
rect 244834 237757 244862 246480
rect 245396 241786 245452 241795
rect 245396 241721 245452 241730
rect 244822 237751 244874 237757
rect 244822 237693 244874 237699
rect 245014 237603 245066 237609
rect 245014 237545 245066 237551
rect 244630 234939 244682 234945
rect 244630 234881 244682 234887
rect 244450 233456 244704 233484
rect 245026 233470 245054 237545
rect 245410 233470 245438 241721
rect 245698 235389 245726 246480
rect 245890 238127 245918 246494
rect 246178 245897 246206 246721
rect 246166 245891 246218 245897
rect 246166 245833 246218 245839
rect 246370 243751 246398 246494
rect 246466 245083 246494 246753
rect 247810 246637 247838 246753
rect 248278 246705 248330 246711
rect 248278 246647 248330 246653
rect 247702 246631 247754 246637
rect 247702 246573 247754 246579
rect 247798 246631 247850 246637
rect 247798 246573 247850 246579
rect 246562 246480 246816 246508
rect 246946 246480 247200 246508
rect 247330 246480 247632 246508
rect 246454 245077 246506 245083
rect 246454 245019 246506 245025
rect 246358 243745 246410 243751
rect 246358 243687 246410 243693
rect 246164 241934 246220 241943
rect 246164 241869 246220 241878
rect 245878 238121 245930 238127
rect 245878 238063 245930 238069
rect 245782 237751 245834 237757
rect 245782 237693 245834 237699
rect 245686 235383 245738 235389
rect 245686 235325 245738 235331
rect 245794 233470 245822 237693
rect 246178 233470 246206 241869
rect 246358 240193 246410 240199
rect 246358 240135 246410 240141
rect 246370 235241 246398 240135
rect 246562 237091 246590 246480
rect 246742 237677 246794 237683
rect 246742 237619 246794 237625
rect 246550 237085 246602 237091
rect 246550 237027 246602 237033
rect 246358 235235 246410 235241
rect 246358 235177 246410 235183
rect 246754 233484 246782 237619
rect 246946 236943 246974 246480
rect 247330 243677 247358 246480
rect 247714 246341 247742 246573
rect 247906 246480 248112 246508
rect 248182 246483 248234 246489
rect 247702 246335 247754 246341
rect 247702 246277 247754 246283
rect 247606 245225 247658 245231
rect 247606 245167 247658 245173
rect 247508 245042 247564 245051
rect 247618 245028 247646 245167
rect 247700 245042 247756 245051
rect 247618 245000 247700 245028
rect 247508 244977 247564 244986
rect 247700 244977 247756 244986
rect 247522 244755 247550 244977
rect 247702 244929 247754 244935
rect 247702 244871 247754 244877
rect 247714 244755 247742 244871
rect 247508 244746 247564 244755
rect 247508 244681 247564 244690
rect 247700 244746 247756 244755
rect 247700 244681 247756 244690
rect 247318 243671 247370 243677
rect 247318 243613 247370 243619
rect 247906 240569 247934 246480
rect 248182 246425 248234 246431
rect 248194 245971 248222 246425
rect 248290 246193 248318 246647
rect 248278 246187 248330 246193
rect 248278 246129 248330 246135
rect 248182 245965 248234 245971
rect 248182 245907 248234 245913
rect 248386 245897 248414 246753
rect 267956 246818 268012 246827
rect 259220 246753 259276 246762
rect 267478 246779 267530 246785
rect 254038 246721 254090 246727
rect 248374 245891 248426 245897
rect 248374 245833 248426 245839
rect 247990 245595 248042 245601
rect 247990 245537 248042 245543
rect 248002 244861 248030 245537
rect 248086 245077 248138 245083
rect 248086 245019 248138 245025
rect 247990 244855 248042 244861
rect 247990 244797 248042 244803
rect 248098 244787 248126 245019
rect 248086 244781 248138 244787
rect 248086 244723 248138 244729
rect 248578 241827 248606 246494
rect 248674 246480 248928 246508
rect 249408 246480 249662 246508
rect 248566 241821 248618 241827
rect 248566 241763 248618 241769
rect 247894 240563 247946 240569
rect 247894 240505 247946 240511
rect 248374 240563 248426 240569
rect 248374 240505 248426 240511
rect 247124 240306 247180 240315
rect 247124 240241 247180 240250
rect 246934 236937 246986 236943
rect 246934 236879 246986 236885
rect 247138 233484 247166 240241
rect 247604 240158 247660 240167
rect 247604 240093 247660 240102
rect 247222 237825 247274 237831
rect 247222 237767 247274 237773
rect 246528 233456 246782 233484
rect 246912 233456 247166 233484
rect 247234 233470 247262 237767
rect 247618 233470 247646 240093
rect 247990 237899 248042 237905
rect 247990 237841 248042 237847
rect 248002 233470 248030 237841
rect 248386 233470 248414 240505
rect 248674 240495 248702 246480
rect 249634 244047 249662 246480
rect 249622 244041 249674 244047
rect 249622 243983 249674 243989
rect 249826 241087 249854 246494
rect 250306 241901 250334 246494
rect 250294 241895 250346 241901
rect 250294 241837 250346 241843
rect 250690 241161 250718 246494
rect 251136 246480 251390 246508
rect 251616 246480 251870 246508
rect 251362 244121 251390 246480
rect 251842 245823 251870 246480
rect 251830 245817 251882 245823
rect 251830 245759 251882 245765
rect 251350 244115 251402 244121
rect 251350 244057 251402 244063
rect 250678 241155 250730 241161
rect 250678 241097 250730 241103
rect 249814 241081 249866 241087
rect 249814 241023 249866 241029
rect 252034 240865 252062 246494
rect 252418 245453 252446 246494
rect 252406 245447 252458 245453
rect 252406 245389 252458 245395
rect 252790 241451 252842 241457
rect 252790 241393 252842 241399
rect 252022 240859 252074 240865
rect 252022 240801 252074 240807
rect 252310 240859 252362 240865
rect 252310 240801 252362 240807
rect 251542 240785 251594 240791
rect 251542 240727 251594 240733
rect 249814 240711 249866 240717
rect 249814 240653 249866 240659
rect 248662 240489 248714 240495
rect 248662 240431 248714 240437
rect 249334 240489 249386 240495
rect 249334 240431 249386 240437
rect 248950 237455 249002 237461
rect 248950 237397 249002 237403
rect 248962 233484 248990 237397
rect 249346 233484 249374 240431
rect 249430 238047 249482 238053
rect 249430 237989 249482 237995
rect 248736 233456 248990 233484
rect 249120 233456 249374 233484
rect 249442 233470 249470 237989
rect 249826 233470 249854 240653
rect 250582 240637 250634 240643
rect 250582 240579 250634 240585
rect 250198 237973 250250 237979
rect 250198 237915 250250 237921
rect 250210 233470 250238 237915
rect 250594 233470 250622 240579
rect 251158 238121 251210 238127
rect 251158 238063 251210 238069
rect 251170 233484 251198 238063
rect 251554 233484 251582 240727
rect 251638 238195 251690 238201
rect 251638 238137 251690 238143
rect 250944 233456 251198 233484
rect 251328 233456 251582 233484
rect 251650 233470 251678 238137
rect 252322 233484 252350 240801
rect 252406 238269 252458 238275
rect 252406 238211 252458 238217
rect 252048 233456 252350 233484
rect 252418 233470 252446 238211
rect 252802 233470 252830 241393
rect 252898 240939 252926 246494
rect 253344 246480 253406 246508
rect 253378 245527 253406 246480
rect 253474 246480 253728 246508
rect 253366 245521 253418 245527
rect 253366 245463 253418 245469
rect 252886 240933 252938 240939
rect 252886 240875 252938 240881
rect 253474 238497 253502 246480
rect 254050 245749 254078 246721
rect 254146 245749 254174 246494
rect 254338 246480 254640 246508
rect 254038 245743 254090 245749
rect 254038 245685 254090 245691
rect 254134 245743 254186 245749
rect 254134 245685 254186 245691
rect 254230 241081 254282 241087
rect 254230 241023 254282 241029
rect 253750 240933 253802 240939
rect 253750 240875 253802 240881
rect 253462 238491 253514 238497
rect 253462 238433 253514 238439
rect 253366 238343 253418 238349
rect 253366 238285 253418 238291
rect 253378 233484 253406 238285
rect 253762 233484 253790 240875
rect 253846 238565 253898 238571
rect 253846 238507 253898 238513
rect 253152 233456 253406 233484
rect 253536 233456 253790 233484
rect 253858 233470 253886 238507
rect 254242 233470 254270 241023
rect 254338 236869 254366 246480
rect 255106 241753 255134 246494
rect 255202 246480 255456 246508
rect 255682 246480 255936 246508
rect 255094 241747 255146 241753
rect 255094 241689 255146 241695
rect 254998 241155 255050 241161
rect 254998 241097 255050 241103
rect 254614 238491 254666 238497
rect 254614 238433 254666 238439
rect 254326 236863 254378 236869
rect 254326 236805 254378 236811
rect 254626 233470 254654 238433
rect 255010 233470 255038 241097
rect 255202 238645 255230 246480
rect 255682 239237 255710 246480
rect 255958 241229 256010 241235
rect 255958 241171 256010 241177
rect 255670 239231 255722 239237
rect 255670 239173 255722 239179
rect 255190 238639 255242 238645
rect 255190 238581 255242 238587
rect 255574 238639 255626 238645
rect 255574 238581 255626 238587
rect 255586 233484 255614 238581
rect 255970 233484 255998 241171
rect 256054 238713 256106 238719
rect 256054 238655 256106 238661
rect 255360 233456 255614 233484
rect 255744 233456 255998 233484
rect 256066 233470 256094 238655
rect 256354 235685 256382 246494
rect 256438 240045 256490 240051
rect 256438 239987 256490 239993
rect 256342 235679 256394 235685
rect 256342 235621 256394 235627
rect 256450 233470 256478 239987
rect 256834 238941 256862 246494
rect 257218 244269 257246 246494
rect 257410 246480 257664 246508
rect 258144 246480 258398 246508
rect 257206 244263 257258 244269
rect 257206 244205 257258 244211
rect 257206 240193 257258 240199
rect 257206 240135 257258 240141
rect 256822 238935 256874 238941
rect 256822 238877 256874 238883
rect 256822 237529 256874 237535
rect 256822 237471 256874 237477
rect 256834 233470 256862 237471
rect 257218 233470 257246 240135
rect 257410 237387 257438 246480
rect 257684 244746 257740 244755
rect 257684 244681 257740 244690
rect 257588 244302 257644 244311
rect 257588 244237 257644 244246
rect 257602 243127 257630 244237
rect 257698 244163 257726 244681
rect 257782 244559 257834 244565
rect 257782 244501 257834 244507
rect 257684 244154 257740 244163
rect 257684 244089 257740 244098
rect 257794 243973 257822 244501
rect 257876 244154 257932 244163
rect 257876 244089 257932 244098
rect 257782 243967 257834 243973
rect 257782 243909 257834 243915
rect 257588 243118 257644 243127
rect 257588 243053 257644 243062
rect 257890 242979 257918 244089
rect 257876 242970 257932 242979
rect 257876 242905 257932 242914
rect 258262 238935 258314 238941
rect 258262 238877 258314 238883
rect 257782 238787 257834 238793
rect 257782 238729 257834 238735
rect 257398 237381 257450 237387
rect 257398 237323 257450 237329
rect 257794 233484 257822 238729
rect 258166 236641 258218 236647
rect 258166 236583 258218 236589
rect 258178 233484 258206 236583
rect 257568 233456 257822 233484
rect 257952 233456 258206 233484
rect 258274 233470 258302 238877
rect 258370 235833 258398 246480
rect 258562 238867 258590 246494
rect 258946 244343 258974 246494
rect 259234 244713 259262 246753
rect 291956 246818 292012 246827
rect 268012 246776 268094 246804
rect 267956 246753 268012 246762
rect 267478 246721 267530 246727
rect 266614 246705 266666 246711
rect 266614 246647 266666 246653
rect 259222 244707 259274 244713
rect 259222 244649 259274 244655
rect 258934 244337 258986 244343
rect 258934 244279 258986 244285
rect 258644 240898 258700 240907
rect 258644 240833 258700 240842
rect 258550 238861 258602 238867
rect 258550 238803 258602 238809
rect 258358 235827 258410 235833
rect 258358 235769 258410 235775
rect 258658 233470 258686 240833
rect 259426 240273 259454 246494
rect 259872 246480 260126 246508
rect 260352 246480 260606 246508
rect 259988 241638 260044 241647
rect 259988 241573 260044 241582
rect 259604 241490 259660 241499
rect 259604 241425 259660 241434
rect 259414 240267 259466 240273
rect 259414 240209 259466 240215
rect 258838 238713 258890 238719
rect 258838 238655 258890 238661
rect 258850 237461 258878 238655
rect 259028 238530 259084 238539
rect 259028 238465 259084 238474
rect 258838 237455 258890 237461
rect 258838 237397 258890 237403
rect 259042 233470 259070 238465
rect 259618 233484 259646 241425
rect 260002 233484 260030 241573
rect 260098 235611 260126 246480
rect 260374 245151 260426 245157
rect 260374 245093 260426 245099
rect 260086 235605 260138 235611
rect 260086 235547 260138 235553
rect 260386 233484 260414 245093
rect 260470 245077 260522 245083
rect 260470 245019 260522 245025
rect 259440 233456 259646 233484
rect 259776 233456 260030 233484
rect 260160 233456 260414 233484
rect 260482 233470 260510 245019
rect 260578 244417 260606 246480
rect 260566 244411 260618 244417
rect 260566 244353 260618 244359
rect 260674 239977 260702 246494
rect 260854 245299 260906 245305
rect 260854 245241 260906 245247
rect 260662 239971 260714 239977
rect 260662 239913 260714 239919
rect 260866 233470 260894 245241
rect 261154 235759 261182 246494
rect 261238 245225 261290 245231
rect 261238 245167 261290 245173
rect 261142 235753 261194 235759
rect 261142 235695 261194 235701
rect 261250 233470 261278 245167
rect 261634 241605 261662 246494
rect 261984 246480 262046 246508
rect 261814 245373 261866 245379
rect 261814 245315 261866 245321
rect 261622 241599 261674 241605
rect 261622 241541 261674 241547
rect 261826 233484 261854 245315
rect 262018 244565 262046 246480
rect 262210 246480 262464 246508
rect 262006 244559 262058 244565
rect 262006 244501 262058 244507
rect 262006 241599 262058 241605
rect 262006 241541 262058 241547
rect 262018 233780 262046 241541
rect 262210 240347 262238 246480
rect 262678 245595 262730 245601
rect 262678 245537 262730 245543
rect 262198 240341 262250 240347
rect 262198 240283 262250 240289
rect 262294 240341 262346 240347
rect 262294 240283 262346 240289
rect 262306 236647 262334 240283
rect 262580 240010 262636 240019
rect 262580 239945 262636 239954
rect 262294 236641 262346 236647
rect 262294 236583 262346 236589
rect 261648 233456 261854 233484
rect 261970 233752 262046 233780
rect 261970 233470 261998 233752
rect 262594 233484 262622 239945
rect 262368 233456 262622 233484
rect 262690 233470 262718 245537
rect 262882 235907 262910 246494
rect 263062 245891 263114 245897
rect 263062 245833 263114 245839
rect 262870 235901 262922 235907
rect 262870 235843 262922 235849
rect 263074 233470 263102 245833
rect 263362 241531 263390 246494
rect 263446 246187 263498 246193
rect 263446 246129 263498 246135
rect 263350 241525 263402 241531
rect 263350 241467 263402 241473
rect 263458 233470 263486 246129
rect 263746 242863 263774 246494
rect 263938 246480 264192 246508
rect 264418 246480 264672 246508
rect 263830 245965 263882 245971
rect 263830 245907 263882 245913
rect 263734 242857 263786 242863
rect 263734 242799 263786 242805
rect 263842 233470 263870 245907
rect 263938 240421 263966 246480
rect 264310 241525 264362 241531
rect 264310 241467 264362 241473
rect 263926 240415 263978 240421
rect 263926 240357 263978 240363
rect 264322 233484 264350 241467
rect 264418 240125 264446 246480
rect 265090 242937 265118 246494
rect 265078 242931 265130 242937
rect 265078 242873 265130 242879
rect 264886 242635 264938 242641
rect 264886 242577 264938 242583
rect 264406 240119 264458 240125
rect 264406 240061 264458 240067
rect 264790 236049 264842 236055
rect 264790 235991 264842 235997
rect 264802 233484 264830 235991
rect 264192 233456 264350 233484
rect 264576 233456 264830 233484
rect 264898 233470 264926 242577
rect 265474 235463 265502 246494
rect 265654 239675 265706 239681
rect 265654 239617 265706 239623
rect 265462 235457 265514 235463
rect 265462 235399 265514 235405
rect 265270 234643 265322 234649
rect 265270 234585 265322 234591
rect 265282 233470 265310 234585
rect 265666 233470 265694 239617
rect 265954 236129 265982 246494
rect 266146 246480 266400 246508
rect 266146 243307 266174 246480
rect 266626 246415 266654 246647
rect 267490 246563 267518 246721
rect 267478 246557 267530 246563
rect 266880 246480 267134 246508
rect 267478 246499 267530 246505
rect 267862 246557 267914 246563
rect 267914 246505 267998 246508
rect 267862 246499 267998 246505
rect 266518 246409 266570 246415
rect 266518 246351 266570 246357
rect 266614 246409 266666 246415
rect 266614 246351 266666 246357
rect 266530 245675 266558 246351
rect 266518 245669 266570 245675
rect 266518 245611 266570 245617
rect 266134 243301 266186 243307
rect 266134 243243 266186 243249
rect 266998 243153 267050 243159
rect 266998 243095 267050 243101
rect 265942 236123 265994 236129
rect 265942 236065 265994 236071
rect 266614 234569 266666 234575
rect 266614 234511 266666 234517
rect 266038 234495 266090 234501
rect 266038 234437 266090 234443
rect 266050 233470 266078 234437
rect 266626 233484 266654 234511
rect 267010 233484 267038 243095
rect 267106 243085 267134 246480
rect 267202 244639 267230 246494
rect 267190 244633 267242 244639
rect 267190 244575 267242 244581
rect 267094 243079 267146 243085
rect 267094 243021 267146 243027
rect 267478 243005 267530 243011
rect 267478 242947 267530 242953
rect 267094 234273 267146 234279
rect 267094 234215 267146 234221
rect 266400 233456 266654 233484
rect 266784 233456 267038 233484
rect 267106 233470 267134 234215
rect 267490 233470 267518 242947
rect 267682 235981 267710 246494
rect 267874 246489 267998 246499
rect 267874 246483 268010 246489
rect 267874 246480 267958 246483
rect 267958 246425 268010 246431
rect 267766 246409 267818 246415
rect 268066 246360 268094 246776
rect 269302 246779 269354 246785
rect 269302 246721 269354 246727
rect 288310 246779 288362 246785
rect 288310 246721 288362 246727
rect 288406 246779 288458 246785
rect 288406 246721 288458 246727
rect 290134 246779 290186 246785
rect 290134 246721 290186 246727
rect 291094 246779 291146 246785
rect 291956 246753 292012 246762
rect 292148 246818 292204 246827
rect 307988 246818 308044 246827
rect 292148 246753 292204 246762
rect 292630 246779 292682 246785
rect 291094 246721 291146 246727
rect 268822 246631 268874 246637
rect 268822 246573 268874 246579
rect 268176 246480 268382 246508
rect 268512 246480 268766 246508
rect 267818 246357 268094 246360
rect 267766 246351 268094 246357
rect 267778 246332 268094 246351
rect 268246 244929 268298 244935
rect 268246 244871 268298 244877
rect 267862 244781 267914 244787
rect 267914 244729 267998 244732
rect 267862 244723 267998 244729
rect 267874 244704 267998 244723
rect 268258 244713 268286 244871
rect 267970 244195 267998 244704
rect 268246 244707 268298 244713
rect 268246 244649 268298 244655
rect 267862 244189 267914 244195
rect 267862 244131 267914 244137
rect 267958 244189 268010 244195
rect 267958 244131 268010 244137
rect 267874 242567 267902 244131
rect 267862 242561 267914 242567
rect 267862 242503 267914 242509
rect 268150 239009 268202 239015
rect 268150 238951 268202 238957
rect 268246 239009 268298 239015
rect 268246 238951 268298 238957
rect 268162 237461 268190 238951
rect 268150 237455 268202 237461
rect 268150 237397 268202 237403
rect 267670 235975 267722 235981
rect 267670 235917 267722 235923
rect 267862 234199 267914 234205
rect 267862 234141 267914 234147
rect 267874 233470 267902 234141
rect 268258 233470 268286 238951
rect 268354 236647 268382 246480
rect 268738 239977 268766 246480
rect 268834 244787 268862 246573
rect 269206 246557 269258 246563
rect 268992 246480 269150 246508
rect 269206 246499 269258 246505
rect 268822 244781 268874 244787
rect 268822 244723 268874 244729
rect 268726 239971 268778 239977
rect 268726 239913 268778 239919
rect 268342 236641 268394 236647
rect 268342 236583 268394 236589
rect 268822 234125 268874 234131
rect 268822 234067 268874 234073
rect 268834 233484 268862 234067
rect 269122 233613 269150 246480
rect 269218 245675 269246 246499
rect 269314 246267 269342 246721
rect 280822 246631 280874 246637
rect 280822 246573 280874 246579
rect 287842 246591 288158 246619
rect 269302 246261 269354 246267
rect 269302 246203 269354 246209
rect 269206 245669 269258 245675
rect 269206 245611 269258 245617
rect 269206 242339 269258 242345
rect 269206 242281 269258 242287
rect 269110 233607 269162 233613
rect 269110 233549 269162 233555
rect 269218 233484 269246 242281
rect 269410 239755 269438 246494
rect 269686 242487 269738 242493
rect 269686 242429 269738 242435
rect 269398 239749 269450 239755
rect 269398 239691 269450 239697
rect 269302 234051 269354 234057
rect 269302 233993 269354 233999
rect 268608 233456 268862 233484
rect 268992 233456 269246 233484
rect 269314 233470 269342 233993
rect 269698 233470 269726 242429
rect 269890 233909 269918 246494
rect 270166 243301 270218 243307
rect 270166 243243 270218 243249
rect 270178 239681 270206 243243
rect 270274 239681 270302 246494
rect 270720 246480 270878 246508
rect 270850 242789 270878 246480
rect 270946 246480 271200 246508
rect 270838 242783 270890 242789
rect 270838 242725 270890 242731
rect 270454 242191 270506 242197
rect 270454 242133 270506 242139
rect 270166 239675 270218 239681
rect 270166 239617 270218 239623
rect 270262 239675 270314 239681
rect 270262 239617 270314 239623
rect 269878 233903 269930 233909
rect 269878 233845 269930 233851
rect 270262 233607 270314 233613
rect 270262 233549 270314 233555
rect 270274 233484 270302 233549
rect 270096 233456 270302 233484
rect 270466 233470 270494 242133
rect 270946 239015 270974 246480
rect 271618 246267 271646 246494
rect 271606 246261 271658 246267
rect 271606 246203 271658 246209
rect 272002 241531 272030 246494
rect 271990 241525 272042 241531
rect 271990 241467 272042 241473
rect 272278 239675 272330 239681
rect 272278 239617 272330 239623
rect 271414 239601 271466 239607
rect 271414 239543 271466 239549
rect 270934 239009 270986 239015
rect 270934 238951 270986 238957
rect 271030 236937 271082 236943
rect 271030 236879 271082 236885
rect 271042 233484 271070 236879
rect 271426 233484 271454 239543
rect 271894 239083 271946 239089
rect 271894 239025 271946 239031
rect 271510 236345 271562 236351
rect 271510 236287 271562 236293
rect 270816 233456 271070 233484
rect 271200 233456 271454 233484
rect 271522 233470 271550 236287
rect 271906 233470 271934 239025
rect 272290 233470 272318 239617
rect 272482 239311 272510 246494
rect 272928 246480 273182 246508
rect 273408 246480 273566 246508
rect 273792 246480 274046 246508
rect 273154 241901 273182 246480
rect 273046 241895 273098 241901
rect 273046 241837 273098 241843
rect 273142 241895 273194 241901
rect 273142 241837 273194 241843
rect 273058 241679 273086 241837
rect 272950 241673 273002 241679
rect 272950 241615 273002 241621
rect 273046 241673 273098 241679
rect 273046 241615 273098 241621
rect 272470 239305 272522 239311
rect 272470 239247 272522 239253
rect 272662 236419 272714 236425
rect 272662 236361 272714 236367
rect 272674 233470 272702 236361
rect 272962 234543 272990 241615
rect 273538 239533 273566 246480
rect 274018 241827 274046 246480
rect 273910 241821 273962 241827
rect 273910 241763 273962 241769
rect 274006 241821 274058 241827
rect 274006 241763 274058 241769
rect 273814 241673 273866 241679
rect 273814 241615 273866 241621
rect 273526 239527 273578 239533
rect 273526 239469 273578 239475
rect 273238 239157 273290 239163
rect 273238 239099 273290 239105
rect 272948 234534 273004 234543
rect 272948 234469 273004 234478
rect 273250 233484 273278 239099
rect 273526 237159 273578 237165
rect 273526 237101 273578 237107
rect 273538 233484 273566 237101
rect 273826 235463 273854 241615
rect 273922 235537 273950 241763
rect 274102 241747 274154 241753
rect 274102 241689 274154 241695
rect 274114 236740 274142 241689
rect 274210 237387 274238 246494
rect 274486 242413 274538 242419
rect 274486 242355 274538 242361
rect 274198 237381 274250 237387
rect 274198 237323 274250 237329
rect 274018 236712 274142 236740
rect 273910 235531 273962 235537
rect 273910 235473 273962 235479
rect 273814 235457 273866 235463
rect 273814 235399 273866 235405
rect 274018 233484 274046 236712
rect 274102 236567 274154 236573
rect 274102 236509 274154 236515
rect 273024 233456 273278 233484
rect 273408 233456 273566 233484
rect 273744 233456 274046 233484
rect 274114 233470 274142 236509
rect 274498 233470 274526 242355
rect 274690 236795 274718 246494
rect 275136 246480 275390 246508
rect 275520 246480 275774 246508
rect 276000 246480 276254 246508
rect 274870 239823 274922 239829
rect 274870 239765 274922 239771
rect 274678 236789 274730 236795
rect 274678 236731 274730 236737
rect 274882 233470 274910 239765
rect 275362 239607 275390 246480
rect 275746 240421 275774 246480
rect 275734 240415 275786 240421
rect 275734 240357 275786 240363
rect 275350 239601 275402 239607
rect 275350 239543 275402 239549
rect 275926 239453 275978 239459
rect 275926 239395 275978 239401
rect 275446 239379 275498 239385
rect 275446 239321 275498 239327
rect 275458 233484 275486 239321
rect 275830 237233 275882 237239
rect 275830 237175 275882 237181
rect 275842 233484 275870 237175
rect 275232 233456 275486 233484
rect 275616 233456 275870 233484
rect 275938 233470 275966 239395
rect 276226 239237 276254 246480
rect 276310 239749 276362 239755
rect 276310 239691 276362 239697
rect 276214 239231 276266 239237
rect 276214 239173 276266 239179
rect 276322 233470 276350 239691
rect 276418 236499 276446 246494
rect 276802 240273 276830 246494
rect 276790 240267 276842 240273
rect 276790 240209 276842 240215
rect 277078 239897 277130 239903
rect 277078 239839 277130 239845
rect 276694 237307 276746 237313
rect 276694 237249 276746 237255
rect 276406 236493 276458 236499
rect 276406 236435 276458 236441
rect 276706 233470 276734 237249
rect 277090 233470 277118 239839
rect 277282 237017 277310 246494
rect 277714 246212 277742 246494
rect 278208 246480 278462 246508
rect 278544 246480 278846 246508
rect 277666 246184 277742 246212
rect 277942 246187 277994 246193
rect 277666 240125 277694 246184
rect 277942 246129 277994 246135
rect 277954 245971 277982 246129
rect 277942 245965 277994 245971
rect 277942 245907 277994 245913
rect 277750 245891 277802 245897
rect 277750 245833 277802 245839
rect 277762 245675 277790 245833
rect 277750 245669 277802 245675
rect 277750 245611 277802 245617
rect 278038 244781 278090 244787
rect 278038 244723 278090 244729
rect 277750 244707 277802 244713
rect 277750 244649 277802 244655
rect 277762 242937 277790 244649
rect 277846 244633 277898 244639
rect 277846 244575 277898 244581
rect 277858 243085 277886 244575
rect 277942 244485 277994 244491
rect 277942 244427 277994 244433
rect 277846 243079 277898 243085
rect 277846 243021 277898 243027
rect 277750 242931 277802 242937
rect 277750 242873 277802 242879
rect 277954 242863 277982 244427
rect 277942 242857 277994 242863
rect 277942 242799 277994 242805
rect 278050 242641 278078 244723
rect 278038 242635 278090 242641
rect 278038 242577 278090 242583
rect 277942 241525 277994 241531
rect 277942 241467 277994 241473
rect 277750 241377 277802 241383
rect 277750 241319 277802 241325
rect 277654 240119 277706 240125
rect 277654 240061 277706 240067
rect 277762 240051 277790 241319
rect 277846 241303 277898 241309
rect 277846 241245 277898 241251
rect 277858 240199 277886 241245
rect 277954 240347 277982 241467
rect 277942 240341 277994 240347
rect 277942 240283 277994 240289
rect 278038 240341 278090 240347
rect 278038 240283 278090 240289
rect 277846 240193 277898 240199
rect 277846 240135 277898 240141
rect 277942 240193 277994 240199
rect 277942 240135 277994 240141
rect 277750 240045 277802 240051
rect 277750 239987 277802 239993
rect 277654 239823 277706 239829
rect 277654 239765 277706 239771
rect 277270 237011 277322 237017
rect 277270 236953 277322 236959
rect 277666 233484 277694 239765
rect 277954 239681 277982 240135
rect 278050 239755 278078 240283
rect 278038 239749 278090 239755
rect 278038 239691 278090 239697
rect 278230 239749 278282 239755
rect 278230 239691 278282 239697
rect 277942 239675 277994 239681
rect 277942 239617 277994 239623
rect 278242 236333 278270 239691
rect 278434 236721 278462 246480
rect 278518 239009 278570 239015
rect 278518 238951 278570 238957
rect 278422 236715 278474 236721
rect 278422 236657 278474 236663
rect 278050 236305 278270 236333
rect 278050 233484 278078 236305
rect 278134 236271 278186 236277
rect 278134 236213 278186 236219
rect 277440 233456 277694 233484
rect 277824 233456 278078 233484
rect 278146 233470 278174 236213
rect 278530 233470 278558 238951
rect 278818 236869 278846 246480
rect 278902 239675 278954 239681
rect 278902 239617 278954 239623
rect 278806 236863 278858 236869
rect 278806 236805 278858 236811
rect 278914 233470 278942 239617
rect 279010 233484 279038 246494
rect 279490 240125 279518 246494
rect 279682 246480 279936 246508
rect 280320 246480 280574 246508
rect 279478 240119 279530 240125
rect 279478 240061 279530 240067
rect 279682 239681 279710 246480
rect 279766 243153 279818 243159
rect 279958 243153 280010 243159
rect 279818 243101 279958 243104
rect 279766 243095 280010 243101
rect 279778 243076 279998 243095
rect 280342 239971 280394 239977
rect 280342 239913 280394 239919
rect 279670 239675 279722 239681
rect 279670 239617 279722 239623
rect 279766 237011 279818 237017
rect 279766 236953 279818 236959
rect 279382 236715 279434 236721
rect 279382 236657 279434 236663
rect 279394 233484 279422 236657
rect 279778 233484 279806 236953
rect 279010 233456 279312 233484
rect 279394 233456 279648 233484
rect 279778 233456 280032 233484
rect 280354 233470 280382 239913
rect 280546 239681 280574 246480
rect 280534 239675 280586 239681
rect 280534 239617 280586 239623
rect 280438 239231 280490 239237
rect 280438 239173 280490 239179
rect 280450 233484 280478 239173
rect 280738 239015 280766 246494
rect 280834 246193 280862 246573
rect 287842 246563 287870 246591
rect 287830 246557 287882 246563
rect 280822 246187 280874 246193
rect 280822 246129 280874 246135
rect 281110 239601 281162 239607
rect 281110 239543 281162 239549
rect 280726 239009 280778 239015
rect 280726 238951 280778 238957
rect 280450 233456 280752 233484
rect 281122 233470 281150 239543
rect 281218 236277 281246 246494
rect 281590 239527 281642 239533
rect 281590 239469 281642 239475
rect 281494 237381 281546 237387
rect 281494 237323 281546 237329
rect 281398 236641 281450 236647
rect 281398 236583 281450 236589
rect 281410 236351 281438 236583
rect 281398 236345 281450 236351
rect 281398 236287 281450 236293
rect 281206 236271 281258 236277
rect 281206 236213 281258 236219
rect 281506 233470 281534 237323
rect 281602 233484 281630 239469
rect 281698 237387 281726 246494
rect 281794 246480 282048 246508
rect 282528 246480 282782 246508
rect 281794 239755 281822 246480
rect 282166 243227 282218 243233
rect 282166 243169 282218 243175
rect 281878 241895 281930 241901
rect 281878 241837 281930 241843
rect 281890 239755 281918 241837
rect 281782 239749 281834 239755
rect 281782 239691 281834 239697
rect 281878 239749 281930 239755
rect 281878 239691 281930 239697
rect 281686 237381 281738 237387
rect 281686 237323 281738 237329
rect 282178 233484 282206 243169
rect 282548 242230 282604 242239
rect 282548 242165 282604 242174
rect 282260 240454 282316 240463
rect 282260 240389 282316 240398
rect 282274 237461 282302 240389
rect 282262 237455 282314 237461
rect 282262 237397 282314 237403
rect 281602 233456 281856 233484
rect 282178 233456 282240 233484
rect 282562 233470 282590 242165
rect 282754 237091 282782 246480
rect 282946 239829 282974 246494
rect 283220 242378 283276 242387
rect 283220 242313 283276 242322
rect 283030 240415 283082 240421
rect 283030 240357 283082 240363
rect 283042 239829 283070 240357
rect 282934 239823 282986 239829
rect 282934 239765 282986 239771
rect 283030 239823 283082 239829
rect 283030 239765 283082 239771
rect 282742 237085 282794 237091
rect 282742 237027 282794 237033
rect 283234 233484 283262 242313
rect 283426 241901 283454 246494
rect 283414 241895 283466 241901
rect 283414 241837 283466 241843
rect 283810 239903 283838 246494
rect 284256 246480 284414 246508
rect 284278 242117 284330 242123
rect 284278 242059 284330 242065
rect 283894 240267 283946 240273
rect 283894 240209 283946 240215
rect 283906 239903 283934 240209
rect 283798 239897 283850 239903
rect 283798 239839 283850 239845
rect 283894 239897 283946 239903
rect 283894 239839 283946 239845
rect 283318 234421 283370 234427
rect 283318 234363 283370 234369
rect 282960 233456 283262 233484
rect 283330 233470 283358 234363
rect 283702 234347 283754 234353
rect 283702 234289 283754 234295
rect 283714 233470 283742 234289
rect 284290 233484 284318 242059
rect 284386 236943 284414 246480
rect 284482 246480 284736 246508
rect 284482 237313 284510 246480
rect 284662 242931 284714 242937
rect 284662 242873 284714 242879
rect 284470 237307 284522 237313
rect 284470 237249 284522 237255
rect 284374 236937 284426 236943
rect 284374 236879 284426 236885
rect 284674 233484 284702 242873
rect 284758 242635 284810 242641
rect 284758 242577 284810 242583
rect 284064 233456 284318 233484
rect 284448 233456 284702 233484
rect 284770 233470 284798 242577
rect 285058 239533 285086 246494
rect 285552 246480 285854 246508
rect 285140 242674 285196 242683
rect 285140 242609 285196 242618
rect 285046 239527 285098 239533
rect 285046 239469 285098 239475
rect 285154 233470 285182 242609
rect 285526 239305 285578 239311
rect 285526 239247 285578 239253
rect 285538 233470 285566 239247
rect 285826 236721 285854 246480
rect 286018 239459 286046 246494
rect 286464 246480 286526 246508
rect 286006 239453 286058 239459
rect 286006 239395 286058 239401
rect 286498 237461 286526 246480
rect 286594 246480 286848 246508
rect 287830 246499 287882 246505
rect 287926 246557 287978 246563
rect 287926 246499 287978 246505
rect 286486 237455 286538 237461
rect 286486 237397 286538 237403
rect 286594 237239 286622 246480
rect 287062 241821 287114 241827
rect 287062 241763 287114 241769
rect 286774 240193 286826 240199
rect 286774 240135 286826 240141
rect 286678 239601 286730 239607
rect 286678 239543 286730 239549
rect 286690 239163 286718 239543
rect 286786 239163 286814 240135
rect 286966 239971 287018 239977
rect 286966 239913 287018 239919
rect 286678 239157 286730 239163
rect 286678 239099 286730 239105
rect 286774 239157 286826 239163
rect 286774 239099 286826 239105
rect 286774 237381 286826 237387
rect 286774 237323 286826 237329
rect 286582 237233 286634 237239
rect 286582 237175 286634 237181
rect 285814 236715 285866 236721
rect 285814 236657 285866 236663
rect 286786 234395 286814 237323
rect 286868 236902 286924 236911
rect 286868 236837 286924 236846
rect 286772 234386 286828 234395
rect 286772 234321 286828 234330
rect 286486 233829 286538 233835
rect 286486 233771 286538 233777
rect 286102 233681 286154 233687
rect 286102 233623 286154 233629
rect 286114 233484 286142 233623
rect 286498 233484 286526 233771
rect 286882 233484 286910 236837
rect 285936 233456 286142 233484
rect 286272 233456 286526 233484
rect 286656 233456 286910 233484
rect 286978 233470 287006 239913
rect 287074 239681 287102 241763
rect 287062 239675 287114 239681
rect 287062 239617 287114 239623
rect 287266 239311 287294 246494
rect 287350 246261 287402 246267
rect 287350 246203 287402 246209
rect 287362 243085 287390 246203
rect 287350 243079 287402 243085
rect 287350 243021 287402 243027
rect 287446 242561 287498 242567
rect 287446 242503 287498 242509
rect 287542 242561 287594 242567
rect 287542 242503 287594 242509
rect 287350 241747 287402 241753
rect 287350 241689 287402 241695
rect 287254 239305 287306 239311
rect 287254 239247 287306 239253
rect 287158 237455 287210 237461
rect 287158 237397 287210 237403
rect 287170 237313 287198 237397
rect 287158 237307 287210 237313
rect 287158 237249 287210 237255
rect 287362 233470 287390 241689
rect 287458 233484 287486 242503
rect 287554 242345 287582 242503
rect 287542 242339 287594 242345
rect 287542 242281 287594 242287
rect 287746 239385 287774 246494
rect 287938 246415 287966 246499
rect 288022 246483 288074 246489
rect 288022 246425 288074 246431
rect 287926 246409 287978 246415
rect 287926 246351 287978 246357
rect 288034 246193 288062 246425
rect 288130 246415 288158 246591
rect 288118 246409 288170 246415
rect 288118 246351 288170 246357
rect 288118 246261 288170 246267
rect 288118 246203 288170 246209
rect 287830 246187 287882 246193
rect 287830 246129 287882 246135
rect 288022 246187 288074 246193
rect 288022 246129 288074 246135
rect 287842 244880 287870 246129
rect 288130 245176 288158 246203
rect 287938 245148 288158 245176
rect 287938 245051 287966 245148
rect 287924 245042 287980 245051
rect 288116 245042 288172 245051
rect 287924 244977 287980 244986
rect 288034 245000 288116 245028
rect 288034 244880 288062 245000
rect 288116 244977 288172 244986
rect 287842 244852 288062 244880
rect 288226 240125 288254 246494
rect 288322 246489 288350 246721
rect 288418 246637 288446 246721
rect 290038 246705 290090 246711
rect 290038 246647 290090 246653
rect 288406 246631 288458 246637
rect 288406 246573 288458 246579
rect 288310 246483 288362 246489
rect 288310 246425 288362 246431
rect 288418 246480 288576 246508
rect 289056 246480 289310 246508
rect 288418 240347 288446 246480
rect 288982 242265 289034 242271
rect 288982 242207 289034 242213
rect 288994 241975 289022 242207
rect 288982 241969 289034 241975
rect 288982 241911 289034 241917
rect 289174 241895 289226 241901
rect 289174 241837 289226 241843
rect 289186 241679 289214 241837
rect 289174 241673 289226 241679
rect 289174 241615 289226 241621
rect 288406 240341 288458 240347
rect 288406 240283 288458 240289
rect 289174 240341 289226 240347
rect 289174 240283 289226 240289
rect 288214 240119 288266 240125
rect 288214 240061 288266 240067
rect 289078 240045 289130 240051
rect 289078 239987 289130 239993
rect 287734 239379 287786 239385
rect 287734 239321 287786 239327
rect 287830 239379 287882 239385
rect 287830 239321 287882 239327
rect 288982 239379 289034 239385
rect 288982 239321 289034 239327
rect 287842 239089 287870 239321
rect 288994 239089 289022 239321
rect 287830 239083 287882 239089
rect 287830 239025 287882 239031
rect 288982 239083 289034 239089
rect 288982 239025 289034 239031
rect 288982 237011 289034 237017
rect 288982 236953 289034 236959
rect 288694 236641 288746 236647
rect 288694 236583 288746 236589
rect 288118 236345 288170 236351
rect 288118 236287 288170 236293
rect 287458 233456 287760 233484
rect 288130 233470 288158 236287
rect 288706 233484 288734 236583
rect 288994 236425 289022 236953
rect 288982 236419 289034 236425
rect 288982 236361 289034 236367
rect 289090 233484 289118 239987
rect 288480 233456 288734 233484
rect 288864 233456 289118 233484
rect 289186 233470 289214 240283
rect 289282 237091 289310 246480
rect 289474 242419 289502 246494
rect 289666 246480 289968 246508
rect 289462 242413 289514 242419
rect 289462 242355 289514 242361
rect 289366 241673 289418 241679
rect 289366 241615 289418 241621
rect 289378 239163 289406 241615
rect 289366 239157 289418 239163
rect 289366 239099 289418 239105
rect 289270 237085 289322 237091
rect 289270 237027 289322 237033
rect 289666 236573 289694 246480
rect 290050 245051 290078 246647
rect 290146 246637 290174 246721
rect 290134 246631 290186 246637
rect 290134 246573 290186 246579
rect 290998 246631 291050 246637
rect 290998 246573 291050 246579
rect 290146 246480 290352 246508
rect 290614 246483 290666 246489
rect 290036 245042 290092 245051
rect 290036 244977 290092 244986
rect 290146 244177 290174 246480
rect 290784 246480 290846 246508
rect 290614 246425 290666 246431
rect 290626 246249 290654 246425
rect 290818 246360 290846 246480
rect 291010 246471 291038 246573
rect 290914 246443 291038 246471
rect 290914 246360 290942 246443
rect 290818 246332 290942 246360
rect 291106 246249 291134 246721
rect 291970 246637 291998 246753
rect 292162 246711 292190 246753
rect 311156 246818 311212 246827
rect 307988 246753 308044 246762
rect 309718 246779 309770 246785
rect 292630 246721 292682 246727
rect 292150 246705 292202 246711
rect 292150 246647 292202 246653
rect 291574 246631 291626 246637
rect 291574 246573 291626 246579
rect 291958 246631 292010 246637
rect 291958 246573 292010 246579
rect 291264 246480 291518 246508
rect 290626 246221 290942 246249
rect 290914 246212 290942 246221
rect 291010 246221 291134 246249
rect 291010 246212 291038 246221
rect 290914 246184 291038 246212
rect 290146 244149 290366 244177
rect 289654 236567 289706 236573
rect 289654 236509 289706 236515
rect 289942 236567 289994 236573
rect 289942 236509 289994 236515
rect 289364 236310 289420 236319
rect 289364 236245 289366 236254
rect 289418 236245 289420 236254
rect 289366 236213 289418 236219
rect 289846 233533 289898 233539
rect 289584 233481 289846 233484
rect 289584 233475 289898 233481
rect 289584 233456 289886 233475
rect 289954 233470 289982 236509
rect 290338 236351 290366 244149
rect 290708 242526 290764 242535
rect 290708 242461 290764 242470
rect 290518 241969 290570 241975
rect 290518 241911 290570 241917
rect 290530 241827 290558 241911
rect 290518 241821 290570 241827
rect 290518 241763 290570 241769
rect 290614 241821 290666 241827
rect 290614 241763 290666 241769
rect 290326 236345 290378 236351
rect 290326 236287 290378 236293
rect 290626 233780 290654 241763
rect 290530 233752 290654 233780
rect 290530 233484 290558 233752
rect 290722 233669 290750 242461
rect 290806 242413 290858 242419
rect 290804 242378 290806 242387
rect 290858 242378 290860 242387
rect 290804 242313 290860 242322
rect 290806 239675 290858 239681
rect 290806 239617 290858 239623
rect 290818 236277 290846 239617
rect 291490 239237 291518 246480
rect 291586 241975 291614 246573
rect 292642 246563 292670 246721
rect 297142 246705 297194 246711
rect 296880 246653 297142 246656
rect 296880 246647 297194 246653
rect 304630 246705 304682 246711
rect 304630 246647 304682 246653
rect 296880 246628 297182 246647
rect 292630 246557 292682 246563
rect 297622 246557 297674 246563
rect 292630 246499 292682 246505
rect 291574 241969 291626 241975
rect 291574 241911 291626 241917
rect 291478 239231 291530 239237
rect 291478 239173 291530 239179
rect 290902 239009 290954 239015
rect 290902 238951 290954 238957
rect 290806 236271 290858 236277
rect 290806 236213 290858 236219
rect 290914 236203 290942 238951
rect 291286 237381 291338 237387
rect 291286 237323 291338 237329
rect 290902 236197 290954 236203
rect 290902 236139 290954 236145
rect 290352 233456 290558 233484
rect 290674 233641 290750 233669
rect 290674 233470 290702 233641
rect 291298 233484 291326 237323
rect 291682 237239 291710 246494
rect 291862 239453 291914 239459
rect 291862 239395 291914 239401
rect 291874 239163 291902 239395
rect 292066 239385 292094 246494
rect 292340 245042 292396 245051
rect 292340 244977 292396 244986
rect 292354 244935 292382 244977
rect 292342 244929 292394 244935
rect 292342 244871 292394 244877
rect 292342 242265 292394 242271
rect 292438 242265 292490 242271
rect 292342 242207 292394 242213
rect 292436 242230 292438 242239
rect 292490 242230 292492 242239
rect 292246 242043 292298 242049
rect 292246 241985 292298 241991
rect 292258 239755 292286 241985
rect 292354 241975 292382 242207
rect 292436 242165 292492 242174
rect 292342 241969 292394 241975
rect 292342 241911 292394 241917
rect 292150 239749 292202 239755
rect 292150 239691 292202 239697
rect 292246 239749 292298 239755
rect 292246 239691 292298 239697
rect 292054 239379 292106 239385
rect 292054 239321 292106 239327
rect 291862 239157 291914 239163
rect 291862 239099 291914 239105
rect 291670 237233 291722 237239
rect 291670 237175 291722 237181
rect 291382 237159 291434 237165
rect 291382 237101 291434 237107
rect 291072 233456 291326 233484
rect 291394 233470 291422 237101
rect 291766 236197 291818 236203
rect 291766 236139 291818 236145
rect 291778 233470 291806 236139
rect 292162 233470 292190 239691
rect 292546 239607 292574 246494
rect 292992 246480 293246 246508
rect 292630 240045 292682 240051
rect 292630 239987 292682 239993
rect 292642 239607 292670 239987
rect 292534 239601 292586 239607
rect 292534 239543 292586 239549
rect 292630 239601 292682 239607
rect 292630 239543 292682 239549
rect 293218 239311 293246 246480
rect 293314 246480 293376 246508
rect 293808 246480 294110 246508
rect 293206 239305 293258 239311
rect 293206 239247 293258 239253
rect 293314 239015 293342 246480
rect 293410 242928 294014 242956
rect 293410 242789 293438 242928
rect 293398 242783 293450 242789
rect 293398 242725 293450 242731
rect 293494 242783 293546 242789
rect 293494 242725 293546 242731
rect 293878 242783 293930 242789
rect 293878 242725 293930 242731
rect 293506 242567 293534 242725
rect 293494 242561 293546 242567
rect 293494 242503 293546 242509
rect 293890 242216 293918 242725
rect 293986 242493 294014 242928
rect 293974 242487 294026 242493
rect 293974 242429 294026 242435
rect 293698 242188 293918 242216
rect 293590 242043 293642 242049
rect 293590 241985 293642 241991
rect 293302 239009 293354 239015
rect 293302 238951 293354 238957
rect 292534 237455 292586 237461
rect 292534 237397 292586 237403
rect 292546 233470 292574 237397
rect 293494 233977 293546 233983
rect 293494 233919 293546 233925
rect 292870 233755 292922 233761
rect 292870 233697 292922 233703
rect 292882 233470 292910 233697
rect 293506 233484 293534 233919
rect 293280 233456 293534 233484
rect 293602 233470 293630 241985
rect 293698 237461 293726 242188
rect 294082 239015 294110 246480
rect 294274 240051 294302 246494
rect 294466 246480 294768 246508
rect 295104 246480 295358 246508
rect 294262 240045 294314 240051
rect 294262 239987 294314 239993
rect 294466 239089 294494 246480
rect 295222 239897 295274 239903
rect 295222 239839 295274 239845
rect 294742 239823 294794 239829
rect 294742 239765 294794 239771
rect 294454 239083 294506 239089
rect 294454 239025 294506 239031
rect 294070 239009 294122 239015
rect 294070 238951 294122 238957
rect 293686 237455 293738 237461
rect 293686 237397 293738 237403
rect 293782 237455 293834 237461
rect 293782 237397 293834 237403
rect 293794 236319 293822 237397
rect 294358 236789 294410 236795
rect 294358 236731 294410 236737
rect 293780 236310 293836 236319
rect 293780 236245 293836 236254
rect 293974 236271 294026 236277
rect 293974 236213 294026 236219
rect 293986 233470 294014 236213
rect 294370 233470 294398 236731
rect 294754 233470 294782 239765
rect 294838 236493 294890 236499
rect 294838 236435 294890 236441
rect 294850 233484 294878 236435
rect 295234 233484 295262 239839
rect 295330 236869 295358 246480
rect 295426 246480 295584 246508
rect 295426 237461 295454 246480
rect 295798 240193 295850 240199
rect 295798 240135 295850 240141
rect 295894 240193 295946 240199
rect 295894 240135 295946 240141
rect 295702 239897 295754 239903
rect 295702 239839 295754 239845
rect 295414 237455 295466 237461
rect 295414 237397 295466 237403
rect 295318 236863 295370 236869
rect 295318 236805 295370 236811
rect 295714 233539 295742 239839
rect 295702 233533 295754 233539
rect 294850 233456 295104 233484
rect 295234 233456 295488 233484
rect 295702 233475 295754 233481
rect 295810 233470 295838 240135
rect 295906 236911 295934 240135
rect 296002 239089 296030 246494
rect 296482 241679 296510 246494
rect 297312 246480 297374 246508
rect 297622 246499 297674 246505
rect 297910 246557 297962 246563
rect 300214 246557 300266 246563
rect 297962 246505 298224 246508
rect 297910 246499 298224 246505
rect 296674 243529 297182 243548
rect 296662 243523 297194 243529
rect 296714 243520 297142 243523
rect 296662 243465 296714 243471
rect 297142 243465 297194 243471
rect 296662 243375 296714 243381
rect 297142 243375 297194 243381
rect 296714 243335 297142 243363
rect 296662 243317 296714 243323
rect 297142 243317 297194 243323
rect 296758 243301 296810 243307
rect 296758 243243 296810 243249
rect 297238 243301 297290 243307
rect 297238 243243 297290 243249
rect 296662 243227 296714 243233
rect 296770 243215 296798 243243
rect 296950 243227 297002 243233
rect 296770 243187 296950 243215
rect 296662 243169 296714 243175
rect 296950 243169 297002 243175
rect 296674 243127 296702 243169
rect 296758 243153 296810 243159
rect 296660 243118 296716 243127
rect 297250 243127 297278 243243
rect 296758 243095 296810 243101
rect 297236 243118 297292 243127
rect 296660 243053 296716 243062
rect 296770 242979 296798 243095
rect 297236 243053 297292 243062
rect 296756 242970 296812 242979
rect 296756 242905 296812 242914
rect 296470 241673 296522 241679
rect 296470 241615 296522 241621
rect 296566 240267 296618 240273
rect 296566 240209 296618 240215
rect 295990 239083 296042 239089
rect 295990 239025 296042 239031
rect 295892 236902 295948 236911
rect 295892 236837 295948 236846
rect 296182 236789 296234 236795
rect 296182 236731 296234 236737
rect 296194 233470 296222 236731
rect 296578 233470 296606 240209
rect 296950 239527 297002 239533
rect 296950 239469 297002 239475
rect 296962 233470 296990 239469
rect 297346 236425 297374 246480
rect 297526 242487 297578 242493
rect 297526 242429 297578 242435
rect 297538 242387 297566 242429
rect 297524 242378 297580 242387
rect 297524 242313 297580 242322
rect 297634 242197 297662 246499
rect 297778 246212 297806 246494
rect 297922 246480 298224 246499
rect 297778 246184 297854 246212
rect 297622 242191 297674 242197
rect 297622 242133 297674 242139
rect 297622 239971 297674 239977
rect 297622 239913 297674 239919
rect 297634 239533 297662 239913
rect 297622 239527 297674 239533
rect 297622 239469 297674 239475
rect 297826 239459 297854 246184
rect 297922 244852 298142 244880
rect 297922 244195 297950 244852
rect 298114 244787 298142 244852
rect 298006 244781 298058 244787
rect 298006 244723 298058 244729
rect 298102 244781 298154 244787
rect 298102 244723 298154 244729
rect 298018 244195 298046 244723
rect 297910 244189 297962 244195
rect 297910 244131 297962 244137
rect 298006 244189 298058 244195
rect 298006 244131 298058 244137
rect 298102 242931 298154 242937
rect 298102 242873 298154 242879
rect 297910 242783 297962 242789
rect 297910 242725 297962 242731
rect 297922 242683 297950 242725
rect 297908 242674 297964 242683
rect 297908 242609 297964 242618
rect 297910 242561 297962 242567
rect 297910 242503 297962 242509
rect 297922 242123 297950 242503
rect 298114 242493 298142 242873
rect 298196 242526 298252 242535
rect 298102 242487 298154 242493
rect 298196 242461 298252 242470
rect 298102 242429 298154 242435
rect 298004 242378 298060 242387
rect 298004 242313 298060 242322
rect 298018 242197 298046 242313
rect 298006 242191 298058 242197
rect 298006 242133 298058 242139
rect 298210 242123 298238 242461
rect 297910 242117 297962 242123
rect 297910 242059 297962 242065
rect 298198 242117 298250 242123
rect 298198 242059 298250 242065
rect 298102 241747 298154 241753
rect 298102 241689 298154 241695
rect 298114 240273 298142 241689
rect 298102 240267 298154 240273
rect 298102 240209 298154 240215
rect 298198 239971 298250 239977
rect 298198 239913 298250 239919
rect 297910 239749 297962 239755
rect 298210 239700 298238 239913
rect 297910 239691 297962 239697
rect 297526 239453 297578 239459
rect 297526 239395 297578 239401
rect 297814 239453 297866 239459
rect 297814 239395 297866 239401
rect 297334 236419 297386 236425
rect 297334 236361 297386 236367
rect 297538 236277 297566 239395
rect 297922 237184 297950 239691
rect 298018 239672 298238 239700
rect 298018 239607 298046 239672
rect 298006 239601 298058 239607
rect 298006 239543 298058 239549
rect 297922 237156 298142 237184
rect 298006 237011 298058 237017
rect 298006 236953 298058 236959
rect 297526 236271 297578 236277
rect 297526 236213 297578 236219
rect 297428 234386 297484 234395
rect 297428 234321 297484 234330
rect 297046 233533 297098 233539
rect 297442 233484 297470 234321
rect 297098 233481 297312 233484
rect 297046 233475 297312 233481
rect 297058 233456 297312 233475
rect 297442 233456 297696 233484
rect 298018 233470 298046 236953
rect 298114 233484 298142 237156
rect 298594 233613 298622 246494
rect 299074 239829 299102 246494
rect 299266 246480 299520 246508
rect 300000 246505 300214 246508
rect 302326 246557 302378 246563
rect 300000 246499 300266 246505
rect 300000 246480 300254 246499
rect 300336 246480 300446 246508
rect 299266 242345 299294 246480
rect 299542 244929 299594 244935
rect 299542 244871 299594 244877
rect 299554 243844 299582 244871
rect 299506 243816 299582 243844
rect 299506 243751 299534 243816
rect 299494 243745 299546 243751
rect 299494 243687 299546 243693
rect 300418 243696 300446 246480
rect 300418 243668 300542 243696
rect 300514 242771 300542 243668
rect 300322 242743 300542 242771
rect 299254 242339 299306 242345
rect 299254 242281 299306 242287
rect 299638 242339 299690 242345
rect 299638 242281 299690 242287
rect 299650 242049 299678 242281
rect 299638 242043 299690 242049
rect 299638 241985 299690 241991
rect 299734 241895 299786 241901
rect 299734 241837 299786 241843
rect 299062 239823 299114 239829
rect 299062 239765 299114 239771
rect 299158 239157 299210 239163
rect 299158 239099 299210 239105
rect 298774 236937 298826 236943
rect 298774 236879 298826 236885
rect 298582 233607 298634 233613
rect 298582 233549 298634 233555
rect 298114 233456 298416 233484
rect 298786 233470 298814 236879
rect 299170 233470 299198 239099
rect 299746 237313 299774 241837
rect 299638 237307 299690 237313
rect 299638 237249 299690 237255
rect 299734 237307 299786 237313
rect 299734 237249 299786 237255
rect 299254 236715 299306 236721
rect 299254 236657 299306 236663
rect 299266 233484 299294 236657
rect 299650 233484 299678 237249
rect 300214 236271 300266 236277
rect 300214 236213 300266 236219
rect 299266 233456 299520 233484
rect 299650 233456 299904 233484
rect 300226 233470 300254 236213
rect 300322 234057 300350 242743
rect 300598 240119 300650 240125
rect 300598 240061 300650 240067
rect 300310 234051 300362 234057
rect 300310 233993 300362 233999
rect 300610 233470 300638 240061
rect 300802 237017 300830 246494
rect 301282 242863 301310 246494
rect 301632 246480 301886 246508
rect 301270 242857 301322 242863
rect 301270 242799 301322 242805
rect 301858 239607 301886 246480
rect 301954 246480 302112 246508
rect 302326 246499 302378 246505
rect 301846 239601 301898 239607
rect 301846 239543 301898 239549
rect 301846 239231 301898 239237
rect 301846 239173 301898 239179
rect 300982 237085 301034 237091
rect 300982 237027 301034 237033
rect 300790 237011 300842 237017
rect 300790 236953 300842 236959
rect 300994 233470 301022 237027
rect 301462 236345 301514 236351
rect 301462 236287 301514 236293
rect 301366 233903 301418 233909
rect 301366 233845 301418 233851
rect 301378 233470 301406 233845
rect 301474 233484 301502 236287
rect 301858 233484 301886 239173
rect 301954 234131 301982 246480
rect 302338 237165 302366 246499
rect 302530 239385 302558 246494
rect 303010 239755 303038 246494
rect 302998 239749 303050 239755
rect 302998 239691 303050 239697
rect 302422 239379 302474 239385
rect 302422 239321 302474 239327
rect 302518 239379 302570 239385
rect 302518 239321 302570 239327
rect 302326 237159 302378 237165
rect 302326 237101 302378 237107
rect 301942 234125 301994 234131
rect 301942 234067 301994 234073
rect 301474 233456 301728 233484
rect 301858 233456 302112 233484
rect 302434 233470 302462 239321
rect 302806 239305 302858 239311
rect 302806 239247 302858 239253
rect 302818 233470 302846 239247
rect 303190 239009 303242 239015
rect 303190 238951 303242 238957
rect 303202 233470 303230 238951
rect 303394 234205 303422 246494
rect 303840 246480 304094 246508
rect 303574 240045 303626 240051
rect 303574 239987 303626 239993
rect 303382 234199 303434 234205
rect 303382 234141 303434 234147
rect 303586 233470 303614 239987
rect 304066 239681 304094 246480
rect 304162 246480 304320 246508
rect 304162 243011 304190 246480
rect 304150 243005 304202 243011
rect 304150 242947 304202 242953
rect 304054 239675 304106 239681
rect 304054 239617 304106 239623
rect 304054 239083 304106 239089
rect 304054 239025 304106 239031
rect 303670 236863 303722 236869
rect 303670 236805 303722 236811
rect 303682 233484 303710 236805
rect 304066 233484 304094 239025
rect 303682 233456 303936 233484
rect 304066 233456 304320 233484
rect 304642 233470 304670 246647
rect 308002 246637 308030 246753
rect 309718 246721 309770 246727
rect 309814 246779 309866 246785
rect 309814 246721 309866 246727
rect 310006 246779 310058 246785
rect 327092 246818 327148 246827
rect 311156 246753 311158 246762
rect 310006 246721 310058 246727
rect 311210 246753 311212 246762
rect 326326 246779 326378 246785
rect 311158 246721 311210 246727
rect 327092 246753 327148 246762
rect 327956 246818 328012 246827
rect 327956 246753 328012 246762
rect 328340 246818 328396 246827
rect 328340 246753 328396 246762
rect 328532 246818 328588 246827
rect 348116 246818 348172 246827
rect 340032 246776 340382 246804
rect 328532 246753 328588 246762
rect 326326 246721 326378 246727
rect 307990 246631 308042 246637
rect 307990 246573 308042 246579
rect 309430 246631 309482 246637
rect 309430 246573 309482 246579
rect 307510 246557 307562 246563
rect 304738 240051 304766 246494
rect 304726 240045 304778 240051
rect 304726 239987 304778 239993
rect 305014 239453 305066 239459
rect 305014 239395 305066 239401
rect 304726 237455 304778 237461
rect 304726 237397 304778 237403
rect 304738 236573 304766 237397
rect 304726 236567 304778 236573
rect 304726 236509 304778 236515
rect 305026 233470 305054 239395
rect 305122 234279 305150 246494
rect 305398 242191 305450 242197
rect 305398 242133 305450 242139
rect 305110 234273 305162 234279
rect 305110 234215 305162 234221
rect 305410 233470 305438 242133
rect 305602 241753 305630 246494
rect 305794 246480 306048 246508
rect 306528 246480 306782 246508
rect 305794 242979 305822 246480
rect 305780 242970 305836 242979
rect 305780 242905 305836 242914
rect 306754 241901 306782 246480
rect 306850 246480 306912 246508
rect 308086 246557 308138 246563
rect 307510 246499 307562 246505
rect 306742 241895 306794 241901
rect 306742 241837 306794 241843
rect 305590 241747 305642 241753
rect 305590 241689 305642 241695
rect 305782 239823 305834 239829
rect 305782 239765 305834 239771
rect 305794 233470 305822 239765
rect 306850 239700 306878 246480
rect 306934 240341 306986 240347
rect 306934 240283 306986 240289
rect 306754 239672 306878 239700
rect 305878 237159 305930 237165
rect 305878 237101 305930 237107
rect 305890 233484 305918 237101
rect 306262 237011 306314 237017
rect 306262 236953 306314 236959
rect 306274 233484 306302 236953
rect 306754 234575 306782 239672
rect 306946 239607 306974 240283
rect 306838 239601 306890 239607
rect 306838 239543 306890 239549
rect 306934 239601 306986 239607
rect 306934 239543 306986 239549
rect 306742 234569 306794 234575
rect 306742 234511 306794 234517
rect 305890 233456 306144 233484
rect 306274 233456 306528 233484
rect 306850 233470 306878 239543
rect 307222 239379 307274 239385
rect 307222 239321 307274 239327
rect 307234 233470 307262 239321
rect 307330 234501 307358 246494
rect 307522 246267 307550 246499
rect 307618 246480 307824 246508
rect 308086 246499 308138 246505
rect 307510 246261 307562 246267
rect 307510 246203 307562 246209
rect 307618 241827 307646 246480
rect 308098 246415 308126 246499
rect 308256 246480 308414 246508
rect 308640 246480 308894 246508
rect 308086 246409 308138 246415
rect 308086 246351 308138 246357
rect 308182 246261 308234 246267
rect 307906 246221 308182 246249
rect 307906 246193 307934 246221
rect 308182 246203 308234 246209
rect 307894 246187 307946 246193
rect 307894 246129 307946 246135
rect 307796 245042 307852 245051
rect 307796 244977 307852 244986
rect 307988 245042 308044 245051
rect 308180 245042 308236 245051
rect 308044 245000 308126 245028
rect 307988 244977 308044 244986
rect 307810 244935 307838 244977
rect 307702 244929 307754 244935
rect 307702 244871 307754 244877
rect 307798 244929 307850 244935
rect 307798 244871 307850 244877
rect 307714 243751 307742 244871
rect 308098 244861 308126 245000
rect 308236 245000 308318 245028
rect 308180 244977 308236 244986
rect 308086 244855 308138 244861
rect 308086 244797 308138 244803
rect 308290 244459 308318 245000
rect 308084 244450 308140 244459
rect 308276 244450 308332 244459
rect 308140 244408 308222 244436
rect 308084 244385 308140 244394
rect 307702 243745 307754 243751
rect 307702 243687 307754 243693
rect 308194 243127 308222 244408
rect 308276 244385 308332 244394
rect 308386 243233 308414 246480
rect 308758 244411 308810 244417
rect 308758 244353 308810 244359
rect 308770 243233 308798 244353
rect 308374 243227 308426 243233
rect 308374 243169 308426 243175
rect 308758 243227 308810 243233
rect 308758 243169 308810 243175
rect 308180 243118 308236 243127
rect 308180 243053 308236 243062
rect 307606 241821 307658 241827
rect 307606 241763 307658 241769
rect 308470 241747 308522 241753
rect 308470 241689 308522 241695
rect 308182 240045 308234 240051
rect 308182 239987 308234 239993
rect 307606 239749 307658 239755
rect 307606 239691 307658 239697
rect 307318 234495 307370 234501
rect 307318 234437 307370 234443
rect 307618 233470 307646 239691
rect 307990 239675 308042 239681
rect 307990 239617 308042 239623
rect 308002 233470 308030 239617
rect 308194 233484 308222 239987
rect 308482 233484 308510 241689
rect 308866 239755 308894 246480
rect 308962 246480 309120 246508
rect 308854 239749 308906 239755
rect 308854 239691 308906 239697
rect 308962 238960 308990 246480
rect 309442 245051 309470 246573
rect 309428 245042 309484 245051
rect 309428 244977 309484 244986
rect 309142 244929 309194 244935
rect 309142 244871 309194 244877
rect 309154 244787 309182 244871
rect 309142 244781 309194 244787
rect 309142 244723 309194 244729
rect 309430 243153 309482 243159
rect 309430 243095 309482 243101
rect 309142 241895 309194 241901
rect 309142 241837 309194 241843
rect 308866 238932 308990 238960
rect 308866 234649 308894 238932
rect 308950 238787 309002 238793
rect 308950 238729 309002 238735
rect 308962 236869 308990 238729
rect 308950 236863 309002 236869
rect 308950 236805 309002 236811
rect 308854 234643 308906 234649
rect 308854 234585 308906 234591
rect 309154 233484 309182 241837
rect 308194 233456 308352 233484
rect 308482 233456 308736 233484
rect 309072 233456 309182 233484
rect 309442 233470 309470 243095
rect 309538 239681 309566 246494
rect 309730 246415 309758 246721
rect 309622 246409 309674 246415
rect 309622 246351 309674 246357
rect 309718 246409 309770 246415
rect 309718 246351 309770 246357
rect 309634 244935 309662 246351
rect 309826 246267 309854 246721
rect 309814 246261 309866 246267
rect 309814 246203 309866 246209
rect 309622 244929 309674 244935
rect 309622 244871 309674 244877
rect 309922 244195 309950 246494
rect 310018 246489 310046 246721
rect 324022 246631 324074 246637
rect 324022 246573 324074 246579
rect 310006 246483 310058 246489
rect 310416 246480 310718 246508
rect 310006 246425 310058 246431
rect 309910 244189 309962 244195
rect 309910 244131 309962 244137
rect 309814 241821 309866 241827
rect 309814 241763 309866 241769
rect 309526 239675 309578 239681
rect 309526 239617 309578 239623
rect 309826 233470 309854 241763
rect 310486 241229 310538 241235
rect 310486 241171 310538 241177
rect 310498 240051 310526 241171
rect 310486 240045 310538 240051
rect 310486 239987 310538 239993
rect 310198 239749 310250 239755
rect 310198 239691 310250 239697
rect 310006 237529 310058 237535
rect 310006 237471 310058 237477
rect 310018 237091 310046 237471
rect 310006 237085 310058 237091
rect 310006 237027 310058 237033
rect 310210 233470 310238 239691
rect 310294 239675 310346 239681
rect 310294 239617 310346 239623
rect 310306 233484 310334 239617
rect 310690 233484 310718 246480
rect 310834 246212 310862 246494
rect 310786 246184 310862 246212
rect 311266 246480 311328 246508
rect 310786 236055 310814 246184
rect 310774 236049 310826 236055
rect 310774 235991 310826 235997
rect 310306 233456 310560 233484
rect 310690 233456 310944 233484
rect 311266 233470 311294 246480
rect 311650 240273 311678 246494
rect 311638 240267 311690 240273
rect 311638 240209 311690 240215
rect 311638 239749 311690 239755
rect 311638 239691 311690 239697
rect 311650 233470 311678 239691
rect 312130 236647 312158 246494
rect 312406 244189 312458 244195
rect 312406 244131 312458 244137
rect 312118 236641 312170 236647
rect 312118 236583 312170 236589
rect 312022 234643 312074 234649
rect 312022 234585 312074 234591
rect 312034 233470 312062 234585
rect 312418 233470 312446 244131
rect 312610 239533 312638 246494
rect 312802 246480 313056 246508
rect 313186 246480 313440 246508
rect 312802 239977 312830 246480
rect 313186 240199 313214 246480
rect 313366 240415 313418 240421
rect 313366 240357 313418 240363
rect 313174 240193 313226 240199
rect 313174 240135 313226 240141
rect 312790 239971 312842 239977
rect 312790 239913 312842 239919
rect 312598 239527 312650 239533
rect 312598 239469 312650 239475
rect 312982 236049 313034 236055
rect 312982 235991 313034 235997
rect 312994 233484 313022 235991
rect 313378 233484 313406 240357
rect 313462 240193 313514 240199
rect 313462 240135 313514 240141
rect 312768 233456 313022 233484
rect 313152 233456 313406 233484
rect 313474 233470 313502 240135
rect 313750 239971 313802 239977
rect 313750 239913 313802 239919
rect 313762 233484 313790 239913
rect 313858 239607 313886 246494
rect 314230 241895 314282 241901
rect 314230 241837 314282 241843
rect 314242 241531 314270 241837
rect 314230 241525 314282 241531
rect 314230 241467 314282 241473
rect 314230 240267 314282 240273
rect 314230 240209 314282 240215
rect 313846 239601 313898 239607
rect 313846 239543 313898 239549
rect 313762 233456 313872 233484
rect 314242 233470 314270 240209
rect 314338 233835 314366 246494
rect 314422 241821 314474 241827
rect 314422 241763 314474 241769
rect 314434 241679 314462 241763
rect 314422 241673 314474 241679
rect 314422 241615 314474 241621
rect 314518 241451 314570 241457
rect 314518 241393 314570 241399
rect 314530 241161 314558 241393
rect 314614 241377 314666 241383
rect 314614 241319 314666 241325
rect 314626 241161 314654 241319
rect 314518 241155 314570 241161
rect 314518 241097 314570 241103
rect 314614 241155 314666 241161
rect 314614 241097 314666 241103
rect 314614 240341 314666 240347
rect 314614 240283 314666 240289
rect 314326 233829 314378 233835
rect 314326 233771 314378 233777
rect 314626 233470 314654 240283
rect 314818 239829 314846 246494
rect 315154 246212 315182 246494
rect 315106 246184 315182 246212
rect 315394 246480 315648 246508
rect 314806 239823 314858 239829
rect 314806 239765 314858 239771
rect 315106 233687 315134 246184
rect 315190 241821 315242 241827
rect 315190 241763 315242 241769
rect 315094 233681 315146 233687
rect 315094 233623 315146 233629
rect 315202 233484 315230 241763
rect 315394 237461 315422 246480
rect 316066 241679 316094 246494
rect 316450 242789 316478 246494
rect 316438 242783 316490 242789
rect 316438 242725 316490 242731
rect 316930 242123 316958 246494
rect 317122 246480 317376 246508
rect 317602 246480 317856 246508
rect 317986 246480 318192 246508
rect 318466 246480 318672 246508
rect 317122 242641 317150 246480
rect 317110 242635 317162 242641
rect 317110 242577 317162 242583
rect 316918 242117 316970 242123
rect 316918 242059 316970 242065
rect 316054 241673 316106 241679
rect 316054 241615 316106 241621
rect 316630 241673 316682 241679
rect 316630 241615 316682 241621
rect 315670 239675 315722 239681
rect 315670 239617 315722 239623
rect 315574 237677 315626 237683
rect 315574 237619 315626 237625
rect 315586 237461 315614 237619
rect 315382 237455 315434 237461
rect 315382 237397 315434 237403
rect 315574 237455 315626 237461
rect 315574 237397 315626 237403
rect 315574 237233 315626 237239
rect 315574 237175 315626 237181
rect 315586 233484 315614 237175
rect 314976 233456 315230 233484
rect 315360 233456 315614 233484
rect 315682 233470 315710 239617
rect 316438 239009 316490 239015
rect 316438 238951 316490 238957
rect 315778 238044 316094 238072
rect 315778 237831 315806 238044
rect 315862 237973 315914 237979
rect 315862 237915 315914 237921
rect 315874 237831 315902 237915
rect 316066 237905 316094 238044
rect 316054 237899 316106 237905
rect 316054 237841 316106 237847
rect 315766 237825 315818 237831
rect 315766 237767 315818 237773
rect 315862 237825 315914 237831
rect 315862 237767 315914 237773
rect 316054 234569 316106 234575
rect 316054 234511 316106 234517
rect 316066 233470 316094 234511
rect 316450 233470 316478 238951
rect 316642 237239 316670 241615
rect 316822 240119 316874 240125
rect 316822 240061 316874 240067
rect 316630 237233 316682 237239
rect 316630 237175 316682 237181
rect 316834 233470 316862 240061
rect 317602 237535 317630 246480
rect 317986 242493 318014 246480
rect 318166 244707 318218 244713
rect 318166 244649 318218 244655
rect 318178 243159 318206 244649
rect 318262 244633 318314 244639
rect 318262 244575 318314 244581
rect 318166 243153 318218 243159
rect 318166 243095 318218 243101
rect 318274 243085 318302 244575
rect 318262 243079 318314 243085
rect 318262 243021 318314 243027
rect 317974 242487 318026 242493
rect 317974 242429 318026 242435
rect 317974 242191 318026 242197
rect 317974 242133 318026 242139
rect 317782 241377 317834 241383
rect 317782 241319 317834 241325
rect 317686 238935 317738 238941
rect 317686 238877 317738 238883
rect 317698 238423 317726 238877
rect 317686 238417 317738 238423
rect 317686 238359 317738 238365
rect 317590 237529 317642 237535
rect 317590 237471 317642 237477
rect 317398 237381 317450 237387
rect 317398 237323 317450 237329
rect 317410 233484 317438 237323
rect 317794 233484 317822 241319
rect 317878 241303 317930 241309
rect 317878 241245 317930 241251
rect 317184 233456 317438 233484
rect 317568 233456 317822 233484
rect 317890 233470 317918 241245
rect 317986 238645 318014 242133
rect 318262 239231 318314 239237
rect 318262 239173 318314 239179
rect 318166 238787 318218 238793
rect 318166 238729 318218 238735
rect 317974 238639 318026 238645
rect 317974 238581 318026 238587
rect 318178 238571 318206 238729
rect 318070 238565 318122 238571
rect 318070 238507 318122 238513
rect 318166 238565 318218 238571
rect 318166 238507 318218 238513
rect 318082 238423 318110 238507
rect 318070 238417 318122 238423
rect 318070 238359 318122 238365
rect 318274 233470 318302 239173
rect 318466 237165 318494 246480
rect 319138 242567 319166 246494
rect 319330 246480 319584 246508
rect 319714 246480 319968 246508
rect 319126 242561 319178 242567
rect 319126 242503 319178 242509
rect 318646 238787 318698 238793
rect 318646 238729 318698 238735
rect 318454 237159 318506 237165
rect 318454 237101 318506 237107
rect 318658 233470 318686 238729
rect 319030 237529 319082 237535
rect 319030 237471 319082 237477
rect 319042 233470 319070 237471
rect 319330 236203 319358 246480
rect 319606 242117 319658 242123
rect 319606 242059 319658 242065
rect 319318 236197 319370 236203
rect 319318 236139 319370 236145
rect 319618 233484 319646 242059
rect 319714 234353 319742 246480
rect 320086 238639 320138 238645
rect 320086 238581 320138 238587
rect 319990 236271 320042 236277
rect 319990 236213 320042 236219
rect 319702 234347 319754 234353
rect 319702 234289 319754 234295
rect 320002 233484 320030 236213
rect 319392 233456 319646 233484
rect 319776 233456 320030 233484
rect 320098 233470 320126 238581
rect 320386 234427 320414 246494
rect 320866 242715 320894 246494
rect 320854 242709 320906 242715
rect 320854 242651 320906 242657
rect 321346 242419 321374 246494
rect 321442 246480 321696 246508
rect 321922 246480 322176 246508
rect 321334 242413 321386 242419
rect 321334 242355 321386 242361
rect 320854 239379 320906 239385
rect 320854 239321 320906 239327
rect 320470 236197 320522 236203
rect 320470 236139 320522 236145
rect 320374 234421 320426 234427
rect 320374 234363 320426 234369
rect 320482 233470 320510 236139
rect 320866 233470 320894 239321
rect 321238 239083 321290 239089
rect 321238 239025 321290 239031
rect 321250 233470 321278 239025
rect 321442 233761 321470 246480
rect 321922 242271 321950 246480
rect 321910 242265 321962 242271
rect 321910 242207 321962 242213
rect 321622 239527 321674 239533
rect 321622 239469 321674 239475
rect 321634 236555 321662 239469
rect 321922 238747 322526 238775
rect 321922 238275 321950 238747
rect 322102 238639 322154 238645
rect 322294 238639 322346 238645
rect 322154 238599 322294 238627
rect 322102 238581 322154 238587
rect 322294 238581 322346 238587
rect 322498 238571 322526 238747
rect 322390 238565 322442 238571
rect 322390 238507 322442 238513
rect 322486 238565 322538 238571
rect 322486 238507 322538 238513
rect 322402 238405 322430 238507
rect 322486 238417 322538 238423
rect 322402 238377 322486 238405
rect 322486 238359 322538 238365
rect 321910 238269 321962 238275
rect 321910 238211 321962 238217
rect 321910 238047 321962 238053
rect 321910 237989 321962 237995
rect 322102 238047 322154 238053
rect 322486 238047 322538 238053
rect 322102 237989 322154 237995
rect 322306 238007 322486 238035
rect 321922 237503 321950 237989
rect 322114 237924 322142 237989
rect 322306 237979 322334 238007
rect 322486 237989 322538 237995
rect 322018 237896 322142 237924
rect 322294 237973 322346 237979
rect 322294 237915 322346 237921
rect 322018 237831 322046 237896
rect 322006 237825 322058 237831
rect 322006 237767 322058 237773
rect 322390 237677 322442 237683
rect 322390 237619 322442 237625
rect 321908 237494 321964 237503
rect 322402 237461 322430 237619
rect 321908 237429 321964 237438
rect 322390 237455 322442 237461
rect 322390 237397 322442 237403
rect 322486 237455 322538 237461
rect 322486 237397 322538 237403
rect 322292 237346 322348 237355
rect 322292 237281 322294 237290
rect 322346 237281 322348 237290
rect 322294 237249 322346 237255
rect 322498 237221 322526 237397
rect 322402 237193 322526 237221
rect 321634 236527 321950 236555
rect 321814 236493 321866 236499
rect 321814 236435 321866 236441
rect 321430 233755 321482 233761
rect 321430 233697 321482 233703
rect 321826 233484 321854 236435
rect 321600 233456 321854 233484
rect 321922 233484 321950 236527
rect 322402 234575 322430 237193
rect 322486 237159 322538 237165
rect 322486 237101 322538 237107
rect 322390 234569 322442 234575
rect 322390 234511 322442 234517
rect 322498 233484 322526 237101
rect 322594 233983 322622 246494
rect 323074 243307 323102 246494
rect 323062 243301 323114 243307
rect 323062 243243 323114 243249
rect 323458 242345 323486 246494
rect 323650 246480 323904 246508
rect 323446 242339 323498 242345
rect 323446 242281 323498 242287
rect 323650 239755 323678 246480
rect 324034 246341 324062 246573
rect 326338 246563 326366 246721
rect 326326 246557 326378 246563
rect 324130 246480 324384 246508
rect 324022 246335 324074 246341
rect 324022 246277 324074 246283
rect 323638 239749 323690 239755
rect 323638 239691 323690 239697
rect 323062 239453 323114 239459
rect 323062 239395 323114 239401
rect 322678 239157 322730 239163
rect 322678 239099 322730 239105
rect 322582 233977 322634 233983
rect 322582 233919 322634 233925
rect 321922 233456 321984 233484
rect 322320 233456 322526 233484
rect 322690 233470 322718 239099
rect 322772 237346 322828 237355
rect 322772 237281 322774 237290
rect 322826 237281 322828 237290
rect 322774 237249 322826 237255
rect 323074 233470 323102 239395
rect 323446 239305 323498 239311
rect 323446 239247 323498 239253
rect 323458 233470 323486 239247
rect 324130 237091 324158 246480
rect 324406 239601 324458 239607
rect 324406 239543 324458 239549
rect 324118 237085 324170 237091
rect 324118 237027 324170 237033
rect 324022 236567 324074 236573
rect 324022 236509 324074 236515
rect 324034 233484 324062 236509
rect 324418 233484 324446 239543
rect 324706 239385 324734 246494
rect 325186 241605 325214 246494
rect 325474 246480 325680 246508
rect 325858 246480 326112 246508
rect 326326 246499 326378 246505
rect 326496 246480 326750 246508
rect 325174 241599 325226 241605
rect 325174 241541 325226 241547
rect 325270 241599 325322 241605
rect 325270 241541 325322 241547
rect 325282 239977 325310 241541
rect 325270 239971 325322 239977
rect 325270 239913 325322 239919
rect 324886 239453 324938 239459
rect 324886 239395 324938 239401
rect 324694 239379 324746 239385
rect 324694 239321 324746 239327
rect 324898 239237 324926 239395
rect 324886 239231 324938 239237
rect 324886 239173 324938 239179
rect 325474 239108 325502 246480
rect 325654 239675 325706 239681
rect 325654 239617 325706 239623
rect 325186 239080 325502 239108
rect 324502 236715 324554 236721
rect 324502 236657 324554 236663
rect 323808 233456 324062 233484
rect 324192 233456 324446 233484
rect 324514 233470 324542 236657
rect 325186 233484 325214 239080
rect 325270 236641 325322 236647
rect 325270 236583 325322 236589
rect 324912 233456 325214 233484
rect 325282 233470 325310 236583
rect 325666 233470 325694 239617
rect 325858 238719 325886 246480
rect 326614 239897 326666 239903
rect 326614 239839 326666 239845
rect 325942 238935 325994 238941
rect 325942 238877 325994 238883
rect 325954 238719 325982 238877
rect 325846 238713 325898 238719
rect 325846 238655 325898 238661
rect 325942 238713 325994 238719
rect 325942 238655 325994 238661
rect 326230 236937 326282 236943
rect 326230 236879 326282 236885
rect 326242 233484 326270 236879
rect 326626 233484 326654 239839
rect 326722 238941 326750 246480
rect 326804 245042 326860 245051
rect 326804 244977 326860 244986
rect 326818 244713 326846 244977
rect 326806 244707 326858 244713
rect 326806 244649 326858 244655
rect 326914 241013 326942 246494
rect 327106 246341 327134 246753
rect 327094 246335 327146 246341
rect 327094 246277 327146 246283
rect 327394 241383 327422 246494
rect 327586 246480 327888 246508
rect 327382 241377 327434 241383
rect 327382 241319 327434 241325
rect 326902 241007 326954 241013
rect 326902 240949 326954 240955
rect 326998 241007 327050 241013
rect 326998 240949 327050 240955
rect 327010 240125 327038 240949
rect 326998 240119 327050 240125
rect 326998 240061 327050 240067
rect 327094 239823 327146 239829
rect 327094 239765 327146 239771
rect 326710 238935 326762 238941
rect 326710 238877 326762 238883
rect 326806 238047 326858 238053
rect 326806 237989 326858 237995
rect 326818 237905 326846 237989
rect 326806 237899 326858 237905
rect 326806 237841 326858 237847
rect 326710 237011 326762 237017
rect 326710 236953 326762 236959
rect 326016 233456 326270 233484
rect 326400 233456 326654 233484
rect 326722 233470 326750 236953
rect 327106 233470 327134 239765
rect 327586 238719 327614 246480
rect 327970 244787 327998 246753
rect 328210 246212 328238 246494
rect 328162 246184 328238 246212
rect 327958 244781 328010 244787
rect 327958 244723 328010 244729
rect 328054 244781 328106 244787
rect 328054 244723 328106 244729
rect 328066 244491 328094 244723
rect 328054 244485 328106 244491
rect 328054 244427 328106 244433
rect 328162 241753 328190 246184
rect 328354 245176 328382 246753
rect 328546 246711 328574 246753
rect 328534 246705 328586 246711
rect 328534 246647 328586 246653
rect 329014 246705 329066 246711
rect 329014 246647 329066 246653
rect 339286 246705 339338 246711
rect 339286 246647 339338 246653
rect 328918 246557 328970 246563
rect 328704 246480 328862 246508
rect 328918 246499 328970 246505
rect 328354 245148 328574 245176
rect 328244 245042 328300 245051
rect 328244 244977 328300 244986
rect 328436 245042 328492 245051
rect 328436 244977 328492 244986
rect 328258 244935 328286 244977
rect 328246 244929 328298 244935
rect 328246 244871 328298 244877
rect 328450 244436 328478 244977
rect 328546 244935 328574 245148
rect 328628 245042 328684 245051
rect 328628 244977 328684 244986
rect 328534 244929 328586 244935
rect 328534 244871 328586 244877
rect 328642 244861 328670 244977
rect 328630 244855 328682 244861
rect 328630 244797 328682 244803
rect 328724 244450 328780 244459
rect 328450 244408 328724 244436
rect 328724 244385 328780 244394
rect 328436 243562 328492 243571
rect 328436 243497 328492 243506
rect 328450 242979 328478 243497
rect 328436 242970 328492 242979
rect 328436 242905 328492 242914
rect 328150 241747 328202 241753
rect 328150 241689 328202 241695
rect 328246 241747 328298 241753
rect 328246 241689 328298 241695
rect 328258 241605 328286 241689
rect 328246 241599 328298 241605
rect 328246 241541 328298 241547
rect 327862 239971 327914 239977
rect 327862 239913 327914 239919
rect 327574 238713 327626 238719
rect 327574 238655 327626 238661
rect 327478 237085 327530 237091
rect 327478 237027 327530 237033
rect 327490 233470 327518 237027
rect 327874 233470 327902 239913
rect 328834 239755 328862 246480
rect 328930 246267 328958 246499
rect 328918 246261 328970 246267
rect 328918 246203 328970 246209
rect 329026 244713 329054 246647
rect 329014 244707 329066 244713
rect 329014 244649 329066 244655
rect 328822 239749 328874 239755
rect 328822 239691 328874 239697
rect 328630 239675 328682 239681
rect 328630 239617 328682 239623
rect 328726 239675 328778 239681
rect 328726 239617 328778 239623
rect 328642 239237 328670 239617
rect 328630 239231 328682 239237
rect 328630 239173 328682 239179
rect 328246 236789 328298 236795
rect 328246 236731 328298 236737
rect 328258 233780 328286 236731
rect 328210 233752 328286 233780
rect 328210 233470 328238 233752
rect 328738 233484 328766 239617
rect 328918 238935 328970 238941
rect 328918 238877 328970 238883
rect 328608 233456 328766 233484
rect 328930 233470 328958 238877
rect 329122 238867 329150 246494
rect 329602 241457 329630 246494
rect 329986 241901 330014 246494
rect 330178 246480 330432 246508
rect 330754 246480 330912 246508
rect 329974 241895 330026 241901
rect 329974 241837 330026 241843
rect 329590 241451 329642 241457
rect 329590 241393 329642 241399
rect 330178 241309 330206 246480
rect 330166 241303 330218 241309
rect 330166 241245 330218 241251
rect 329302 240119 329354 240125
rect 329302 240061 329354 240067
rect 329110 238861 329162 238867
rect 329110 238803 329162 238809
rect 329314 233470 329342 240061
rect 330070 239749 330122 239755
rect 330070 239691 330122 239697
rect 329686 237159 329738 237165
rect 329686 237101 329738 237107
rect 329698 233470 329726 237101
rect 330082 233470 330110 239691
rect 330646 238861 330698 238867
rect 330646 238803 330698 238809
rect 330658 233484 330686 238803
rect 330754 238423 330782 246480
rect 331030 241303 331082 241309
rect 331030 241245 331082 241251
rect 330742 238417 330794 238423
rect 330742 238359 330794 238365
rect 331042 233484 331070 241245
rect 331330 239459 331358 246494
rect 331510 241599 331562 241605
rect 331510 241541 331562 241547
rect 331318 239453 331370 239459
rect 331318 239395 331370 239401
rect 331126 238713 331178 238719
rect 331126 238655 331178 238661
rect 330432 233456 330686 233484
rect 330816 233456 331070 233484
rect 331138 233470 331166 238655
rect 331522 233470 331550 241541
rect 331714 241235 331742 246494
rect 331702 241229 331754 241235
rect 331702 241171 331754 241177
rect 331894 238935 331946 238941
rect 331894 238877 331946 238883
rect 331798 238639 331850 238645
rect 331798 238581 331850 238587
rect 331606 238565 331658 238571
rect 331606 238507 331658 238513
rect 331618 238275 331646 238507
rect 331606 238269 331658 238275
rect 331606 238211 331658 238217
rect 331810 236740 331838 238581
rect 331714 236712 331838 236740
rect 331714 236647 331742 236712
rect 331702 236641 331754 236647
rect 331702 236583 331754 236589
rect 331906 233470 331934 238877
rect 332194 238793 332222 246494
rect 332386 246480 332640 246508
rect 332770 246480 333024 246508
rect 332182 238787 332234 238793
rect 332182 238729 332234 238735
rect 332278 238787 332330 238793
rect 332278 238729 332330 238735
rect 332290 238664 332318 238729
rect 332098 238645 332318 238664
rect 332086 238639 332318 238645
rect 332138 238636 332318 238639
rect 332086 238581 332138 238587
rect 332386 237535 332414 246480
rect 332770 241161 332798 246480
rect 333442 242123 333470 246494
rect 333430 242117 333482 242123
rect 333430 242059 333482 242065
rect 333718 241451 333770 241457
rect 333718 241393 333770 241399
rect 332950 241377 333002 241383
rect 332950 241319 333002 241325
rect 333334 241377 333386 241383
rect 333334 241319 333386 241325
rect 332758 241155 332810 241161
rect 332758 241097 332810 241103
rect 332374 237529 332426 237535
rect 332374 237471 332426 237477
rect 332758 237529 332810 237535
rect 332758 237471 332810 237477
rect 332770 236943 332798 237471
rect 332758 236937 332810 236943
rect 332758 236879 332810 236885
rect 332854 236937 332906 236943
rect 332854 236879 332906 236885
rect 332278 236345 332330 236351
rect 332278 236287 332330 236293
rect 332290 233470 332318 236287
rect 332866 233484 332894 236879
rect 332640 233456 332894 233484
rect 332962 233484 332990 241319
rect 332962 233456 333024 233484
rect 333346 233470 333374 241319
rect 333730 233470 333758 241393
rect 333922 236869 333950 246494
rect 334210 246480 334416 246508
rect 334498 246480 334752 246508
rect 334978 246480 335232 246508
rect 334102 238639 334154 238645
rect 334102 238581 334154 238587
rect 333910 236863 333962 236869
rect 333910 236805 333962 236811
rect 334114 233470 334142 238581
rect 334210 236277 334238 246480
rect 334498 240144 334526 246480
rect 334402 240116 334526 240144
rect 334402 240051 334430 240116
rect 334390 240045 334442 240051
rect 334390 239987 334442 239993
rect 334486 240045 334538 240051
rect 334486 239987 334538 239993
rect 334198 236271 334250 236277
rect 334198 236213 334250 236219
rect 334498 233470 334526 239987
rect 334978 238571 335006 246480
rect 335156 243710 335212 243719
rect 335156 243645 335212 243654
rect 334966 238565 335018 238571
rect 334966 238507 335018 238513
rect 335062 236271 335114 236277
rect 335062 236213 335114 236219
rect 335074 233484 335102 236213
rect 334848 233456 335102 233484
rect 335170 233484 335198 243645
rect 335650 242197 335678 246494
rect 335926 244263 335978 244269
rect 335926 244205 335978 244211
rect 335638 242191 335690 242197
rect 335638 242133 335690 242139
rect 335350 238565 335402 238571
rect 335350 238507 335402 238513
rect 335254 238417 335306 238423
rect 335254 238359 335306 238365
rect 335266 236277 335294 238359
rect 335362 237503 335390 238507
rect 335348 237494 335404 237503
rect 335348 237429 335404 237438
rect 335254 236271 335306 236277
rect 335254 236213 335306 236219
rect 335542 235679 335594 235685
rect 335542 235621 335594 235627
rect 335170 233456 335232 233484
rect 335554 233470 335582 235621
rect 335938 233470 335966 244205
rect 336130 236203 336158 246494
rect 336514 241531 336542 246494
rect 336960 246480 337022 246508
rect 336694 244337 336746 244343
rect 336694 244279 336746 244285
rect 336502 241525 336554 241531
rect 336502 241467 336554 241473
rect 336118 236197 336170 236203
rect 336118 236139 336170 236145
rect 336310 235827 336362 235833
rect 336310 235769 336362 235775
rect 336322 233470 336350 235769
rect 336706 233470 336734 244279
rect 336994 238497 337022 246480
rect 337186 246480 337440 246508
rect 337186 239089 337214 246480
rect 337270 243227 337322 243233
rect 337270 243169 337322 243175
rect 337174 239083 337226 239089
rect 337174 239025 337226 239031
rect 336982 238491 337034 238497
rect 336982 238433 337034 238439
rect 336982 235605 337034 235611
rect 336982 235547 337034 235553
rect 336994 233780 337022 235547
rect 336994 233752 337070 233780
rect 337042 233470 337070 233752
rect 337282 233484 337310 243169
rect 337858 241087 337886 246494
rect 338134 244559 338186 244565
rect 338134 244501 338186 244507
rect 337846 241081 337898 241087
rect 337846 241023 337898 241029
rect 337750 235753 337802 235759
rect 337750 235695 337802 235701
rect 337282 233456 337440 233484
rect 337762 233470 337790 235695
rect 338146 233470 338174 244501
rect 338242 236573 338270 246494
rect 338614 244781 338666 244787
rect 338614 244723 338666 244729
rect 338326 241895 338378 241901
rect 338326 241837 338378 241843
rect 338338 241013 338366 241837
rect 338326 241007 338378 241013
rect 338326 240949 338378 240955
rect 338230 236567 338282 236573
rect 338230 236509 338282 236515
rect 338518 235901 338570 235907
rect 338518 235843 338570 235849
rect 338530 233470 338558 235843
rect 338626 233484 338654 244723
rect 338722 238349 338750 246494
rect 338914 246480 339168 246508
rect 338914 239533 338942 246480
rect 339298 246341 339326 246647
rect 339862 246631 339914 246637
rect 339862 246573 339914 246579
rect 340150 246631 340202 246637
rect 340150 246573 340202 246579
rect 339394 246480 339648 246508
rect 339286 246335 339338 246341
rect 339286 246277 339338 246283
rect 339190 241599 339242 241605
rect 339190 241541 339242 241547
rect 339202 239755 339230 241541
rect 339394 240939 339422 246480
rect 339874 246341 339902 246573
rect 339862 246335 339914 246341
rect 339862 246277 339914 246283
rect 339958 246335 340010 246341
rect 339958 246277 340010 246283
rect 339970 246064 339998 246277
rect 340162 246193 340190 246573
rect 340150 246187 340202 246193
rect 340150 246129 340202 246135
rect 340246 246187 340298 246193
rect 340246 246129 340298 246135
rect 339874 246036 339998 246064
rect 339874 245971 339902 246036
rect 340258 245971 340286 246129
rect 339862 245965 339914 245971
rect 339862 245907 339914 245913
rect 340246 245965 340298 245971
rect 340246 245907 340298 245913
rect 339574 243153 339626 243159
rect 340354 243141 340382 246776
rect 348116 246753 348118 246762
rect 348170 246753 348172 246762
rect 348596 246818 348652 246827
rect 367604 246818 367660 246827
rect 348596 246753 348598 246762
rect 348118 246721 348170 246727
rect 348650 246753 348652 246762
rect 348886 246779 348938 246785
rect 348598 246721 348650 246727
rect 348886 246721 348938 246727
rect 350326 246779 350378 246785
rect 367604 246753 367660 246762
rect 367988 246818 368044 246827
rect 367988 246753 368044 246762
rect 369428 246818 369484 246827
rect 369908 246818 369964 246827
rect 369428 246753 369484 246762
rect 369814 246779 369866 246785
rect 350326 246721 350378 246727
rect 339574 243095 339626 243101
rect 340258 243113 340382 243141
rect 339382 240933 339434 240939
rect 339382 240875 339434 240881
rect 339478 240933 339530 240939
rect 339478 240875 339530 240881
rect 339190 239749 339242 239755
rect 339190 239691 339242 239697
rect 338902 239527 338954 239533
rect 338902 239469 338954 239475
rect 338710 238343 338762 238349
rect 338710 238285 338762 238291
rect 339490 236943 339518 240875
rect 339478 236937 339530 236943
rect 339478 236879 339530 236885
rect 338996 235866 339052 235875
rect 338996 235801 339052 235810
rect 339010 233484 339038 235801
rect 339586 233484 339614 243095
rect 339778 241753 339902 241772
rect 339766 241747 339914 241753
rect 339818 241744 339862 241747
rect 339766 241689 339818 241695
rect 339862 241689 339914 241695
rect 340258 239089 340286 243113
rect 340342 243079 340394 243085
rect 340342 243021 340394 243027
rect 339862 239083 339914 239089
rect 339862 239025 339914 239031
rect 340246 239083 340298 239089
rect 340246 239025 340298 239031
rect 339874 237239 339902 239025
rect 339862 237233 339914 237239
rect 339862 237175 339914 237181
rect 339958 236123 340010 236129
rect 339958 236065 340010 236071
rect 338626 233456 338928 233484
rect 339010 233456 339264 233484
rect 339586 233456 339648 233484
rect 339970 233470 339998 236065
rect 340354 233470 340382 243021
rect 340450 238201 340478 246494
rect 340930 239163 340958 246494
rect 341108 243858 341164 243867
rect 341108 243793 341164 243802
rect 340918 239157 340970 239163
rect 340918 239099 340970 239105
rect 340438 238195 340490 238201
rect 340438 238137 340490 238143
rect 340726 235975 340778 235981
rect 340726 235917 340778 235923
rect 340738 233470 340766 235917
rect 341122 233470 341150 243793
rect 341314 239385 341342 246494
rect 341506 246480 341760 246508
rect 341986 246480 342240 246508
rect 341302 239379 341354 239385
rect 341302 239321 341354 239327
rect 341506 238275 341534 246480
rect 341588 244006 341644 244015
rect 341588 243941 341644 243950
rect 341494 238269 341546 238275
rect 341494 238211 341546 238217
rect 341204 235274 341260 235283
rect 341204 235209 341260 235218
rect 341218 233484 341246 235209
rect 341602 233484 341630 243941
rect 341986 239311 342014 246480
rect 342548 243118 342604 243127
rect 342548 243053 342604 243062
rect 341974 239305 342026 239311
rect 341974 239247 342026 239253
rect 342164 235570 342220 235579
rect 342164 235505 342220 235514
rect 341218 233456 341472 233484
rect 341602 233456 341856 233484
rect 342178 233470 342206 235505
rect 342562 233470 342590 243053
rect 342658 240865 342686 246494
rect 342646 240859 342698 240865
rect 342646 240801 342698 240807
rect 343042 236647 343070 246494
rect 343316 244154 343372 244163
rect 343316 244089 343372 244098
rect 343030 236641 343082 236647
rect 343030 236583 343082 236589
rect 342932 235422 342988 235431
rect 342932 235357 342988 235366
rect 342946 233470 342974 235357
rect 343330 233470 343358 244089
rect 343522 238127 343550 246494
rect 343714 246480 343968 246508
rect 344194 246480 344448 246508
rect 343714 239607 343742 246480
rect 343796 244302 343852 244311
rect 343796 244237 343852 244246
rect 343702 239601 343754 239607
rect 343702 239543 343754 239549
rect 343510 238121 343562 238127
rect 343510 238063 343562 238069
rect 343412 235718 343468 235727
rect 343412 235653 343468 235662
rect 343426 233484 343454 235653
rect 343810 233484 343838 244237
rect 344194 240791 344222 246480
rect 344468 244746 344524 244755
rect 344468 244681 344524 244690
rect 344182 240785 344234 240791
rect 344182 240727 344234 240733
rect 344372 235126 344428 235135
rect 344372 235061 344428 235070
rect 343426 233456 343680 233484
rect 343810 233456 344064 233484
rect 344386 233470 344414 235061
rect 344482 233484 344510 244681
rect 344770 236721 344798 246494
rect 345250 238053 345278 246494
rect 345526 243375 345578 243381
rect 345526 243317 345578 243323
rect 345238 238047 345290 238053
rect 345238 237989 345290 237995
rect 344758 236715 344810 236721
rect 344758 236657 344810 236663
rect 345142 234717 345194 234723
rect 345142 234659 345194 234665
rect 344482 233456 344784 233484
rect 345154 233470 345182 234659
rect 345538 233470 345566 243317
rect 345730 240643 345758 246494
rect 345922 246480 346176 246508
rect 346306 246480 346560 246508
rect 345718 240637 345770 240643
rect 345718 240579 345770 240585
rect 345922 238793 345950 246480
rect 346004 243562 346060 243571
rect 346004 243497 346060 243506
rect 345910 238787 345962 238793
rect 345910 238729 345962 238735
rect 345620 236162 345676 236171
rect 345620 236097 345676 236106
rect 345634 233484 345662 236097
rect 346018 233484 346046 243497
rect 346306 237979 346334 246480
rect 346678 243449 346730 243455
rect 346678 243391 346730 243397
rect 346294 237973 346346 237979
rect 346294 237915 346346 237921
rect 346580 236014 346636 236023
rect 346580 235949 346636 235958
rect 345634 233456 345888 233484
rect 346018 233456 346272 233484
rect 346594 233470 346622 235949
rect 346690 233484 346718 243391
rect 346978 239237 347006 246494
rect 347254 246335 347306 246341
rect 347254 246277 347306 246283
rect 347266 245971 347294 246277
rect 347350 246187 347402 246193
rect 347350 246129 347402 246135
rect 347362 246045 347390 246129
rect 347350 246039 347402 246045
rect 347350 245981 347402 245987
rect 347254 245965 347306 245971
rect 347254 245907 347306 245913
rect 347458 240717 347486 246494
rect 347542 246483 347594 246489
rect 347542 246425 347594 246431
rect 347554 246193 347582 246425
rect 347542 246187 347594 246193
rect 347542 246129 347594 246135
rect 347732 243266 347788 243275
rect 347732 243201 347788 243210
rect 347446 240711 347498 240717
rect 347446 240653 347498 240659
rect 346966 239231 347018 239237
rect 346966 239173 347018 239179
rect 347350 234791 347402 234797
rect 347350 234733 347402 234739
rect 346690 233456 346992 233484
rect 347362 233470 347390 234733
rect 347746 233470 347774 243201
rect 347938 237535 347966 246494
rect 348034 246480 348288 246508
rect 348706 246480 348768 246508
rect 348034 238571 348062 246480
rect 348212 245042 348268 245051
rect 348212 244977 348268 244986
rect 348226 244861 348254 244977
rect 348214 244855 348266 244861
rect 348214 244797 348266 244803
rect 348596 244746 348652 244755
rect 348418 244704 348596 244732
rect 348418 244607 348446 244704
rect 348596 244681 348652 244690
rect 348404 244598 348460 244607
rect 348404 244533 348460 244542
rect 348404 242970 348460 242979
rect 348404 242905 348460 242914
rect 348022 238565 348074 238571
rect 348022 238507 348074 238513
rect 347926 237529 347978 237535
rect 347926 237471 347978 237477
rect 347830 235087 347882 235093
rect 347830 235029 347882 235035
rect 347842 233484 347870 235029
rect 348418 233484 348446 242905
rect 348706 239903 348734 246480
rect 348898 245051 348926 246721
rect 350134 246631 350186 246637
rect 350134 246573 350186 246579
rect 348884 245042 348940 245051
rect 348884 244977 348940 244986
rect 348884 242082 348940 242091
rect 348884 242017 348940 242026
rect 348694 239897 348746 239903
rect 348694 239839 348746 239845
rect 348790 234865 348842 234871
rect 348790 234807 348842 234813
rect 347842 233456 348096 233484
rect 348418 233456 348480 233484
rect 348802 233470 348830 234807
rect 348898 233484 348926 242017
rect 349186 240495 349214 246494
rect 349174 240489 349226 240495
rect 349174 240431 349226 240437
rect 349570 237017 349598 246494
rect 349942 243597 349994 243603
rect 349942 243539 349994 243545
rect 349558 237011 349610 237017
rect 349558 236953 349610 236959
rect 349558 235013 349610 235019
rect 349558 234955 349610 234961
rect 348898 233456 349200 233484
rect 349570 233470 349598 234955
rect 349954 233470 349982 243539
rect 350050 239829 350078 246494
rect 350146 246341 350174 246573
rect 350338 246489 350366 246721
rect 352342 246705 352394 246711
rect 352342 246647 352394 246653
rect 350614 246557 350666 246563
rect 350614 246499 350666 246505
rect 350326 246483 350378 246489
rect 350326 246425 350378 246431
rect 350134 246335 350186 246341
rect 350134 246277 350186 246283
rect 350482 246212 350510 246494
rect 350434 246184 350510 246212
rect 350626 246193 350654 246499
rect 350722 246480 350976 246508
rect 350614 246187 350666 246193
rect 350434 240569 350462 246184
rect 350614 246129 350666 246135
rect 350518 241969 350570 241975
rect 350518 241911 350570 241917
rect 350422 240563 350474 240569
rect 350422 240505 350474 240511
rect 350038 239823 350090 239829
rect 350038 239765 350090 239771
rect 350038 235161 350090 235167
rect 350038 235103 350090 235109
rect 350050 233484 350078 235103
rect 350530 233484 350558 241911
rect 350722 237091 350750 246480
rect 351298 237905 351326 246494
rect 351478 243523 351530 243529
rect 351478 243465 351530 243471
rect 351380 239122 351436 239131
rect 351380 239057 351436 239066
rect 351394 238719 351422 239057
rect 351382 238713 351434 238719
rect 351382 238655 351434 238661
rect 351286 237899 351338 237905
rect 351286 237841 351338 237847
rect 350710 237085 350762 237091
rect 350710 237027 350762 237033
rect 350998 235309 351050 235315
rect 350998 235251 351050 235257
rect 350050 233456 350304 233484
rect 350530 233456 350688 233484
rect 351010 233470 351038 235251
rect 351490 233484 351518 243465
rect 351778 239977 351806 246494
rect 352150 243967 352202 243973
rect 352150 243909 352202 243915
rect 351766 239971 351818 239977
rect 351766 239913 351818 239919
rect 351766 234939 351818 234945
rect 351766 234881 351818 234887
rect 351408 233456 351518 233484
rect 351778 233470 351806 234881
rect 352162 233470 352190 243909
rect 352258 240167 352286 246494
rect 352354 246267 352382 246647
rect 352450 246480 352704 246508
rect 353026 246480 353088 246508
rect 352342 246261 352394 246267
rect 352342 246203 352394 246209
rect 352244 240158 352300 240167
rect 352244 240093 352300 240102
rect 352450 236795 352478 246480
rect 352630 243893 352682 243899
rect 352630 243835 352682 243841
rect 352438 236789 352490 236795
rect 352438 236731 352490 236737
rect 352244 234978 352300 234987
rect 352244 234913 352300 234922
rect 352258 233484 352286 234913
rect 352642 233484 352670 243835
rect 353026 237831 353054 246480
rect 353506 239681 353534 246494
rect 353590 243819 353642 243825
rect 353590 243761 353642 243767
rect 353494 239675 353546 239681
rect 353494 239617 353546 239623
rect 353014 237825 353066 237831
rect 353014 237767 353066 237773
rect 353206 235235 353258 235241
rect 353206 235177 353258 235183
rect 352258 233456 352512 233484
rect 352642 233456 352896 233484
rect 353218 233470 353246 235177
rect 353602 233470 353630 243761
rect 353986 240315 354014 246494
rect 354358 243745 354410 243751
rect 354358 243687 354410 243693
rect 353972 240306 354028 240315
rect 353972 240241 354028 240250
rect 353974 235383 354026 235389
rect 353974 235325 354026 235331
rect 353986 233470 354014 235325
rect 354370 233470 354398 243687
rect 354466 237683 354494 246494
rect 354562 246480 354816 246508
rect 355042 246480 355296 246508
rect 354562 240125 354590 246480
rect 354838 243671 354890 243677
rect 354838 243613 354890 243619
rect 354550 240119 354602 240125
rect 354550 240061 354602 240067
rect 354454 237677 354506 237683
rect 354454 237619 354506 237625
rect 354452 234534 354508 234543
rect 354452 234469 354508 234478
rect 354466 233484 354494 234469
rect 354850 233484 354878 243613
rect 355042 241943 355070 246480
rect 355028 241934 355084 241943
rect 355028 241869 355084 241878
rect 355714 237165 355742 246494
rect 355798 244041 355850 244047
rect 355798 243983 355850 243989
rect 355702 237159 355754 237165
rect 355702 237101 355754 237107
rect 355414 235531 355466 235537
rect 355414 235473 355466 235479
rect 354466 233456 354720 233484
rect 354850 233456 355104 233484
rect 355426 233470 355454 235473
rect 355810 233470 355838 243983
rect 356194 237757 356222 246494
rect 356278 244115 356330 244121
rect 356278 244057 356330 244063
rect 356182 237751 356234 237757
rect 356182 237693 356234 237699
rect 356182 235457 356234 235463
rect 356182 235399 356234 235405
rect 356194 233470 356222 235399
rect 356290 233484 356318 244057
rect 356578 241605 356606 246494
rect 356770 246480 357024 246508
rect 357250 246480 357504 246508
rect 356662 245817 356714 245823
rect 356662 245759 356714 245765
rect 356566 241599 356618 241605
rect 356566 241541 356618 241547
rect 356674 233484 356702 245759
rect 356770 241795 356798 246480
rect 357142 245447 357194 245453
rect 357142 245389 357194 245395
rect 356756 241786 356812 241795
rect 356756 241721 356812 241730
rect 357154 233484 357182 245389
rect 357250 238867 357278 246480
rect 357622 245521 357674 245527
rect 357622 245463 357674 245469
rect 357238 238861 357290 238867
rect 357238 238803 357290 238809
rect 356290 233456 356592 233484
rect 356674 233456 356928 233484
rect 357154 233456 357312 233484
rect 357634 233470 357662 245463
rect 357826 237609 357854 246494
rect 358006 245743 358058 245749
rect 358006 245685 358058 245691
rect 357814 237603 357866 237609
rect 357814 237545 357866 237551
rect 358018 233470 358046 245685
rect 358306 241309 358334 246494
rect 358486 245003 358538 245009
rect 358486 244945 358538 244951
rect 358294 241303 358346 241309
rect 358294 241245 358346 241251
rect 358390 237307 358442 237313
rect 358390 237249 358442 237255
rect 358402 233470 358430 237249
rect 358498 233484 358526 244945
rect 358786 238793 358814 246494
rect 358978 246480 359232 246508
rect 359362 246480 359616 246508
rect 358978 238983 359006 246480
rect 359362 241531 359390 246480
rect 359350 241525 359402 241531
rect 359350 241467 359402 241473
rect 360034 241351 360062 246494
rect 360118 241969 360170 241975
rect 360118 241911 360170 241917
rect 360130 241753 360158 241911
rect 360118 241747 360170 241753
rect 360118 241689 360170 241695
rect 360020 241342 360076 241351
rect 360020 241277 360076 241286
rect 360214 239971 360266 239977
rect 360214 239913 360266 239919
rect 358964 238974 359020 238983
rect 358964 238909 359020 238918
rect 358774 238787 358826 238793
rect 358774 238729 358826 238735
rect 358870 238713 358922 238719
rect 358870 238655 358922 238661
rect 358882 233484 358910 238655
rect 359830 237825 359882 237831
rect 359830 237767 359882 237773
rect 359252 236606 359308 236615
rect 359252 236541 359308 236550
rect 359266 233484 359294 236541
rect 358498 233456 358800 233484
rect 358882 233456 359136 233484
rect 359266 233456 359520 233484
rect 359842 233470 359870 237767
rect 360226 233470 360254 239913
rect 360514 238941 360542 246494
rect 360706 246480 361008 246508
rect 361090 246480 361344 246508
rect 361570 246480 361824 246508
rect 360598 240119 360650 240125
rect 360598 240061 360650 240067
rect 360502 238935 360554 238941
rect 360502 238877 360554 238883
rect 360610 233470 360638 240061
rect 360706 238835 360734 246480
rect 360982 241525 361034 241531
rect 360982 241467 361034 241473
rect 360692 238826 360748 238835
rect 360692 238761 360748 238770
rect 360994 233470 361022 241467
rect 361090 236351 361118 246480
rect 361570 241203 361598 246480
rect 361942 241599 361994 241605
rect 361942 241541 361994 241547
rect 361556 241194 361612 241203
rect 361556 241129 361612 241138
rect 361558 239453 361610 239459
rect 361558 239395 361610 239401
rect 361078 236345 361130 236351
rect 361078 236287 361130 236293
rect 361570 233484 361598 239395
rect 361954 233484 361982 241541
rect 362038 241303 362090 241309
rect 362038 241245 362090 241251
rect 361344 233456 361598 233484
rect 361728 233456 361982 233484
rect 362050 233470 362078 241245
rect 362242 240939 362270 246494
rect 362422 241007 362474 241013
rect 362422 240949 362474 240955
rect 362230 240933 362282 240939
rect 362230 240875 362282 240881
rect 362434 233470 362462 240949
rect 362722 238687 362750 246494
rect 362902 241451 362954 241457
rect 362902 241393 362954 241399
rect 362914 241087 362942 241393
rect 362902 241081 362954 241087
rect 363106 241055 363134 246494
rect 363298 246480 363552 246508
rect 363874 246480 364032 246508
rect 363190 241451 363242 241457
rect 363190 241393 363242 241399
rect 362902 241023 362954 241029
rect 363092 241046 363148 241055
rect 363092 240981 363148 240990
rect 362708 238678 362764 238687
rect 362708 238613 362764 238622
rect 362806 237899 362858 237905
rect 362806 237841 362858 237847
rect 362818 233470 362846 237841
rect 363202 233470 363230 241393
rect 363298 241383 363326 246480
rect 363286 241377 363338 241383
rect 363286 241319 363338 241325
rect 363766 241229 363818 241235
rect 363766 241171 363818 241177
rect 363778 233484 363806 241171
rect 363874 238391 363902 246480
rect 364150 241377 364202 241383
rect 364150 241319 364202 241325
rect 363860 238382 363916 238391
rect 363860 238317 363916 238326
rect 364162 233484 364190 241319
rect 364246 241155 364298 241161
rect 364246 241097 364298 241103
rect 363552 233456 363806 233484
rect 363936 233456 364190 233484
rect 364258 233470 364286 241097
rect 364354 241087 364382 246494
rect 364342 241081 364394 241087
rect 364342 241023 364394 241029
rect 364834 240759 364862 246494
rect 365014 240785 365066 240791
rect 364820 240750 364876 240759
rect 365014 240727 365066 240733
rect 364820 240685 364876 240694
rect 364630 240637 364682 240643
rect 364630 240579 364682 240585
rect 364642 233470 364670 240579
rect 365026 233470 365054 240727
rect 365314 238645 365342 246494
rect 365760 246480 365822 246508
rect 365398 240563 365450 240569
rect 365398 240505 365450 240511
rect 365302 238639 365354 238645
rect 365302 238581 365354 238587
rect 365410 233470 365438 240505
rect 365794 238243 365822 246480
rect 365890 246480 366144 246508
rect 365890 240051 365918 246480
rect 365974 240933 366026 240939
rect 365974 240875 366026 240881
rect 365878 240045 365930 240051
rect 365878 239987 365930 239993
rect 365780 238234 365836 238243
rect 365780 238169 365836 238178
rect 365986 233484 366014 240875
rect 366358 240859 366410 240865
rect 366358 240801 366410 240807
rect 366370 233484 366398 240801
rect 366562 240611 366590 246494
rect 366548 240602 366604 240611
rect 366548 240537 366604 240546
rect 366454 240489 366506 240495
rect 366454 240431 366506 240437
rect 365760 233456 366014 233484
rect 366144 233456 366398 233484
rect 366466 233470 366494 240431
rect 366838 238935 366890 238941
rect 366838 238877 366890 238883
rect 366850 233470 366878 238877
rect 367042 238423 367070 246494
rect 367522 245897 367550 246494
rect 367618 246341 367646 246753
rect 367714 246480 367872 246508
rect 367606 246335 367658 246341
rect 367606 246277 367658 246283
rect 367510 245891 367562 245897
rect 367510 245833 367562 245839
rect 367222 240711 367274 240717
rect 367222 240653 367274 240659
rect 367030 238417 367082 238423
rect 367030 238359 367082 238365
rect 367234 233470 367262 240653
rect 367604 240602 367660 240611
rect 367604 240537 367660 240546
rect 367618 233470 367646 240537
rect 367714 234649 367742 246480
rect 368002 246193 368030 246753
rect 368470 246631 368522 246637
rect 368470 246573 368522 246579
rect 369046 246631 369098 246637
rect 369046 246573 369098 246579
rect 368098 246480 368352 246508
rect 367990 246187 368042 246193
rect 367990 246129 368042 246135
rect 368098 245971 368126 246480
rect 368374 246409 368426 246415
rect 368374 246351 368426 246357
rect 368386 245971 368414 246351
rect 368086 245965 368138 245971
rect 368086 245907 368138 245913
rect 368374 245965 368426 245971
rect 368374 245907 368426 245913
rect 368482 245620 368510 246573
rect 368566 245817 368618 245823
rect 368566 245759 368618 245765
rect 368386 245592 368510 245620
rect 368386 245051 368414 245592
rect 368372 245042 368428 245051
rect 368372 244977 368428 244986
rect 368470 244929 368522 244935
rect 368470 244871 368522 244877
rect 368482 244607 368510 244871
rect 368468 244598 368524 244607
rect 368468 244533 368524 244542
rect 368578 244459 368606 245759
rect 368564 244450 368620 244459
rect 368564 244385 368620 244394
rect 368770 244195 368798 246494
rect 369058 245051 369086 246573
rect 369442 246563 369470 246753
rect 369908 246753 369910 246762
rect 369814 246721 369866 246727
rect 369962 246753 369964 246762
rect 370196 246818 370252 246827
rect 370196 246753 370252 246762
rect 370676 246818 370732 246827
rect 370676 246753 370732 246762
rect 377204 246818 377260 246827
rect 388244 246818 388300 246827
rect 377204 246753 377260 246762
rect 378646 246779 378698 246785
rect 369910 246721 369962 246727
rect 369826 246637 369854 246721
rect 369814 246631 369866 246637
rect 369814 246573 369866 246579
rect 369430 246557 369482 246563
rect 369430 246499 369482 246505
rect 369718 246557 369770 246563
rect 369718 246499 369770 246505
rect 369250 245675 369278 246494
rect 369238 245669 369290 245675
rect 369238 245611 369290 245617
rect 369044 245042 369100 245051
rect 369044 244977 369100 244986
rect 368854 244855 368906 244861
rect 368854 244797 368906 244803
rect 368866 244607 368894 244797
rect 369140 244746 369196 244755
rect 369140 244681 369196 244690
rect 368852 244598 368908 244607
rect 368852 244533 368908 244542
rect 368758 244189 368810 244195
rect 369154 244163 369182 244681
rect 368758 244131 368810 244137
rect 369140 244154 369196 244163
rect 369140 244089 369196 244098
rect 368182 238861 368234 238867
rect 368182 238803 368234 238809
rect 367702 234643 367754 234649
rect 367702 234585 367754 234591
rect 368194 233484 368222 238803
rect 368566 238787 368618 238793
rect 368566 238729 368618 238735
rect 368578 237387 368606 238729
rect 368662 238639 368714 238645
rect 368662 238581 368714 238587
rect 368566 237381 368618 237387
rect 368566 237323 368618 237329
rect 368566 234495 368618 234501
rect 368566 234437 368618 234443
rect 368578 233484 368606 234437
rect 367968 233456 368222 233484
rect 368352 233456 368606 233484
rect 368674 233470 368702 238581
rect 369430 238491 369482 238497
rect 369430 238433 369482 238439
rect 369046 237307 369098 237313
rect 369046 237249 369098 237255
rect 369058 233470 369086 237249
rect 369442 233470 369470 238433
rect 369634 236055 369662 246494
rect 369730 245971 369758 246499
rect 369826 246480 370080 246508
rect 369718 245965 369770 245971
rect 369718 245907 369770 245913
rect 369826 245601 369854 246480
rect 370210 246193 370238 246753
rect 370690 246637 370718 246753
rect 377218 246711 377246 246753
rect 392564 246818 392620 246827
rect 388244 246753 388300 246762
rect 389494 246779 389546 246785
rect 378646 246721 378698 246727
rect 377206 246705 377258 246711
rect 377206 246647 377258 246653
rect 370678 246631 370730 246637
rect 370678 246573 370730 246579
rect 370306 246480 370560 246508
rect 370198 246187 370250 246193
rect 370198 246129 370250 246135
rect 369814 245595 369866 245601
rect 369814 245537 369866 245543
rect 370306 240421 370334 246480
rect 370294 240415 370346 240421
rect 370294 240357 370346 240363
rect 370978 240019 371006 246494
rect 371362 240199 371390 246494
rect 371842 241975 371870 246494
rect 372034 246480 372288 246508
rect 372418 246480 372672 246508
rect 372898 246480 373152 246508
rect 373282 246480 373584 246508
rect 372034 245379 372062 246480
rect 372022 245373 372074 245379
rect 372022 245315 372074 245321
rect 371830 241969 371882 241975
rect 371830 241911 371882 241917
rect 372418 240273 372446 246480
rect 372898 245231 372926 246480
rect 372886 245225 372938 245231
rect 372886 245167 372938 245173
rect 373282 240347 373310 246480
rect 374050 245305 374078 246494
rect 374038 245299 374090 245305
rect 374038 245241 374090 245247
rect 374434 241827 374462 246494
rect 374626 246480 374880 246508
rect 375106 246480 375360 246508
rect 374626 245083 374654 246480
rect 374614 245077 374666 245083
rect 374614 245019 374666 245025
rect 374422 241821 374474 241827
rect 374422 241763 374474 241769
rect 375106 241679 375134 246480
rect 375778 245157 375806 246494
rect 375766 245151 375818 245157
rect 375766 245093 375818 245099
rect 375094 241673 375146 241679
rect 376162 241647 376190 246494
rect 375094 241615 375146 241621
rect 376148 241638 376204 241647
rect 373942 241599 373994 241605
rect 376148 241573 376204 241582
rect 373942 241541 373994 241547
rect 373954 241309 373982 241541
rect 373558 241303 373610 241309
rect 373558 241245 373610 241251
rect 373942 241303 373994 241309
rect 373942 241245 373994 241251
rect 373570 241087 373598 241245
rect 373558 241081 373610 241087
rect 373558 241023 373610 241029
rect 373270 240341 373322 240347
rect 373270 240283 373322 240289
rect 372406 240267 372458 240273
rect 372406 240209 372458 240215
rect 376438 240267 376490 240273
rect 376438 240209 376490 240215
rect 371350 240193 371402 240199
rect 371350 240135 371402 240141
rect 373078 240193 373130 240199
rect 373078 240135 373130 240141
rect 370964 240010 371020 240019
rect 370964 239945 371020 239954
rect 372598 238713 372650 238719
rect 372598 238655 372650 238661
rect 371638 238417 371690 238423
rect 371638 238359 371690 238365
rect 370390 238343 370442 238349
rect 370390 238285 370442 238291
rect 369814 238269 369866 238275
rect 369814 238211 369866 238217
rect 369622 236049 369674 236055
rect 369622 235991 369674 235997
rect 369826 233470 369854 238211
rect 370402 233484 370430 238285
rect 370870 238195 370922 238201
rect 370870 238137 370922 238143
rect 370774 236863 370826 236869
rect 370774 236805 370826 236811
rect 370786 233484 370814 236805
rect 370176 233456 370430 233484
rect 370560 233456 370814 233484
rect 370882 233470 370910 238137
rect 371254 238047 371306 238053
rect 371254 237989 371306 237995
rect 371266 233470 371294 237989
rect 371650 233470 371678 238359
rect 372022 238121 372074 238127
rect 372022 238063 372074 238069
rect 372034 233470 372062 238063
rect 372610 233484 372638 238655
rect 372982 237455 373034 237461
rect 372982 237397 373034 237403
rect 372994 233484 373022 237397
rect 372384 233456 372638 233484
rect 372768 233456 373022 233484
rect 373090 233470 373118 240135
rect 375670 239897 375722 239903
rect 375670 239839 375722 239845
rect 374806 239675 374858 239681
rect 374806 239617 374858 239623
rect 373846 239601 373898 239607
rect 373846 239543 373898 239549
rect 373462 237529 373514 237535
rect 373462 237471 373514 237477
rect 373474 233470 373502 237471
rect 373858 233470 373886 239543
rect 374230 237603 374282 237609
rect 374230 237545 374282 237551
rect 374242 233470 374270 237545
rect 374818 233484 374846 239617
rect 375190 239083 375242 239089
rect 375190 239025 375242 239031
rect 375202 233484 375230 239025
rect 375286 237973 375338 237979
rect 375286 237915 375338 237921
rect 374592 233456 374846 233484
rect 374976 233456 375230 233484
rect 375298 233470 375326 237915
rect 375682 233470 375710 239839
rect 376054 239749 376106 239755
rect 376054 239691 376106 239697
rect 375958 238861 376010 238867
rect 375958 238803 376010 238809
rect 375970 238571 375998 238803
rect 375958 238565 376010 238571
rect 375958 238507 376010 238513
rect 376066 233470 376094 239691
rect 376450 233470 376478 240209
rect 376642 237387 376670 246494
rect 376834 246480 377088 246508
rect 377314 246480 377568 246508
rect 377698 246480 377904 246508
rect 376834 241499 376862 246480
rect 377014 241747 377066 241753
rect 377014 241689 377066 241695
rect 376820 241490 376876 241499
rect 376820 241425 376876 241434
rect 376630 237381 376682 237387
rect 376630 237323 376682 237329
rect 377026 233484 377054 241689
rect 377206 240045 377258 240051
rect 377206 239987 377258 239993
rect 377218 233780 377246 239987
rect 377314 239015 377342 246480
rect 377494 239157 377546 239163
rect 377494 239099 377546 239105
rect 377302 239009 377354 239015
rect 377302 238951 377354 238957
rect 376800 233456 377054 233484
rect 377170 233752 377246 233780
rect 377170 233470 377198 233752
rect 377506 233470 377534 239099
rect 377698 238539 377726 246480
rect 378370 241901 378398 246494
rect 378658 246415 378686 246721
rect 388258 246711 388286 246753
rect 392564 246753 392620 246762
rect 392948 246818 393004 246827
rect 393428 246818 393484 246827
rect 392948 246753 393004 246762
rect 393046 246779 393098 246785
rect 389494 246721 389546 246727
rect 388246 246705 388298 246711
rect 383184 246628 383486 246656
rect 388246 246647 388298 246653
rect 389014 246705 389066 246711
rect 389014 246647 389066 246653
rect 378646 246409 378698 246415
rect 378646 246351 378698 246357
rect 378358 241895 378410 241901
rect 378358 241837 378410 241843
rect 378850 240907 378878 246494
rect 379042 246480 379296 246508
rect 379426 246480 379680 246508
rect 378836 240898 378892 240907
rect 378836 240833 378892 240842
rect 378262 240415 378314 240421
rect 378262 240357 378314 240363
rect 377878 240341 377930 240347
rect 377878 240283 377930 240289
rect 377684 238530 377740 238539
rect 377684 238465 377740 238474
rect 377890 233470 377918 240283
rect 378274 233470 378302 240357
rect 378742 240119 378794 240125
rect 378742 240061 378794 240067
rect 378646 239971 378698 239977
rect 378646 239913 378698 239919
rect 378658 239459 378686 239913
rect 378646 239453 378698 239459
rect 378646 239395 378698 239401
rect 378754 239311 378782 240061
rect 378742 239305 378794 239311
rect 378742 239247 378794 239253
rect 378646 239231 378698 239237
rect 378646 239173 378698 239179
rect 378658 233470 378686 239173
rect 379042 238793 379070 246480
rect 379222 241821 379274 241827
rect 379222 241763 379274 241769
rect 379030 238787 379082 238793
rect 379030 238729 379082 238735
rect 379234 233484 379262 241763
rect 379426 234839 379454 246480
rect 379606 241673 379658 241679
rect 379606 241615 379658 241621
rect 379412 234830 379468 234839
rect 379412 234765 379468 234774
rect 379618 233484 379646 241615
rect 380098 241531 380126 246494
rect 380086 241525 380138 241531
rect 380086 241467 380138 241473
rect 380578 239829 380606 246494
rect 380854 239897 380906 239903
rect 380854 239839 380906 239845
rect 380566 239823 380618 239829
rect 380566 239765 380618 239771
rect 380086 239379 380138 239385
rect 380086 239321 380138 239327
rect 379702 238787 379754 238793
rect 379702 238729 379754 238735
rect 379008 233456 379262 233484
rect 379392 233456 379646 233484
rect 379714 233470 379742 238729
rect 379990 237159 380042 237165
rect 379990 237101 380042 237107
rect 380002 234501 380030 237101
rect 379990 234495 380042 234501
rect 379990 234437 380042 234443
rect 380098 233470 380126 239321
rect 380470 239009 380522 239015
rect 380470 238951 380522 238957
rect 380182 237307 380234 237313
rect 380182 237249 380234 237255
rect 380194 237165 380222 237249
rect 380182 237159 380234 237165
rect 380182 237101 380234 237107
rect 380482 233470 380510 238951
rect 380866 233470 380894 239839
rect 380962 237831 380990 246494
rect 381154 246480 381408 246508
rect 381888 246480 382142 246508
rect 380950 237825 381002 237831
rect 380950 237767 381002 237773
rect 381154 236869 381182 246480
rect 381814 240119 381866 240125
rect 381814 240061 381866 240067
rect 381430 238935 381482 238941
rect 381430 238877 381482 238883
rect 381142 236863 381194 236869
rect 381142 236805 381194 236811
rect 381442 233484 381470 238877
rect 381826 233484 381854 240061
rect 381910 236715 381962 236721
rect 381910 236657 381962 236663
rect 381216 233456 381470 233484
rect 381600 233456 381854 233484
rect 381922 233470 381950 236657
rect 382114 233484 382142 246480
rect 382306 237905 382334 246494
rect 382690 239681 382718 246494
rect 383350 246409 383402 246415
rect 383350 246351 383402 246357
rect 383062 246187 383114 246193
rect 383062 246129 383114 246135
rect 383158 246187 383210 246193
rect 383158 246129 383210 246135
rect 383074 245749 383102 246129
rect 383170 245897 383198 246129
rect 383158 245891 383210 245897
rect 383158 245833 383210 245839
rect 383062 245743 383114 245749
rect 383062 245685 383114 245691
rect 383062 244263 383114 244269
rect 383062 244205 383114 244211
rect 383074 241795 383102 244205
rect 383060 241786 383116 241795
rect 383060 241721 383116 241730
rect 383060 240158 383116 240167
rect 383060 240093 383062 240102
rect 383114 240093 383116 240102
rect 383062 240061 383114 240067
rect 383060 240010 383116 240019
rect 383060 239945 383062 239954
rect 383114 239945 383116 239954
rect 383062 239913 383114 239919
rect 382678 239675 382730 239681
rect 382678 239617 382730 239623
rect 383254 239675 383306 239681
rect 383254 239617 383306 239623
rect 383062 239527 383114 239533
rect 383266 239515 383294 239617
rect 383114 239487 383294 239515
rect 383062 239469 383114 239475
rect 383060 239122 383116 239131
rect 382882 239080 383060 239108
rect 382294 237899 382346 237905
rect 382294 237841 382346 237847
rect 382882 233484 382910 239080
rect 383060 239057 383116 239066
rect 383362 238867 383390 246351
rect 383458 244269 383486 246628
rect 388534 246631 388586 246637
rect 388534 246573 388586 246579
rect 383602 246415 383630 246494
rect 383842 246480 384096 246508
rect 383590 246409 383642 246415
rect 383590 246351 383642 246357
rect 383446 244263 383498 244269
rect 383446 244205 383498 244211
rect 383554 241596 383774 241624
rect 383554 241531 383582 241596
rect 383542 241525 383594 241531
rect 383542 241467 383594 241473
rect 383638 241525 383690 241531
rect 383638 241467 383690 241473
rect 383350 238861 383402 238867
rect 383350 238803 383402 238809
rect 383062 238713 383114 238719
rect 383060 238678 383062 238687
rect 383114 238678 383116 238687
rect 383060 238613 383116 238622
rect 383062 234347 383114 234353
rect 383062 234289 383114 234295
rect 382114 233456 382320 233484
rect 382704 233456 382910 233484
rect 383074 233470 383102 234289
rect 383650 233484 383678 241467
rect 383424 233456 383678 233484
rect 383746 233484 383774 241596
rect 383842 239237 383870 246480
rect 383830 239231 383882 239237
rect 383830 239173 383882 239179
rect 384118 237899 384170 237905
rect 384118 237841 384170 237847
rect 383746 233456 383808 233484
rect 384130 233470 384158 237841
rect 384418 234353 384446 246494
rect 384610 246480 384912 246508
rect 384610 238571 384638 246480
rect 385268 243414 385324 243423
rect 385268 243349 385324 243358
rect 384886 239823 384938 239829
rect 384886 239765 384938 239771
rect 384598 238565 384650 238571
rect 384598 238507 384650 238513
rect 384502 237825 384554 237831
rect 384502 237767 384554 237773
rect 384406 234347 384458 234353
rect 384406 234289 384458 234295
rect 384514 233470 384542 237767
rect 384898 233470 384926 239765
rect 385282 233470 385310 243349
rect 385378 238793 385406 246494
rect 385570 246480 385824 246508
rect 385954 246480 386208 246508
rect 385570 241531 385598 246480
rect 385558 241525 385610 241531
rect 385558 241467 385610 241473
rect 385366 238787 385418 238793
rect 385366 238729 385418 238735
rect 385954 237313 385982 246480
rect 386626 239385 386654 246494
rect 386998 240267 387050 240273
rect 386998 240209 387050 240215
rect 386806 240193 386858 240199
rect 386806 240135 386858 240141
rect 386614 239379 386666 239385
rect 386614 239321 386666 239327
rect 386710 239379 386762 239385
rect 386710 239321 386762 239327
rect 386722 239163 386750 239321
rect 386818 239237 386846 240135
rect 387010 239755 387038 240209
rect 386998 239749 387050 239755
rect 386998 239691 387050 239697
rect 386806 239231 386858 239237
rect 386806 239173 386858 239179
rect 386710 239157 386762 239163
rect 386710 239099 386762 239105
rect 387106 238645 387134 246494
rect 387586 239015 387614 246494
rect 387682 246480 387936 246508
rect 388162 246480 388416 246508
rect 387574 239009 387626 239015
rect 387574 238951 387626 238957
rect 387094 238639 387146 238645
rect 387094 238581 387146 238587
rect 385942 237307 385994 237313
rect 385942 237249 385994 237255
rect 387682 237239 387710 246480
rect 388162 239903 388190 246480
rect 388546 245051 388574 246573
rect 388726 245817 388778 245823
rect 388726 245759 388778 245765
rect 388738 245051 388766 245759
rect 388532 245042 388588 245051
rect 388532 244977 388588 244986
rect 388724 245042 388780 245051
rect 388724 244977 388780 244986
rect 388534 244855 388586 244861
rect 388534 244797 388586 244803
rect 388546 244755 388574 244797
rect 388532 244746 388588 244755
rect 388532 244681 388588 244690
rect 388150 239897 388202 239903
rect 388150 239839 388202 239845
rect 388834 238497 388862 246494
rect 389026 245051 389054 246647
rect 389012 245042 389068 245051
rect 389012 244977 389068 244986
rect 389218 238941 389246 246494
rect 389506 246489 389534 246721
rect 392578 246711 392606 246753
rect 392566 246705 392618 246711
rect 392566 246647 392618 246653
rect 389782 246557 389834 246563
rect 389782 246499 389834 246505
rect 389494 246483 389546 246489
rect 389494 246425 389546 246431
rect 389206 238935 389258 238941
rect 389206 238877 389258 238883
rect 388822 238491 388874 238497
rect 388822 238433 388874 238439
rect 389698 238275 389726 246494
rect 389794 245231 389822 246499
rect 389890 246480 390144 246508
rect 390370 246480 390624 246508
rect 389782 245225 389834 245231
rect 389782 245167 389834 245173
rect 389782 244929 389834 244935
rect 389782 244871 389834 244877
rect 389794 244713 389822 244871
rect 389782 244707 389834 244713
rect 389782 244649 389834 244655
rect 389890 240167 389918 246480
rect 389876 240158 389932 240167
rect 389876 240093 389932 240102
rect 390370 238349 390398 246480
rect 390358 238343 390410 238349
rect 390358 238285 390410 238291
rect 389686 238269 389738 238275
rect 389686 238211 389738 238217
rect 387670 237233 387722 237239
rect 387670 237175 387722 237181
rect 390946 236721 390974 246494
rect 391426 238095 391454 246494
rect 391906 238201 391934 246494
rect 392098 246480 392352 246508
rect 392482 246480 392736 246508
rect 391990 246261 392042 246267
rect 391990 246203 392042 246209
rect 392002 245971 392030 246203
rect 391990 245965 392042 245971
rect 391990 245907 392042 245913
rect 392098 239459 392126 246480
rect 392086 239453 392138 239459
rect 392086 239395 392138 239401
rect 391894 238195 391946 238201
rect 391894 238137 391946 238143
rect 391412 238086 391468 238095
rect 392482 238053 392510 246480
rect 392962 245749 392990 246753
rect 393046 246721 393098 246727
rect 393334 246779 393386 246785
rect 393428 246753 393484 246762
rect 403318 246779 403370 246785
rect 393334 246721 393386 246727
rect 393058 246267 393086 246721
rect 393046 246261 393098 246267
rect 393046 246203 393098 246209
rect 392950 245743 393002 245749
rect 392950 245685 393002 245691
rect 391412 238021 391468 238030
rect 392470 238047 392522 238053
rect 392470 237989 392522 237995
rect 393154 237947 393182 246494
rect 393346 246193 393374 246721
rect 393442 246711 393470 246753
rect 403318 246721 403370 246727
rect 393430 246705 393482 246711
rect 393430 246647 393482 246653
rect 393334 246187 393386 246193
rect 393334 246129 393386 246135
rect 393634 238423 393662 246494
rect 394114 239311 394142 246494
rect 394210 246480 394464 246508
rect 394690 246480 394944 246508
rect 394102 239305 394154 239311
rect 394102 239247 394154 239253
rect 393622 238417 393674 238423
rect 393622 238359 393674 238365
rect 394210 238127 394238 246480
rect 394198 238121 394250 238127
rect 394198 238063 394250 238069
rect 393140 237938 393196 237947
rect 393140 237873 393196 237882
rect 394690 237799 394718 246480
rect 395362 238687 395390 246494
rect 395842 241901 395870 246494
rect 395830 241895 395882 241901
rect 395830 241837 395882 241843
rect 395348 238678 395404 238687
rect 395348 238613 395404 238622
rect 394676 237790 394732 237799
rect 394676 237725 394732 237734
rect 396226 237461 396254 246494
rect 396418 246480 396672 246508
rect 396898 246480 397152 246508
rect 396418 239681 396446 246480
rect 396406 239675 396458 239681
rect 396406 239617 396458 239623
rect 396898 239237 396926 246480
rect 397474 241309 397502 246494
rect 397462 241303 397514 241309
rect 397462 241245 397514 241251
rect 396886 239231 396938 239237
rect 396886 239173 396938 239179
rect 397954 237535 397982 246494
rect 398434 241087 398462 246494
rect 398626 246480 398880 246508
rect 399010 246480 399264 246508
rect 398422 241081 398474 241087
rect 398422 241023 398474 241029
rect 398626 239607 398654 246480
rect 399010 241013 399038 246480
rect 398998 241007 399050 241013
rect 398998 240949 399050 240955
rect 398614 239601 398666 239607
rect 398614 239543 398666 239549
rect 399682 237609 399710 246494
rect 400162 241457 400190 246494
rect 400150 241451 400202 241457
rect 400150 241393 400202 241399
rect 400642 239089 400670 246494
rect 400738 246480 400992 246508
rect 401218 246480 401472 246508
rect 400738 241235 400766 246480
rect 400918 245965 400970 245971
rect 400918 245907 400970 245913
rect 400930 244755 400958 245907
rect 400916 244746 400972 244755
rect 400916 244681 400972 244690
rect 400726 241229 400778 241235
rect 400726 241171 400778 241177
rect 400630 239083 400682 239089
rect 400630 239025 400682 239031
rect 401218 237979 401246 246480
rect 401494 245891 401546 245897
rect 401494 245833 401546 245839
rect 401506 245051 401534 245833
rect 401492 245042 401548 245051
rect 401492 244977 401548 244986
rect 401890 241383 401918 246494
rect 401878 241377 401930 241383
rect 401878 241319 401930 241325
rect 402370 240019 402398 246494
rect 402754 241161 402782 246494
rect 403200 246480 403262 246508
rect 402742 241155 402794 241161
rect 402742 241097 402794 241103
rect 403234 240273 403262 246480
rect 403330 245051 403358 246721
rect 403798 246705 403850 246711
rect 403798 246647 403850 246653
rect 403426 246480 403680 246508
rect 403316 245042 403372 245051
rect 403316 244977 403372 244986
rect 403426 240643 403454 246480
rect 403810 244607 403838 246647
rect 404374 246557 404426 246563
rect 404374 246499 404426 246505
rect 403894 246187 403946 246193
rect 403894 246129 403946 246135
rect 403906 244755 403934 246129
rect 403892 244746 403948 244755
rect 403892 244681 403948 244690
rect 403796 244598 403852 244607
rect 403796 244533 403852 244542
rect 403414 240637 403466 240643
rect 403414 240579 403466 240585
rect 403222 240267 403274 240273
rect 403222 240209 403274 240215
rect 404098 240199 404126 246494
rect 404386 245051 404414 246499
rect 404372 245042 404428 245051
rect 404372 244977 404428 244986
rect 404372 244746 404428 244755
rect 404372 244681 404374 244690
rect 404426 244681 404428 244690
rect 404374 244649 404426 244655
rect 404482 240791 404510 246494
rect 404962 241753 404990 246494
rect 405142 246483 405194 246489
rect 405142 246425 405194 246431
rect 405250 246480 405408 246508
rect 405538 246480 405792 246508
rect 406114 246480 406272 246508
rect 405154 245051 405182 246425
rect 405140 245042 405196 245051
rect 405140 244977 405196 244986
rect 404950 241747 405002 241753
rect 404950 241689 405002 241695
rect 404470 240785 404522 240791
rect 404470 240727 404522 240733
rect 405250 240569 405278 246480
rect 405238 240563 405290 240569
rect 405238 240505 405290 240511
rect 404086 240193 404138 240199
rect 404086 240135 404138 240141
rect 405538 240051 405566 246480
rect 406114 240939 406142 246480
rect 406102 240933 406154 240939
rect 406102 240875 406154 240881
rect 405526 240045 405578 240051
rect 402356 240010 402412 240019
rect 405526 239987 405578 239993
rect 402356 239945 402412 239954
rect 406690 239385 406718 246494
rect 407062 245225 407114 245231
rect 407062 245167 407114 245173
rect 407074 245051 407102 245167
rect 407060 245042 407116 245051
rect 407060 244977 407116 244986
rect 407170 240865 407198 246494
rect 407158 240859 407210 240865
rect 407158 240801 407210 240807
rect 407554 240347 407582 246494
rect 407746 246480 408000 246508
rect 408226 246480 408480 246508
rect 407746 240495 407774 246480
rect 407734 240489 407786 240495
rect 407734 240431 407786 240437
rect 408226 240421 408254 246480
rect 408898 240717 408926 246494
rect 409174 246261 409226 246267
rect 409174 246203 409226 246209
rect 409186 245051 409214 246203
rect 409172 245042 409228 245051
rect 409172 244977 409228 244986
rect 409282 241827 409310 246494
rect 409270 241821 409322 241827
rect 409270 241763 409322 241769
rect 408886 240711 408938 240717
rect 408886 240653 408938 240659
rect 409762 240611 409790 246494
rect 409954 246480 410208 246508
rect 410434 246480 410688 246508
rect 409954 241679 409982 246480
rect 409942 241673 409994 241679
rect 409942 241615 409994 241621
rect 409748 240602 409804 240611
rect 409748 240537 409804 240546
rect 408214 240415 408266 240421
rect 408214 240357 408266 240363
rect 407542 240341 407594 240347
rect 407542 240283 407594 240289
rect 406678 239379 406730 239385
rect 406678 239321 406730 239327
rect 401206 237973 401258 237979
rect 401206 237915 401258 237921
rect 410434 237905 410462 246480
rect 410422 237899 410474 237905
rect 410422 237841 410474 237847
rect 411010 237831 411038 246494
rect 411490 240463 411518 246494
rect 411476 240454 411532 240463
rect 411476 240389 411532 240398
rect 410998 237825 411050 237831
rect 410998 237767 411050 237773
rect 411970 237651 411998 246494
rect 411956 237642 412012 237651
rect 399670 237603 399722 237609
rect 411956 237577 412012 237586
rect 420598 237603 420650 237609
rect 399670 237545 399722 237551
rect 420598 237545 420650 237551
rect 397942 237529 397994 237535
rect 397942 237471 397994 237477
rect 396214 237455 396266 237461
rect 396214 237397 396266 237403
rect 390934 236715 390986 236721
rect 390934 236657 390986 236663
rect 420610 236467 420638 237545
rect 497506 236763 497534 251605
rect 625186 249153 625214 253381
rect 613462 249147 613514 249153
rect 613462 249089 613514 249095
rect 625174 249147 625226 249153
rect 625174 249089 625226 249095
rect 504022 246113 504074 246119
rect 504022 246055 504074 246061
rect 504034 242091 504062 246055
rect 509782 246039 509834 246045
rect 509782 245981 509834 245987
rect 509794 242239 509822 245981
rect 613474 244861 613502 249089
rect 608182 244855 608234 244861
rect 608182 244797 608234 244803
rect 613462 244855 613514 244861
rect 613462 244797 613514 244803
rect 509780 242230 509836 242239
rect 509780 242165 509836 242174
rect 504020 242082 504076 242091
rect 504020 242017 504076 242026
rect 497492 236754 497548 236763
rect 497492 236689 497548 236698
rect 420596 236458 420652 236467
rect 420596 236393 420652 236402
rect 420610 233470 420638 236393
rect 497506 233470 497534 236689
rect 504034 233484 504062 242017
rect 509794 233484 509822 242165
rect 549238 237677 549290 237683
rect 549238 237619 549290 237625
rect 549250 236203 549278 237619
rect 608194 237609 608222 244797
rect 639298 237961 639326 256341
rect 639766 238343 639818 238349
rect 639766 238285 639818 238291
rect 639202 237933 639326 237961
rect 639382 237973 639434 237979
rect 637942 237899 637994 237905
rect 637942 237841 637994 237847
rect 637366 237751 637418 237757
rect 637366 237693 637418 237699
rect 608182 237603 608234 237609
rect 608182 237545 608234 237551
rect 541462 236197 541514 236203
rect 541462 236139 541514 236145
rect 549238 236197 549290 236203
rect 549238 236139 549290 236145
rect 541474 234691 541502 236139
rect 541460 234682 541516 234691
rect 541460 234617 541516 234626
rect 549250 233484 549278 236139
rect 637378 233780 637406 237693
rect 637846 237603 637898 237609
rect 637846 237545 637898 237551
rect 637330 233752 637406 233780
rect 637076 233646 637132 233655
rect 637076 233581 637132 233590
rect 504034 233456 505584 233484
rect 509794 233456 510384 233484
rect 549024 233456 549278 233484
rect 637090 233484 637118 233581
rect 637330 233484 637358 233752
rect 637090 233470 637358 233484
rect 637556 233498 637612 233507
rect 637090 233456 637344 233470
rect 214292 233433 214348 233442
rect 637858 233484 637886 237545
rect 637954 233507 637982 237841
rect 638902 237825 638954 237831
rect 638902 237767 638954 237773
rect 638710 236197 638762 236203
rect 638710 236139 638762 236145
rect 638722 233803 638750 236139
rect 638132 233794 638188 233803
rect 638132 233729 638188 233738
rect 638708 233794 638764 233803
rect 638708 233729 638764 233738
rect 637612 233456 637886 233484
rect 637940 233498 637996 233507
rect 637556 233433 637612 233442
rect 638146 233484 638174 233729
rect 638516 233646 638572 233655
rect 638516 233581 638572 233590
rect 638530 233484 638558 233581
rect 638914 233484 638942 237767
rect 639202 236203 639230 237933
rect 639382 237915 639434 237921
rect 639394 237776 639422 237915
rect 639298 237748 639422 237776
rect 639190 236197 639242 236203
rect 639190 236139 639242 236145
rect 637996 233456 638064 233484
rect 638146 233456 638448 233484
rect 638530 233456 638942 233484
rect 638996 233498 639052 233507
rect 637940 233433 637996 233442
rect 639298 233484 639326 237748
rect 639052 233456 639326 233484
rect 638996 233433 639052 233442
rect 639778 232892 639806 238285
rect 649570 237831 649598 927373
rect 649666 801383 649694 987609
rect 649750 986631 649802 986637
rect 649750 986573 649802 986579
rect 649652 801374 649708 801383
rect 649652 801309 649708 801318
rect 649654 748869 649706 748875
rect 649654 748811 649706 748817
rect 649558 237825 649610 237831
rect 649558 237767 649610 237773
rect 639552 232864 639806 232892
rect 645718 232941 645770 232947
rect 645718 232883 645770 232889
rect 218998 54305 219050 54311
rect 212372 54270 212428 54279
rect 212372 54205 212428 54214
rect 214388 54270 214444 54279
rect 214444 54228 214512 54256
rect 218928 54253 218998 54256
rect 218928 54247 219050 54253
rect 221014 54305 221066 54311
rect 221014 54247 221066 54253
rect 216322 54237 216350 54242
rect 216310 54231 216362 54237
rect 214388 54205 214444 54214
rect 212386 53793 212414 54205
rect 218928 54228 219038 54247
rect 216310 54173 216362 54179
rect 219190 54157 219242 54163
rect 214772 54122 214828 54131
rect 214828 54080 214896 54108
rect 219242 54105 219312 54108
rect 219190 54099 219312 54105
rect 218998 54083 219050 54089
rect 214772 54057 214828 54066
rect 219202 54080 219312 54099
rect 218998 54025 219050 54031
rect 218806 54009 218858 54015
rect 216596 53974 216652 53983
rect 216652 53932 216720 53960
rect 218806 53951 218858 53957
rect 216596 53909 216652 53918
rect 216790 53861 216842 53867
rect 216790 53803 216842 53809
rect 216980 53826 217036 53835
rect 212374 53787 212426 53793
rect 212374 53729 212426 53735
rect 210754 53636 211008 53664
rect 210358 53491 210410 53497
rect 210358 53433 210410 53439
rect 209878 51715 209930 51721
rect 209878 51657 209930 51663
rect 209492 48942 209548 48951
rect 209492 48877 209548 48886
rect 209014 48829 209066 48835
rect 209014 48771 209066 48777
rect 208918 48681 208970 48687
rect 208918 48623 208970 48629
rect 208822 48533 208874 48539
rect 208822 48475 208874 48481
rect 208726 48385 208778 48391
rect 208726 48327 208778 48333
rect 207862 46757 207914 46763
rect 207862 46699 207914 46705
rect 207766 46313 207818 46319
rect 207766 46255 207818 46261
rect 206902 42169 206954 42175
rect 206902 42111 206954 42117
rect 187604 41838 187660 41847
rect 187344 41796 187604 41824
rect 194324 41838 194380 41847
rect 194064 41796 194324 41824
rect 187604 41773 187660 41782
rect 194324 41773 194380 41782
rect 210754 40811 210782 53636
rect 211186 53368 211214 53650
rect 211378 53368 211406 53650
rect 211570 53571 211598 53650
rect 211558 53565 211610 53571
rect 211558 53507 211610 53513
rect 211186 53340 211262 53368
rect 211378 53340 211454 53368
rect 211234 52387 211262 53340
rect 211222 52381 211274 52387
rect 211222 52323 211274 52329
rect 211426 45283 211454 53340
rect 211714 45357 211742 53650
rect 211906 51911 211934 53650
rect 211892 51902 211948 51911
rect 211892 51837 211948 51846
rect 211702 45351 211754 45357
rect 211702 45293 211754 45299
rect 211414 45277 211466 45283
rect 211414 45219 211466 45225
rect 212098 45103 212126 53650
rect 212304 53636 212414 53664
rect 212182 52677 212234 52683
rect 212182 52619 212234 52625
rect 212194 52091 212222 52619
rect 212386 52091 212414 53636
rect 212182 52085 212234 52091
rect 212182 52027 212234 52033
rect 212374 52085 212426 52091
rect 212374 52027 212426 52033
rect 212084 45094 212140 45103
rect 212084 45029 212140 45038
rect 212482 42397 212510 53650
rect 212674 52059 212702 53650
rect 212660 52050 212716 52059
rect 212660 51985 212716 51994
rect 212866 44955 212894 53650
rect 213058 53539 213086 53650
rect 213216 53636 213278 53664
rect 213044 53530 213100 53539
rect 213044 53465 213100 53474
rect 212852 44946 212908 44955
rect 212852 44881 212908 44890
rect 213250 43285 213278 53636
rect 213394 53405 213422 53650
rect 213346 53377 213422 53405
rect 213346 53201 213374 53377
rect 213586 53368 213614 53650
rect 213730 53636 213792 53664
rect 213586 53340 213662 53368
rect 213334 53195 213386 53201
rect 213334 53137 213386 53143
rect 213430 52085 213482 52091
rect 213430 52027 213482 52033
rect 213442 51869 213470 52027
rect 213430 51863 213482 51869
rect 213430 51805 213482 51811
rect 213238 43279 213290 43285
rect 213238 43221 213290 43227
rect 212470 42391 212522 42397
rect 212470 42333 212522 42339
rect 213634 42101 213662 53340
rect 213730 51795 213758 53636
rect 213718 51789 213770 51795
rect 213718 51731 213770 51737
rect 213922 45209 213950 53650
rect 214114 51721 214142 53650
rect 214102 51715 214154 51721
rect 214102 51657 214154 51663
rect 213910 45203 213962 45209
rect 213910 45145 213962 45151
rect 213622 42095 213674 42101
rect 213622 42037 213674 42043
rect 214306 42027 214334 53650
rect 214690 45135 214718 53650
rect 214678 45129 214730 45135
rect 214678 45071 214730 45077
rect 215074 45061 215102 53650
rect 215266 53391 215294 53650
rect 215424 53636 215486 53664
rect 215252 53382 215308 53391
rect 215252 53317 215308 53326
rect 215062 45055 215114 45061
rect 215062 44997 215114 45003
rect 215458 44987 215486 53636
rect 215602 53479 215630 53650
rect 215554 53451 215630 53479
rect 215554 53275 215582 53451
rect 215794 53405 215822 53650
rect 215938 53636 216000 53664
rect 215938 53539 215966 53636
rect 215924 53530 215980 53539
rect 215924 53465 215980 53474
rect 215746 53377 215822 53405
rect 215542 53269 215594 53275
rect 215542 53211 215594 53217
rect 215746 53127 215774 53377
rect 215734 53121 215786 53127
rect 216022 53121 216074 53127
rect 215734 53063 215786 53069
rect 216020 53086 216022 53095
rect 216074 53086 216076 53095
rect 216020 53021 216076 53030
rect 216130 52461 216158 53650
rect 216118 52455 216170 52461
rect 216118 52397 216170 52403
rect 216514 47725 216542 53650
rect 216598 53565 216650 53571
rect 216802 53539 216830 53803
rect 217036 53784 217104 53812
rect 216980 53761 217036 53770
rect 216598 53507 216650 53513
rect 216788 53530 216844 53539
rect 216610 51795 216638 53507
rect 216788 53465 216844 53474
rect 216598 51789 216650 51795
rect 216598 51731 216650 51737
rect 216898 50389 216926 53650
rect 217282 52609 217310 53650
rect 217474 53423 217502 53650
rect 217632 53636 217694 53664
rect 217462 53417 217514 53423
rect 217462 53359 217514 53365
rect 217270 52603 217322 52609
rect 217270 52545 217322 52551
rect 217270 51197 217322 51203
rect 217270 51139 217322 51145
rect 216886 50383 216938 50389
rect 216886 50325 216938 50331
rect 217282 50241 217310 51139
rect 217270 50235 217322 50241
rect 217270 50177 217322 50183
rect 216502 47719 216554 47725
rect 216502 47661 216554 47667
rect 217666 47651 217694 53636
rect 217810 53497 217838 53650
rect 217798 53491 217850 53497
rect 217798 53433 217850 53439
rect 218002 53368 218030 53650
rect 217954 53340 218030 53368
rect 218146 53636 218208 53664
rect 217654 47645 217706 47651
rect 217654 47587 217706 47593
rect 217954 47577 217982 53340
rect 218146 53053 218174 53636
rect 218134 53047 218186 53053
rect 218134 52989 218186 52995
rect 217942 47571 217994 47577
rect 217942 47513 217994 47519
rect 218338 47503 218366 53650
rect 218326 47497 218378 47503
rect 218326 47439 218378 47445
rect 218530 46467 218558 53650
rect 218722 47429 218750 53650
rect 218818 53423 218846 53951
rect 219010 53497 219038 54025
rect 219190 53935 219242 53941
rect 219190 53877 219242 53883
rect 218998 53491 219050 53497
rect 218998 53433 219050 53439
rect 218806 53417 218858 53423
rect 218806 53359 218858 53365
rect 219106 47799 219134 53650
rect 219202 53571 219230 53877
rect 219190 53565 219242 53571
rect 219190 53507 219242 53513
rect 219490 49649 219518 53650
rect 219682 53349 219710 53650
rect 219826 53571 219854 53650
rect 219814 53565 219866 53571
rect 220018 53539 220046 53650
rect 219814 53507 219866 53513
rect 220004 53530 220060 53539
rect 220004 53465 220060 53474
rect 220210 53368 220238 53650
rect 219670 53343 219722 53349
rect 219670 53285 219722 53291
rect 219862 53343 219914 53349
rect 219862 53285 219914 53291
rect 220162 53340 220238 53368
rect 220354 53636 220416 53664
rect 219874 52905 219902 53285
rect 219862 52899 219914 52905
rect 219862 52841 219914 52847
rect 219478 49643 219530 49649
rect 219478 49585 219530 49591
rect 220162 47947 220190 53340
rect 220354 53243 220382 53636
rect 220340 53234 220396 53243
rect 220340 53169 220396 53178
rect 220546 48909 220574 53650
rect 220738 48951 220766 53650
rect 220930 52683 220958 53650
rect 221026 53571 221054 54247
rect 221136 53793 221246 53812
rect 221136 53787 221258 53793
rect 221136 53784 221206 53787
rect 221206 53729 221258 53735
rect 293782 53713 293834 53719
rect 221014 53565 221066 53571
rect 221014 53507 221066 53513
rect 220918 52677 220970 52683
rect 220918 52619 220970 52625
rect 220724 48942 220780 48951
rect 220534 48903 220586 48909
rect 220724 48877 220780 48886
rect 220534 48845 220586 48851
rect 220150 47941 220202 47947
rect 220150 47883 220202 47889
rect 221314 47873 221342 53650
rect 221506 49871 221534 53650
rect 221494 49865 221546 49871
rect 221494 49807 221546 49813
rect 221698 48761 221726 53650
rect 221782 52307 221834 52313
rect 221782 52249 221834 52255
rect 221794 51647 221822 52249
rect 221890 51763 221918 53650
rect 222048 53636 222110 53664
rect 221876 51754 221932 51763
rect 221876 51689 221932 51698
rect 221782 51641 221834 51647
rect 221782 51583 221834 51589
rect 222082 48835 222110 53636
rect 222226 53368 222254 53650
rect 222418 53368 222446 53650
rect 222226 53340 222302 53368
rect 222274 48835 222302 53340
rect 222370 53340 222446 53368
rect 222562 53636 222624 53664
rect 222070 48829 222122 48835
rect 222070 48771 222122 48777
rect 222262 48829 222314 48835
rect 222262 48771 222314 48777
rect 221686 48755 221738 48761
rect 221686 48697 221738 48703
rect 222370 48687 222398 53340
rect 222562 52207 222590 53636
rect 222548 52198 222604 52207
rect 222548 52133 222604 52142
rect 222358 48681 222410 48687
rect 222358 48623 222410 48629
rect 222754 48539 222782 53650
rect 222946 48909 222974 53650
rect 222934 48903 222986 48909
rect 222934 48845 222986 48851
rect 222742 48533 222794 48539
rect 222742 48475 222794 48481
rect 223138 48095 223166 53650
rect 223330 51615 223358 53650
rect 223316 51606 223372 51615
rect 223316 51541 223372 51550
rect 223126 48089 223178 48095
rect 223126 48031 223178 48037
rect 223522 48021 223550 53650
rect 223714 48983 223742 53650
rect 223702 48977 223754 48983
rect 223702 48919 223754 48925
rect 223906 48391 223934 53650
rect 224098 48761 224126 53650
rect 224256 53636 224318 53664
rect 224290 50315 224318 53636
rect 224626 53368 224654 53650
rect 224578 53340 224654 53368
rect 224278 50309 224330 50315
rect 224278 50251 224330 50257
rect 224086 48755 224138 48761
rect 224086 48697 224138 48703
rect 223894 48385 223946 48391
rect 223894 48327 223946 48333
rect 224578 48169 224606 53340
rect 224566 48163 224618 48169
rect 224566 48105 224618 48111
rect 223510 48015 223562 48021
rect 223510 47957 223562 47963
rect 221302 47867 221354 47873
rect 221302 47809 221354 47815
rect 219094 47793 219146 47799
rect 219094 47735 219146 47741
rect 218710 47423 218762 47429
rect 218710 47365 218762 47371
rect 224962 46763 224990 53650
rect 225346 49797 225374 53650
rect 225730 52165 225758 53650
rect 225718 52159 225770 52165
rect 225718 52101 225770 52107
rect 225334 49791 225386 49797
rect 225334 49733 225386 49739
rect 226114 48243 226142 53650
rect 226464 53636 226526 53664
rect 226102 48237 226154 48243
rect 226102 48179 226154 48185
rect 224950 46757 225002 46763
rect 224950 46699 225002 46705
rect 225046 46757 225098 46763
rect 225046 46699 225098 46705
rect 218518 46461 218570 46467
rect 218518 46403 218570 46409
rect 225058 46319 225086 46699
rect 226498 46689 226526 53636
rect 226594 53636 226848 53664
rect 226594 49723 226622 53636
rect 227170 52239 227198 53650
rect 227446 52381 227498 52387
rect 227446 52323 227498 52329
rect 227158 52233 227210 52239
rect 227158 52175 227210 52181
rect 227458 51351 227486 52323
rect 227554 51943 227582 53650
rect 227542 51937 227594 51943
rect 227542 51879 227594 51885
rect 227446 51345 227498 51351
rect 227446 51287 227498 51293
rect 226582 49717 226634 49723
rect 226582 49659 226634 49665
rect 227938 46763 227966 53650
rect 228322 50685 228350 53650
rect 228418 53636 228672 53664
rect 228802 53636 229056 53664
rect 228310 50679 228362 50685
rect 228310 50621 228362 50627
rect 228418 50463 228446 53636
rect 228802 50759 228830 53636
rect 228790 50753 228842 50759
rect 228790 50695 228842 50701
rect 229378 50537 229406 53650
rect 229762 50611 229790 53650
rect 229750 50605 229802 50611
rect 229750 50547 229802 50553
rect 229366 50531 229418 50537
rect 229366 50473 229418 50479
rect 228406 50457 228458 50463
rect 228406 50399 228458 50405
rect 229652 50422 229708 50431
rect 229652 50357 229708 50366
rect 229666 48983 229694 50357
rect 229654 48977 229706 48983
rect 229654 48919 229706 48925
rect 230146 46911 230174 53650
rect 230134 46905 230186 46911
rect 230134 46847 230186 46853
rect 227926 46757 227978 46763
rect 227926 46699 227978 46705
rect 226486 46683 226538 46689
rect 226486 46625 226538 46631
rect 230530 46541 230558 53650
rect 230626 53636 230880 53664
rect 231010 53636 231264 53664
rect 230626 50833 230654 53636
rect 231010 50907 231038 53636
rect 230998 50901 231050 50907
rect 230998 50843 231050 50849
rect 230614 50827 230666 50833
rect 230614 50769 230666 50775
rect 231586 46837 231614 53650
rect 231970 50981 231998 53650
rect 232354 51129 232382 53650
rect 232342 51123 232394 51129
rect 232342 51065 232394 51071
rect 232738 51055 232766 53650
rect 232834 53636 233088 53664
rect 233314 53636 233472 53664
rect 232726 51049 232778 51055
rect 232726 50991 232778 50997
rect 231958 50975 232010 50981
rect 231958 50917 232010 50923
rect 232834 49945 232862 53636
rect 232822 49939 232874 49945
rect 232822 49881 232874 49887
rect 233314 47133 233342 53636
rect 233794 51277 233822 53650
rect 233782 51271 233834 51277
rect 233782 51213 233834 51219
rect 233302 47127 233354 47133
rect 233302 47069 233354 47075
rect 231574 46831 231626 46837
rect 231574 46773 231626 46779
rect 234178 46615 234206 53650
rect 234562 50167 234590 53650
rect 234550 50161 234602 50167
rect 234550 50103 234602 50109
rect 234946 50093 234974 53650
rect 235042 53636 235296 53664
rect 235426 53636 235680 53664
rect 234934 50087 234986 50093
rect 234934 50029 234986 50035
rect 235042 48613 235070 53636
rect 235426 51203 235454 53636
rect 235414 51197 235466 51203
rect 235414 51139 235466 51145
rect 236002 50241 236030 53650
rect 236386 51499 236414 53650
rect 236374 51493 236426 51499
rect 236374 51435 236426 51441
rect 235990 50235 236042 50241
rect 235990 50177 236042 50183
rect 235030 48607 235082 48613
rect 235030 48549 235082 48555
rect 234166 46609 234218 46615
rect 234166 46551 234218 46557
rect 230518 46535 230570 46541
rect 230518 46477 230570 46483
rect 225046 46313 225098 46319
rect 225046 46255 225098 46261
rect 236770 46245 236798 53650
rect 237154 51425 237182 53650
rect 237250 53636 237504 53664
rect 237634 53636 237888 53664
rect 237142 51419 237194 51425
rect 237142 51361 237194 51367
rect 237250 50019 237278 53636
rect 237634 51573 237662 53636
rect 237622 51567 237674 51573
rect 237622 51509 237674 51515
rect 238210 51319 238238 53650
rect 238196 51310 238252 51319
rect 238196 51245 238252 51254
rect 237238 50013 237290 50019
rect 237238 49955 237290 49961
rect 238594 47355 238622 53650
rect 238582 47349 238634 47355
rect 238582 47291 238634 47297
rect 238978 47059 239006 53650
rect 239362 47207 239390 53650
rect 239458 53636 239712 53664
rect 239842 53636 240096 53664
rect 239350 47201 239402 47207
rect 239350 47143 239402 47149
rect 238966 47053 239018 47059
rect 238966 46995 239018 47001
rect 239458 46393 239486 53636
rect 239446 46387 239498 46393
rect 239446 46329 239498 46335
rect 236758 46239 236810 46245
rect 236758 46181 236810 46187
rect 239842 46171 239870 53636
rect 240418 47281 240446 53650
rect 240406 47275 240458 47281
rect 240406 47217 240458 47223
rect 240802 46985 240830 53650
rect 241186 48465 241214 53650
rect 241174 48459 241226 48465
rect 241174 48401 241226 48407
rect 241570 48317 241598 53650
rect 241920 53636 241982 53664
rect 241558 48311 241610 48317
rect 241558 48253 241610 48259
rect 241954 48211 241982 53636
rect 242050 53636 242304 53664
rect 242050 48655 242078 53636
rect 242036 48646 242092 48655
rect 242036 48581 242092 48590
rect 241940 48202 241996 48211
rect 241940 48137 241996 48146
rect 242626 47915 242654 53650
rect 243010 48507 243038 53650
rect 243394 51467 243422 53650
rect 243380 51458 243436 51467
rect 243380 51393 243436 51402
rect 242996 48498 243052 48507
rect 242996 48433 243052 48442
rect 243778 48359 243806 53650
rect 243874 53636 244128 53664
rect 293782 53655 293834 53661
rect 243874 51647 243902 53636
rect 287938 51721 288062 51740
rect 287926 51715 288074 51721
rect 287978 51712 288022 51715
rect 287926 51657 287978 51663
rect 288022 51657 288074 51663
rect 292054 51715 292106 51721
rect 292054 51657 292106 51663
rect 243862 51641 243914 51647
rect 243862 51583 243914 51589
rect 292066 51573 292094 51657
rect 292054 51567 292106 51573
rect 292054 51509 292106 51515
rect 243764 48350 243820 48359
rect 243764 48285 243820 48294
rect 242612 47906 242668 47915
rect 242612 47841 242668 47850
rect 240790 46979 240842 46985
rect 240790 46921 240842 46927
rect 239830 46165 239882 46171
rect 239830 46107 239882 46113
rect 293794 45875 293822 53655
rect 330934 53639 330986 53645
rect 330934 53581 330986 53587
rect 308086 53269 308138 53275
rect 308138 53217 308222 53220
rect 308086 53211 308222 53217
rect 308098 53201 308222 53211
rect 308098 53195 308234 53201
rect 308098 53192 308182 53195
rect 308182 53137 308234 53143
rect 330946 51647 330974 53581
rect 403126 53565 403178 53571
rect 403126 53507 403178 53513
rect 348406 53269 348458 53275
rect 348458 53217 348542 53220
rect 348406 53211 348542 53217
rect 348418 53201 348542 53211
rect 348418 53195 348554 53201
rect 348418 53192 348502 53195
rect 348502 53137 348554 53143
rect 403138 51740 403166 53507
rect 452182 53491 452234 53497
rect 452182 53433 452234 53439
rect 420502 53269 420554 53275
rect 443542 53269 443594 53275
rect 420554 53229 420638 53257
rect 420502 53211 420554 53217
rect 420610 53127 420638 53229
rect 443458 53217 443542 53220
rect 443458 53211 443594 53217
rect 443458 53192 443582 53211
rect 443458 53127 443486 53192
rect 420598 53121 420650 53127
rect 420598 53063 420650 53069
rect 443446 53121 443498 53127
rect 443446 53063 443498 53069
rect 423382 51937 423434 51943
rect 403234 51860 403454 51888
rect 423382 51879 423434 51885
rect 432790 51937 432842 51943
rect 432790 51879 432842 51885
rect 403234 51740 403262 51860
rect 348406 51715 348458 51721
rect 403138 51712 403262 51740
rect 403318 51715 403370 51721
rect 348406 51657 348458 51663
rect 403318 51657 403370 51663
rect 330934 51641 330986 51647
rect 330934 51583 330986 51589
rect 348310 51641 348362 51647
rect 348418 51629 348446 51657
rect 348502 51641 348554 51647
rect 348418 51601 348502 51629
rect 348310 51583 348362 51589
rect 348502 51583 348554 51589
rect 372022 51641 372074 51647
rect 403330 51592 403358 51657
rect 372074 51589 372158 51592
rect 372022 51583 372158 51589
rect 302422 51567 302474 51573
rect 302518 51567 302570 51573
rect 302474 51527 302518 51555
rect 302422 51509 302474 51515
rect 302518 51509 302570 51515
rect 322582 51567 322634 51573
rect 322582 51509 322634 51515
rect 322594 51425 322622 51509
rect 322582 51419 322634 51425
rect 322582 51361 322634 51367
rect 293782 45869 293834 45875
rect 293782 45811 293834 45817
rect 302326 45869 302378 45875
rect 302326 45811 302378 45817
rect 215446 44981 215498 44987
rect 215446 44923 215498 44929
rect 302338 42143 302366 45811
rect 327286 45351 327338 45357
rect 327286 45293 327338 45299
rect 302516 43318 302572 43327
rect 302516 43253 302572 43262
rect 302324 42134 302380 42143
rect 302530 42120 302558 43253
rect 310102 42391 310154 42397
rect 310102 42333 310154 42339
rect 306740 42134 306796 42143
rect 302530 42092 302688 42120
rect 302324 42069 302380 42078
rect 306796 42092 307008 42120
rect 310114 42106 310142 42333
rect 306740 42069 306796 42078
rect 214294 42021 214346 42027
rect 214294 41963 214346 41969
rect 327298 40811 327326 45293
rect 328054 45277 328106 45283
rect 328054 45219 328106 45225
rect 328066 40959 328094 45219
rect 348322 42915 348350 51583
rect 372034 51573 372158 51583
rect 403138 51573 403358 51592
rect 372034 51567 372170 51573
rect 372034 51564 372118 51567
rect 372118 51509 372170 51515
rect 403126 51567 403358 51573
rect 403178 51564 403358 51567
rect 403126 51509 403178 51515
rect 348310 42909 348362 42915
rect 348310 42851 348362 42857
rect 357430 42909 357482 42915
rect 357430 42851 357482 42857
rect 357442 42106 357470 42851
rect 403426 41879 403454 51860
rect 423394 51721 423422 51879
rect 423382 51715 423434 51721
rect 423382 51657 423434 51663
rect 432802 51647 432830 51879
rect 432790 51641 432842 51647
rect 432790 51583 432842 51589
rect 446902 45203 446954 45209
rect 446902 45145 446954 45151
rect 416564 43318 416620 43327
rect 411010 43285 411102 43304
rect 410998 43279 411102 43285
rect 411050 43276 411102 43279
rect 416564 43253 416620 43262
rect 410998 43221 411050 43227
rect 405238 42169 405290 42175
rect 405290 42117 405552 42120
rect 405238 42111 405552 42117
rect 405250 42092 405552 42111
rect 416578 42106 416606 43253
rect 446914 43211 446942 45145
rect 452194 43581 452222 53433
rect 466486 53417 466538 53423
rect 466486 53359 466538 53365
rect 463702 53269 463754 53275
rect 463702 53211 463754 53217
rect 463606 53195 463658 53201
rect 463714 53183 463742 53211
rect 463658 53155 463742 53183
rect 463606 53137 463658 53143
rect 452662 51641 452714 51647
rect 452714 51589 452798 51592
rect 452662 51583 452798 51589
rect 452674 51573 452798 51583
rect 452674 51567 452810 51573
rect 452674 51564 452758 51567
rect 452758 51509 452810 51515
rect 466498 49076 466526 53359
rect 517846 53343 517898 53349
rect 517846 53285 517898 53291
rect 483862 53269 483914 53275
rect 483862 53211 483914 53217
rect 483874 53053 483902 53211
rect 483862 53047 483914 53053
rect 483862 52989 483914 52995
rect 514006 53047 514058 53053
rect 514006 52989 514058 52995
rect 483862 51937 483914 51943
rect 483862 51879 483914 51885
rect 493846 51937 493898 51943
rect 493846 51879 493898 51885
rect 483874 51721 483902 51879
rect 469558 51715 469610 51721
rect 469378 51675 469558 51703
rect 469378 51647 469406 51675
rect 469558 51657 469610 51663
rect 483862 51715 483914 51721
rect 483862 51657 483914 51663
rect 469366 51641 469418 51647
rect 469366 51583 469418 51589
rect 493858 51573 493886 51879
rect 493846 51567 493898 51573
rect 493846 51509 493898 51515
rect 466498 49048 466622 49076
rect 466594 46139 466622 49048
rect 514018 47577 514046 52989
rect 514006 47571 514058 47577
rect 514006 47513 514058 47519
rect 466580 46130 466636 46139
rect 466580 46065 466636 46074
rect 506806 45129 506858 45135
rect 506806 45071 506858 45077
rect 506710 45055 506762 45061
rect 506710 44997 506762 45003
rect 452182 43575 452234 43581
rect 452182 43517 452234 43523
rect 461110 43575 461162 43581
rect 461110 43517 461162 43523
rect 446902 43205 446954 43211
rect 446902 43147 446954 43153
rect 454966 43205 455018 43211
rect 461122 43179 461150 43517
rect 454966 43147 455018 43153
rect 461108 43170 461164 43179
rect 403414 41873 403466 41879
rect 361460 41838 361516 41847
rect 364628 41838 364684 41847
rect 361516 41796 361776 41824
rect 361460 41773 361516 41782
rect 364684 41796 364944 41824
rect 403414 41815 403466 41821
rect 364628 41773 364684 41782
rect 328052 40950 328108 40959
rect 328052 40885 328108 40894
rect 210740 40802 210796 40811
rect 210740 40737 210796 40746
rect 327284 40802 327340 40811
rect 327284 40737 327340 40746
rect 454978 40367 455006 43147
rect 461108 43105 461164 43114
rect 465620 43170 465676 43179
rect 465676 43128 465842 43156
rect 465620 43105 465676 43114
rect 471092 42134 471148 42143
rect 460066 42101 460368 42120
rect 460054 42095 460368 42101
rect 460106 42092 460368 42095
rect 471148 42092 471408 42120
rect 471092 42069 471148 42078
rect 460054 42037 460106 42043
rect 463700 41838 463756 41847
rect 463756 41796 464016 41824
rect 506722 41805 506750 44997
rect 506818 41953 506846 45071
rect 517858 43327 517886 53285
rect 639682 51943 639710 232864
rect 645730 232471 645758 232883
rect 645716 232462 645772 232471
rect 645716 232397 645772 232406
rect 645142 232349 645194 232355
rect 645140 232314 645142 232323
rect 645526 232349 645578 232355
rect 645194 232314 645196 232323
rect 645526 232291 645578 232297
rect 645140 232249 645196 232258
rect 645142 231609 645194 231615
rect 645140 231574 645142 231583
rect 645194 231574 645196 231583
rect 645196 231532 645278 231560
rect 645140 231509 645196 231518
rect 645142 231165 645194 231171
rect 645140 231130 645142 231139
rect 645194 231130 645196 231139
rect 645140 231065 645196 231074
rect 645142 230721 645194 230727
rect 645140 230686 645142 230695
rect 645194 230686 645196 230695
rect 645140 230621 645196 230630
rect 640726 99371 640778 99377
rect 640726 99313 640778 99319
rect 544342 51937 544394 51943
rect 544342 51879 544394 51885
rect 552790 51937 552842 51943
rect 552790 51879 552842 51885
rect 625750 51937 625802 51943
rect 625750 51879 625802 51885
rect 639670 51937 639722 51943
rect 639670 51879 639722 51885
rect 544354 51647 544382 51879
rect 552802 51721 552830 51879
rect 610498 51721 610718 51740
rect 552790 51715 552842 51721
rect 552790 51657 552842 51663
rect 610486 51715 610718 51721
rect 610538 51712 610718 51715
rect 610486 51657 610538 51663
rect 610690 51647 610718 51712
rect 625762 51647 625790 51879
rect 544342 51641 544394 51647
rect 544342 51583 544394 51589
rect 610678 51641 610730 51647
rect 610678 51583 610730 51589
rect 625750 51641 625802 51647
rect 625750 51583 625802 51589
rect 525910 47571 525962 47577
rect 525910 47513 525962 47519
rect 517844 43318 517900 43327
rect 517844 43253 517900 43262
rect 520628 43318 520684 43327
rect 520628 43253 520684 43262
rect 520642 42106 520670 43253
rect 525922 42120 525950 47513
rect 526966 44981 527018 44987
rect 526966 44923 527018 44929
rect 526978 42143 527006 44923
rect 526964 42134 527020 42143
rect 525922 42092 526176 42120
rect 526964 42069 527020 42078
rect 528980 42134 529036 42143
rect 529036 42092 529296 42120
rect 528980 42069 529036 42078
rect 514870 42021 514922 42027
rect 521590 42021 521642 42027
rect 514922 41969 515136 41972
rect 514870 41963 515136 41969
rect 521642 41969 521856 41972
rect 521590 41963 521856 41969
rect 506806 41947 506858 41953
rect 514882 41944 515136 41963
rect 521602 41944 521856 41963
rect 506806 41889 506858 41895
rect 518530 41805 518832 41824
rect 506710 41799 506762 41805
rect 463700 41773 463756 41782
rect 506710 41741 506762 41747
rect 518518 41799 518832 41805
rect 518570 41796 518832 41799
rect 518518 41741 518570 41747
rect 640738 40663 640766 99313
rect 645154 48761 645182 230621
rect 645250 48835 645278 231532
rect 645334 231165 645386 231171
rect 645334 231107 645386 231113
rect 645346 48909 645374 231107
rect 645430 79687 645482 79693
rect 645430 79629 645482 79635
rect 645442 78551 645470 79629
rect 645428 78542 645484 78551
rect 645428 78477 645484 78486
rect 645538 51869 645566 232291
rect 645620 210410 645676 210419
rect 645620 210345 645676 210354
rect 645526 51863 645578 51869
rect 645526 51805 645578 51811
rect 645334 48903 645386 48909
rect 645334 48845 645386 48851
rect 645238 48829 645290 48835
rect 645238 48771 645290 48777
rect 645142 48755 645194 48761
rect 645142 48697 645194 48703
rect 645634 46467 645662 210345
rect 645730 51795 645758 232397
rect 649666 232355 649694 748811
rect 649762 707551 649790 986573
rect 649748 707542 649804 707551
rect 649748 707477 649804 707486
rect 649750 702767 649802 702773
rect 649750 702709 649802 702715
rect 649762 237979 649790 702709
rect 649858 660635 649886 994597
rect 658006 989295 658058 989301
rect 658006 989237 658058 989243
rect 650134 987741 650186 987747
rect 650134 987683 650186 987689
rect 650038 987593 650090 987599
rect 650038 987535 650090 987541
rect 649942 984929 649994 984935
rect 649942 984871 649994 984877
rect 649954 754615 649982 984871
rect 650050 895215 650078 987535
rect 650036 895206 650092 895215
rect 650036 895141 650092 895150
rect 650146 848299 650174 987683
rect 650998 986409 651050 986415
rect 650998 986351 651050 986357
rect 650132 848290 650188 848299
rect 650132 848225 650188 848234
rect 649940 754606 649996 754615
rect 649940 754541 649996 754550
rect 649844 660626 649900 660635
rect 649844 660561 649900 660570
rect 649846 656739 649898 656745
rect 649846 656681 649898 656687
rect 649750 237973 649802 237979
rect 649750 237915 649802 237921
rect 649858 232947 649886 656681
rect 649942 613523 649994 613529
rect 649942 613465 649994 613471
rect 649954 238349 649982 613465
rect 650038 567421 650090 567427
rect 650038 567363 650090 567369
rect 649942 238343 649994 238349
rect 649942 238285 649994 238291
rect 649846 232941 649898 232947
rect 649846 232883 649898 232889
rect 649654 232349 649706 232355
rect 649654 232291 649706 232297
rect 650050 230727 650078 567363
rect 650134 521319 650186 521325
rect 650134 521261 650186 521267
rect 650146 237757 650174 521261
rect 650230 478177 650282 478183
rect 650230 478119 650282 478125
rect 650134 237751 650186 237757
rect 650134 237693 650186 237699
rect 650242 237609 650270 478119
rect 650326 391745 650378 391751
rect 650326 391687 650378 391693
rect 650230 237603 650282 237609
rect 650230 237545 650282 237551
rect 650338 231171 650366 391687
rect 650422 345643 650474 345649
rect 650422 345585 650474 345591
rect 650434 237905 650462 345585
rect 650518 299615 650570 299621
rect 650518 299557 650570 299563
rect 650422 237899 650474 237905
rect 650422 237841 650474 237847
rect 650530 231615 650558 299557
rect 651010 237683 651038 986351
rect 655124 976754 655180 976763
rect 655124 976689 655180 976698
rect 654452 953370 654508 953379
rect 654452 953305 654508 953314
rect 654466 941941 654494 953305
rect 655138 944679 655166 976689
rect 655220 965062 655276 965071
rect 655220 964997 655276 965006
rect 655234 944901 655262 964997
rect 655222 944895 655274 944901
rect 655222 944837 655274 944843
rect 655126 944673 655178 944679
rect 655126 944615 655178 944621
rect 658018 942089 658046 989237
rect 660886 986557 660938 986563
rect 660886 986499 660938 986505
rect 658006 942083 658058 942089
rect 658006 942025 658058 942031
rect 654454 941935 654506 941941
rect 654454 941877 654506 941883
rect 660898 941201 660926 986499
rect 660982 986483 661034 986489
rect 660982 986425 661034 986431
rect 660994 942015 661022 986425
rect 674518 983671 674570 983677
rect 674518 983613 674570 983619
rect 674326 983597 674378 983603
rect 674326 983539 674378 983545
rect 674338 967587 674366 983539
rect 674324 967578 674380 967587
rect 674324 967513 674380 967522
rect 674530 967439 674558 983613
rect 674996 967578 675052 967587
rect 674996 967513 675052 967522
rect 674516 967430 674572 967439
rect 674516 967365 674572 967374
rect 675010 960573 675038 967513
rect 675778 966403 675806 966736
rect 675764 966394 675820 966403
rect 675764 966329 675820 966338
rect 675682 965811 675710 966070
rect 675668 965802 675724 965811
rect 675668 965737 675724 965746
rect 675202 965421 675408 965449
rect 675202 964923 675230 965421
rect 675188 964914 675244 964923
rect 675188 964849 675244 964858
rect 675778 963295 675806 963595
rect 675764 963286 675820 963295
rect 675764 963221 675820 963230
rect 675106 963022 675408 963050
rect 675106 962555 675134 963022
rect 675092 962546 675148 962555
rect 675092 962481 675148 962490
rect 675106 962385 675408 962413
rect 675106 962259 675134 962385
rect 675092 962250 675148 962259
rect 675092 962185 675148 962194
rect 675394 961519 675422 961778
rect 675380 961510 675436 961519
rect 675380 961445 675436 961454
rect 675380 961362 675436 961371
rect 675380 961297 675436 961306
rect 675394 961186 675422 961297
rect 675010 960559 675504 960573
rect 675010 960545 675518 960559
rect 675490 960187 675518 960545
rect 675476 960178 675532 960187
rect 675476 960113 675532 960122
rect 675778 959151 675806 959262
rect 675764 959142 675820 959151
rect 675764 959077 675820 959086
rect 675394 958221 675422 958744
rect 675094 958215 675146 958221
rect 675094 958157 675146 958163
rect 675382 958215 675434 958221
rect 675382 958157 675434 958163
rect 669526 954737 669578 954743
rect 669526 954679 669578 954685
rect 660982 942009 661034 942015
rect 660982 941951 661034 941957
rect 660886 941195 660938 941201
rect 660886 941137 660938 941143
rect 654452 929838 654508 929847
rect 654452 929773 654508 929782
rect 654466 927511 654494 929773
rect 654454 927505 654506 927511
rect 654454 927447 654506 927453
rect 666742 927505 666794 927511
rect 666742 927447 666794 927453
rect 653972 918146 654028 918155
rect 653972 918081 654028 918090
rect 653986 915893 654014 918081
rect 653974 915887 654026 915893
rect 653974 915829 654026 915835
rect 660982 915887 661034 915893
rect 660982 915829 661034 915835
rect 654452 906454 654508 906463
rect 654452 906389 654508 906398
rect 654466 904423 654494 906389
rect 654454 904417 654506 904423
rect 654454 904359 654506 904365
rect 653972 882922 654028 882931
rect 653972 882857 654028 882866
rect 653986 881335 654014 882857
rect 653974 881329 654026 881335
rect 653974 881271 654026 881277
rect 660886 881329 660938 881335
rect 660886 881271 660938 881277
rect 654452 871230 654508 871239
rect 654452 871165 654508 871174
rect 654466 869865 654494 871165
rect 654454 869859 654506 869865
rect 654454 869801 654506 869807
rect 654164 859538 654220 859547
rect 654164 859473 654220 859482
rect 654178 858321 654206 859473
rect 654166 858315 654218 858321
rect 654166 858257 654218 858263
rect 653972 836006 654028 836015
rect 653972 835941 654028 835950
rect 653986 835233 654014 835941
rect 653974 835227 654026 835233
rect 653974 835169 654026 835175
rect 653972 824314 654028 824323
rect 653972 824249 654028 824258
rect 653986 823763 654014 824249
rect 653974 823757 654026 823763
rect 653974 823699 654026 823705
rect 654452 812622 654508 812631
rect 654452 812557 654508 812566
rect 654466 812219 654494 812557
rect 654454 812213 654506 812219
rect 654454 812155 654506 812161
rect 654068 789090 654124 789099
rect 654068 789025 654124 789034
rect 654082 786319 654110 789025
rect 654070 786313 654122 786319
rect 654070 786255 654122 786261
rect 654068 777398 654124 777407
rect 654068 777333 654124 777342
rect 654082 774775 654110 777333
rect 654070 774769 654122 774775
rect 654070 774711 654122 774717
rect 653972 765558 654028 765567
rect 653972 765493 654028 765502
rect 653986 763305 654014 765493
rect 653974 763299 654026 763305
rect 653974 763241 654026 763247
rect 653972 742174 654028 742183
rect 653972 742109 654028 742118
rect 653986 740217 654014 742109
rect 653974 740211 654026 740217
rect 653974 740153 654026 740159
rect 655220 730482 655276 730491
rect 655220 730417 655276 730426
rect 654260 718642 654316 718651
rect 654260 718577 654316 718586
rect 654274 717203 654302 718577
rect 654262 717197 654314 717203
rect 654262 717139 654314 717145
rect 654452 695258 654508 695267
rect 654452 695193 654508 695202
rect 654466 694115 654494 695193
rect 654454 694109 654506 694115
rect 654454 694051 654506 694057
rect 654452 671726 654508 671735
rect 654452 671661 654508 671670
rect 654466 671101 654494 671661
rect 654454 671095 654506 671101
rect 654454 671037 654506 671043
rect 654260 648342 654316 648351
rect 654260 648277 654316 648286
rect 654274 648087 654302 648277
rect 654262 648081 654314 648087
rect 654262 648023 654314 648029
rect 654356 624810 654412 624819
rect 654356 624745 654412 624754
rect 654370 622113 654398 624745
rect 654358 622107 654410 622113
rect 654358 622049 654410 622055
rect 654358 613449 654410 613455
rect 654358 613391 654410 613397
rect 654370 613127 654398 613391
rect 654356 613118 654412 613127
rect 654356 613053 654412 613062
rect 654452 601426 654508 601435
rect 654452 601361 654508 601370
rect 654466 599099 654494 601361
rect 654454 599093 654506 599099
rect 654454 599035 654506 599041
rect 655124 589586 655180 589595
rect 655124 589521 655180 589530
rect 654452 577894 654508 577903
rect 654452 577829 654508 577838
rect 654466 576085 654494 577829
rect 654454 576079 654506 576085
rect 654454 576021 654506 576027
rect 654358 567347 654410 567353
rect 654358 567289 654410 567295
rect 654370 566211 654398 567289
rect 654356 566202 654412 566211
rect 654356 566137 654412 566146
rect 654452 554510 654508 554519
rect 654452 554445 654508 554454
rect 654466 552997 654494 554445
rect 654454 552991 654506 552997
rect 654454 552933 654506 552939
rect 654164 542670 654220 542679
rect 654164 542605 654220 542614
rect 654178 541601 654206 542605
rect 654166 541595 654218 541601
rect 654166 541537 654218 541543
rect 654068 530978 654124 530987
rect 654068 530913 654124 530922
rect 654082 529983 654110 530913
rect 654070 529977 654122 529983
rect 654070 529919 654122 529925
rect 654070 519395 654122 519401
rect 654070 519337 654122 519343
rect 654082 519295 654110 519337
rect 654068 519286 654124 519295
rect 654068 519221 654124 519230
rect 654260 484062 654316 484071
rect 654260 483997 654316 484006
rect 654274 483881 654302 483997
rect 654262 483875 654314 483881
rect 654262 483817 654314 483823
rect 654454 472257 654506 472263
rect 654452 472222 654454 472231
rect 654506 472222 654508 472231
rect 654452 472157 654508 472166
rect 654452 460530 654508 460539
rect 654452 460465 654508 460474
rect 654466 457981 654494 460465
rect 654454 457975 654506 457981
rect 654454 457917 654506 457923
rect 654356 448838 654412 448847
rect 654356 448773 654412 448782
rect 654370 446437 654398 448773
rect 654358 446431 654410 446437
rect 654358 446373 654410 446379
rect 654452 436998 654508 437007
rect 654452 436933 654508 436942
rect 654466 434967 654494 436933
rect 654454 434961 654506 434967
rect 654454 434903 654506 434909
rect 654454 426229 654506 426235
rect 654454 426171 654506 426177
rect 654466 425463 654494 426171
rect 654452 425454 654508 425463
rect 654452 425389 654508 425398
rect 653876 413614 653932 413623
rect 653876 413549 653932 413558
rect 653890 411879 653918 413549
rect 653878 411873 653930 411879
rect 653878 411815 653930 411821
rect 655138 409141 655166 589521
rect 655234 584817 655262 730417
rect 660898 721939 660926 881271
rect 660994 767523 661022 915829
rect 663958 904417 664010 904423
rect 663958 904359 664010 904365
rect 663766 869859 663818 869865
rect 663766 869801 663818 869807
rect 661078 858315 661130 858321
rect 661078 858257 661130 858263
rect 660982 767517 661034 767523
rect 660982 767459 661034 767465
rect 660982 737325 661034 737331
rect 660982 737267 661034 737273
rect 660886 721933 660938 721939
rect 660886 721875 660938 721881
rect 655412 683566 655468 683575
rect 655412 683501 655468 683510
rect 655316 636650 655372 636659
rect 655316 636585 655372 636594
rect 655222 584811 655274 584817
rect 655222 584753 655274 584759
rect 655220 495754 655276 495763
rect 655220 495689 655276 495698
rect 655126 409135 655178 409141
rect 655126 409077 655178 409083
rect 654452 401774 654508 401783
rect 654452 401709 654508 401718
rect 654466 400409 654494 401709
rect 654454 400403 654506 400409
rect 654454 400345 654506 400351
rect 654452 390082 654508 390091
rect 654452 390017 654508 390026
rect 654466 388865 654494 390017
rect 654454 388859 654506 388865
rect 654454 388801 654506 388807
rect 654454 380127 654506 380133
rect 654454 380069 654506 380075
rect 654466 378547 654494 380069
rect 654452 378538 654508 378547
rect 654452 378473 654508 378482
rect 654452 366550 654508 366559
rect 654452 366485 654508 366494
rect 654466 365851 654494 366485
rect 654454 365845 654506 365851
rect 654454 365787 654506 365793
rect 654452 343166 654508 343175
rect 654452 343101 654508 343110
rect 654466 342763 654494 343101
rect 654454 342757 654506 342763
rect 654454 342699 654506 342705
rect 654454 332323 654506 332329
rect 654454 332265 654506 332271
rect 654466 331631 654494 332265
rect 654452 331622 654508 331631
rect 654452 331557 654508 331566
rect 655124 319782 655180 319791
rect 655234 319749 655262 495689
rect 655330 495573 655358 636585
rect 655426 541527 655454 683501
rect 660886 555877 660938 555883
rect 660886 555819 660938 555825
rect 655414 541521 655466 541527
rect 655414 541463 655466 541469
rect 656372 507446 656428 507455
rect 656372 507381 656428 507390
rect 656386 506969 656414 507381
rect 656374 506963 656426 506969
rect 656374 506905 656426 506911
rect 655318 495567 655370 495573
rect 655318 495509 655370 495515
rect 655316 354858 655372 354867
rect 655316 354793 655372 354802
rect 655124 319717 655180 319726
rect 655222 319743 655274 319749
rect 654454 284963 654506 284969
rect 654454 284905 654506 284911
rect 654466 284715 654494 284905
rect 654452 284706 654508 284715
rect 654452 284641 654508 284650
rect 650998 237677 651050 237683
rect 650998 237619 651050 237625
rect 650518 231609 650570 231615
rect 650518 231551 650570 231557
rect 650326 231165 650378 231171
rect 650326 231107 650378 231113
rect 650038 230721 650090 230727
rect 650038 230663 650090 230669
rect 647924 210410 647980 210419
rect 647924 210345 647980 210354
rect 647938 210303 647966 210345
rect 647926 210297 647978 210303
rect 647926 210239 647978 210245
rect 647062 167229 647114 167235
rect 647062 167171 647114 167177
rect 646292 166602 646348 166611
rect 646292 166537 646348 166546
rect 646306 164275 646334 166537
rect 647074 166019 647102 167171
rect 647924 166306 647980 166315
rect 647924 166241 647980 166250
rect 647060 166010 647116 166019
rect 647060 165945 647116 165954
rect 646294 164269 646346 164275
rect 646294 164211 646346 164217
rect 647938 164201 647966 166241
rect 647926 164195 647978 164201
rect 647926 164137 647978 164143
rect 655138 138449 655166 319717
rect 655222 319685 655274 319691
rect 655220 307942 655276 307951
rect 655220 307877 655276 307886
rect 655234 138597 655262 307877
rect 655330 184403 655358 354793
rect 655412 296250 655468 296259
rect 655412 296185 655468 296194
rect 655318 184397 655370 184403
rect 655318 184339 655370 184345
rect 655222 138591 655274 138597
rect 655222 138533 655274 138539
rect 655126 138443 655178 138449
rect 655126 138385 655178 138391
rect 655426 135637 655454 296185
rect 660898 284969 660926 555819
rect 660994 472263 661022 737267
rect 661090 720903 661118 858257
rect 661174 763299 661226 763305
rect 661174 763241 661226 763247
rect 661078 720897 661130 720903
rect 661078 720839 661130 720845
rect 661078 671095 661130 671101
rect 661078 671037 661130 671043
rect 661090 540787 661118 671037
rect 661186 630697 661214 763241
rect 663778 722531 663806 869801
rect 663862 780541 663914 780547
rect 663862 780483 663914 780489
rect 663766 722525 663818 722531
rect 663766 722467 663818 722473
rect 661174 630691 661226 630697
rect 661174 630633 661226 630639
rect 663766 601979 663818 601985
rect 663766 601921 663818 601927
rect 661174 541595 661226 541601
rect 661174 541537 661226 541543
rect 661078 540781 661130 540787
rect 661078 540723 661130 540729
rect 660982 472257 661034 472263
rect 660982 472199 661034 472205
rect 661078 457975 661130 457981
rect 661078 457917 661130 457923
rect 660982 365845 661034 365851
rect 660982 365787 661034 365793
rect 660886 284963 660938 284969
rect 660886 284905 660938 284911
rect 660994 183959 661022 365787
rect 661090 274091 661118 457917
rect 661186 364963 661214 541537
rect 661174 364957 661226 364963
rect 661174 364899 661226 364905
rect 663778 332329 663806 601921
rect 663874 519401 663902 780483
rect 663970 765895 663998 904359
rect 666646 865345 666698 865351
rect 666646 865287 666698 865293
rect 664054 812213 664106 812219
rect 664054 812155 664106 812161
rect 663958 765889 664010 765895
rect 663958 765831 664010 765837
rect 663958 717197 664010 717203
rect 663958 717139 664010 717145
rect 663970 585483 663998 717139
rect 664066 675911 664094 812155
rect 664054 675905 664106 675911
rect 664054 675847 664106 675853
rect 663958 585477 664010 585483
rect 663958 585419 664010 585425
rect 666658 567353 666686 865287
rect 666754 766931 666782 927447
rect 666838 786313 666890 786319
rect 666838 786255 666890 786261
rect 666742 766925 666794 766931
rect 666742 766867 666794 766873
rect 666742 641125 666794 641131
rect 666742 641067 666794 641073
rect 666646 567347 666698 567353
rect 666646 567289 666698 567295
rect 663958 552991 664010 552997
rect 663958 552933 664010 552939
rect 663862 519395 663914 519401
rect 663862 519337 663914 519343
rect 663862 446431 663914 446437
rect 663862 446373 663914 446379
rect 663766 332323 663818 332329
rect 663766 332265 663818 332271
rect 663874 274979 663902 446373
rect 663970 363927 663998 552933
rect 664054 434961 664106 434967
rect 664054 434903 664106 434909
rect 663958 363921 664010 363927
rect 663958 363863 664010 363869
rect 663862 274973 663914 274979
rect 663862 274915 663914 274921
rect 661078 274085 661130 274091
rect 661078 274027 661130 274033
rect 664066 273351 664094 434903
rect 666646 400403 666698 400409
rect 666646 400345 666698 400351
rect 664054 273345 664106 273351
rect 664054 273287 664106 273293
rect 666658 229543 666686 400345
rect 666754 380133 666782 641067
rect 666850 631807 666878 786255
rect 666934 774769 666986 774775
rect 666934 774711 666986 774717
rect 666946 632547 666974 774711
rect 666934 632541 666986 632547
rect 666934 632483 666986 632489
rect 666838 631801 666890 631807
rect 666838 631743 666890 631749
rect 669538 613455 669566 954679
rect 673942 953997 673994 954003
rect 673942 953939 673994 953945
rect 673844 942566 673900 942575
rect 673844 942501 673900 942510
rect 673174 872893 673226 872899
rect 673174 872835 673226 872841
rect 673078 869193 673130 869199
rect 673078 869135 673130 869141
rect 669718 835227 669770 835233
rect 669718 835169 669770 835175
rect 669622 686265 669674 686271
rect 669622 686207 669674 686213
rect 669526 613449 669578 613455
rect 669526 613391 669578 613397
rect 666838 599093 666890 599099
rect 666838 599035 666890 599041
rect 666850 409215 666878 599035
rect 669526 506963 669578 506969
rect 669526 506905 669578 506911
rect 666934 483875 666986 483881
rect 666934 483817 666986 483823
rect 666838 409209 666890 409215
rect 666838 409151 666890 409157
rect 666742 380127 666794 380133
rect 666742 380069 666794 380075
rect 666742 342757 666794 342763
rect 666742 342699 666794 342705
rect 666646 229537 666698 229543
rect 666646 229479 666698 229485
rect 660982 183953 661034 183959
rect 660982 183895 661034 183901
rect 666754 182923 666782 342699
rect 666946 318343 666974 483817
rect 669538 318935 669566 506905
rect 669634 426235 669662 686207
rect 669730 676725 669758 835169
rect 672502 823757 672554 823763
rect 672502 823699 672554 823705
rect 672310 784315 672362 784321
rect 672310 784257 672362 784263
rect 671926 783501 671978 783507
rect 671926 783443 671978 783449
rect 671938 710543 671966 783443
rect 672118 763521 672170 763527
rect 672118 763463 672170 763469
rect 672022 734439 672074 734445
rect 672022 734381 672074 734387
rect 671926 710537 671978 710543
rect 671926 710479 671978 710485
rect 669814 694109 669866 694115
rect 669814 694051 669866 694057
rect 669718 676719 669770 676725
rect 669718 676661 669770 676667
rect 669718 622107 669770 622113
rect 669718 622049 669770 622055
rect 669730 496535 669758 622049
rect 669826 541453 669854 694051
rect 672034 664367 672062 734381
rect 672130 718503 672158 763463
rect 672214 760413 672266 760419
rect 672214 760355 672266 760361
rect 672116 718494 672172 718503
rect 672116 718429 672172 718438
rect 672130 681387 672158 718429
rect 672226 717055 672254 760355
rect 672214 717049 672266 717055
rect 672214 716991 672266 716997
rect 672322 711579 672350 784257
rect 672406 782539 672458 782545
rect 672406 782481 672458 782487
rect 672418 743029 672446 782481
rect 672406 743023 672458 743029
rect 672406 742965 672458 742971
rect 672406 740211 672458 740217
rect 672406 740153 672458 740159
rect 672310 711573 672362 711579
rect 672310 711515 672362 711521
rect 672310 692925 672362 692931
rect 672310 692867 672362 692873
rect 672118 681381 672170 681387
rect 672118 681323 672170 681329
rect 672022 664361 672074 664367
rect 672022 664303 672074 664309
rect 672214 648007 672266 648013
rect 672214 647949 672266 647955
rect 671926 627953 671978 627959
rect 671926 627895 671978 627901
rect 671638 602941 671690 602947
rect 671638 602883 671690 602889
rect 669814 541447 669866 541453
rect 669814 541389 669866 541395
rect 671650 528059 671678 602883
rect 671830 599315 671882 599321
rect 671830 599257 671882 599263
rect 671734 583405 671786 583411
rect 671734 583347 671786 583353
rect 671746 535607 671774 583347
rect 671734 535601 671786 535607
rect 671734 535543 671786 535549
rect 671842 528947 671870 599257
rect 671938 583411 671966 627895
rect 672022 627879 672074 627885
rect 672022 627821 672074 627827
rect 672034 586223 672062 627821
rect 672118 597169 672170 597175
rect 672118 597111 672170 597117
rect 672022 586217 672074 586223
rect 672022 586159 672074 586165
rect 671926 583405 671978 583411
rect 671926 583347 671978 583353
rect 672022 581925 672074 581931
rect 672022 581867 672074 581873
rect 671926 581851 671978 581857
rect 671926 581793 671978 581799
rect 671938 539899 671966 581793
rect 671926 539893 671978 539899
rect 671926 539835 671978 539841
rect 672034 535681 672062 581867
rect 672022 535675 672074 535681
rect 672022 535617 672074 535623
rect 672130 529539 672158 597111
rect 672226 572903 672254 647949
rect 672322 618043 672350 692867
rect 672310 618037 672362 618043
rect 672310 617979 672362 617985
rect 672310 602497 672362 602503
rect 672310 602439 672362 602445
rect 672214 572897 672266 572903
rect 672214 572839 672266 572845
rect 672322 563505 672350 602439
rect 672418 587481 672446 740153
rect 672514 677539 672542 823699
rect 672790 783131 672842 783137
rect 672790 783073 672842 783079
rect 672598 782983 672650 782989
rect 672598 782925 672650 782931
rect 672610 708471 672638 782925
rect 672694 763299 672746 763305
rect 672694 763241 672746 763247
rect 672706 720311 672734 763241
rect 672802 748801 672830 783073
rect 672886 779949 672938 779955
rect 672886 779891 672938 779897
rect 672790 748795 672842 748801
rect 672790 748737 672842 748743
rect 672790 732367 672842 732373
rect 672790 732309 672842 732315
rect 672694 720305 672746 720311
rect 672694 720247 672746 720253
rect 672694 719047 672746 719053
rect 672694 718989 672746 718995
rect 672598 708465 672650 708471
rect 672598 708407 672650 708413
rect 672502 677533 672554 677539
rect 672502 677475 672554 677481
rect 672706 676799 672734 718989
rect 672694 676793 672746 676799
rect 672694 676735 672746 676741
rect 672802 665255 672830 732309
rect 672898 707435 672926 779891
rect 672982 778617 673034 778623
rect 672982 778559 673034 778565
rect 672886 707429 672938 707435
rect 672886 707371 672938 707377
rect 672994 706843 673022 778559
rect 673090 752395 673118 869135
rect 673186 755503 673214 872835
rect 673366 872153 673418 872159
rect 673366 872095 673418 872101
rect 673270 867861 673322 867867
rect 673270 867803 673322 867809
rect 673172 755494 673228 755503
rect 673172 755429 673228 755438
rect 673076 752386 673132 752395
rect 673076 752321 673132 752330
rect 673282 751655 673310 867803
rect 673378 753283 673406 872095
rect 673858 765123 673886 942501
rect 673954 939615 673982 953939
rect 675106 953527 675134 958157
rect 675394 957819 675422 958078
rect 675380 957810 675436 957819
rect 675380 957745 675436 957754
rect 675490 957037 675518 957412
rect 675190 957031 675242 957037
rect 675190 956973 675242 956979
rect 675478 957031 675530 957037
rect 675478 956973 675530 956979
rect 675092 953518 675148 953527
rect 675092 953453 675148 953462
rect 675202 953379 675230 956973
rect 675490 956043 675518 956228
rect 675476 956034 675532 956043
rect 675476 955969 675532 955978
rect 675394 954743 675422 955044
rect 675382 954737 675434 954743
rect 675382 954679 675434 954685
rect 675490 954003 675518 954378
rect 675478 953997 675530 954003
rect 675478 953939 675530 953945
rect 675188 953370 675244 953379
rect 675188 953305 675244 953314
rect 675490 952079 675518 952528
rect 674038 952073 674090 952079
rect 674038 952015 674090 952021
rect 675478 952073 675530 952079
rect 675478 952015 675530 952021
rect 673940 939606 673996 939615
rect 673940 939541 673996 939550
rect 674050 939055 674078 952015
rect 674516 945378 674572 945387
rect 674516 945313 674572 945322
rect 674530 944901 674558 945313
rect 674518 944895 674570 944901
rect 674518 944837 674570 944843
rect 674516 944786 674572 944795
rect 674516 944721 674572 944730
rect 674530 944679 674558 944721
rect 674518 944673 674570 944679
rect 674518 944615 674570 944621
rect 674900 944046 674956 944055
rect 674900 943981 674956 943990
rect 674516 942862 674572 942871
rect 674516 942797 674572 942806
rect 674530 942089 674558 942797
rect 674518 942083 674570 942089
rect 674518 942025 674570 942031
rect 674422 942009 674474 942015
rect 674420 941974 674422 941983
rect 674474 941974 674476 941983
rect 674914 941941 674942 943981
rect 674420 941909 674476 941918
rect 674902 941935 674954 941941
rect 674902 941877 674954 941883
rect 674422 941195 674474 941201
rect 674420 941160 674422 941169
rect 674474 941160 674476 941169
rect 674420 941095 674476 941104
rect 674038 939049 674090 939055
rect 674038 938991 674090 938997
rect 676822 939049 676874 939055
rect 676822 938991 676874 938997
rect 676834 936655 676862 938991
rect 676820 936646 676876 936655
rect 676820 936581 676876 936590
rect 679796 928654 679852 928663
rect 679796 928589 679852 928598
rect 679810 928071 679838 928589
rect 679796 928062 679852 928071
rect 679796 927997 679852 928006
rect 679810 927437 679838 927997
rect 679798 927431 679850 927437
rect 679798 927373 679850 927379
rect 675778 877011 675806 877523
rect 675764 877002 675820 877011
rect 675764 876937 675820 876946
rect 675394 876567 675422 876900
rect 675380 876558 675436 876567
rect 675380 876493 675436 876502
rect 675394 875975 675422 876234
rect 675380 875966 675436 875975
rect 675380 875901 675436 875910
rect 675092 875818 675148 875827
rect 675092 875753 675148 875762
rect 675106 871715 675134 875753
rect 675188 875670 675244 875679
rect 675188 875605 675244 875614
rect 674038 871709 674090 871715
rect 674038 871651 674090 871657
rect 675094 871709 675146 871715
rect 675094 871651 675146 871657
rect 674050 789205 674078 871651
rect 675202 871493 675230 875605
rect 675490 874051 675518 874384
rect 675476 874042 675532 874051
rect 675476 873977 675532 873986
rect 675394 873459 675422 873866
rect 675380 873450 675436 873459
rect 675380 873385 675436 873394
rect 675394 872899 675422 873200
rect 675382 872893 675434 872899
rect 675382 872835 675434 872841
rect 675490 872159 675518 872534
rect 675478 872153 675530 872159
rect 675478 872095 675530 872101
rect 675394 871715 675422 872016
rect 675382 871709 675434 871715
rect 675382 871651 675434 871657
rect 674230 871487 674282 871493
rect 674230 871429 674282 871435
rect 675190 871487 675242 871493
rect 675190 871429 675242 871435
rect 675382 871487 675434 871493
rect 675382 871429 675434 871435
rect 674134 866529 674186 866535
rect 674134 866471 674186 866477
rect 674038 789199 674090 789205
rect 674038 789141 674090 789147
rect 674146 773115 674174 866471
rect 674242 782545 674270 871429
rect 675394 871350 675422 871429
rect 675394 869907 675422 870092
rect 675380 869898 675436 869907
rect 675380 869833 675436 869842
rect 675490 869199 675518 869500
rect 675478 869193 675530 869199
rect 675478 869135 675530 869141
rect 675394 868385 675422 868875
rect 674518 868379 674570 868385
rect 674518 868321 674570 868327
rect 675382 868379 675434 868385
rect 675382 868321 675434 868327
rect 674230 782539 674282 782545
rect 674230 782481 674282 782487
rect 674530 777555 674558 868321
rect 675394 867867 675422 868242
rect 675382 867861 675434 867867
rect 675382 867803 675434 867809
rect 675394 866535 675422 867058
rect 675382 866529 675434 866535
rect 675382 866471 675434 866477
rect 675394 865351 675422 865839
rect 675382 865345 675434 865351
rect 675382 865287 675434 865293
rect 675778 864727 675806 865208
rect 675764 864718 675820 864727
rect 675764 864653 675820 864662
rect 675394 862951 675422 863358
rect 675380 862942 675436 862951
rect 675380 862877 675436 862886
rect 675094 789199 675146 789205
rect 675094 789141 675146 789147
rect 675106 783137 675134 789141
rect 675682 788063 675710 788322
rect 675668 788054 675724 788063
rect 675668 787989 675724 787998
rect 675490 787175 675518 787656
rect 675476 787166 675532 787175
rect 675476 787101 675532 787110
rect 675778 786731 675806 787035
rect 675764 786722 675820 786731
rect 675764 786657 675820 786666
rect 675778 784807 675806 785214
rect 675764 784798 675820 784807
rect 675764 784733 675820 784742
rect 675490 784321 675518 784622
rect 675478 784315 675530 784321
rect 675478 784257 675530 784263
rect 675394 783507 675422 783999
rect 675382 783501 675434 783507
rect 675382 783443 675434 783449
rect 675094 783131 675146 783137
rect 675094 783073 675146 783079
rect 675394 782989 675422 783364
rect 675478 783131 675530 783137
rect 675478 783073 675530 783079
rect 675382 782983 675434 782989
rect 675382 782925 675434 782931
rect 675490 782803 675518 783073
rect 675478 782539 675530 782545
rect 675478 782481 675530 782487
rect 675490 782180 675518 782481
rect 675490 780663 675518 780848
rect 675476 780654 675532 780663
rect 675476 780589 675532 780598
rect 675094 780541 675146 780547
rect 675094 780483 675146 780489
rect 674516 777546 674572 777555
rect 674516 777481 674572 777490
rect 675106 777069 675134 780483
rect 675394 779955 675422 780330
rect 675382 779949 675434 779955
rect 675382 779891 675434 779897
rect 675778 779183 675806 779664
rect 675764 779174 675820 779183
rect 675764 779109 675820 779118
rect 675394 778623 675422 779031
rect 675382 778617 675434 778623
rect 675382 778559 675434 778565
rect 675778 777407 675806 777814
rect 675764 777398 675820 777407
rect 675764 777333 675820 777342
rect 675094 777063 675146 777069
rect 675094 777005 675146 777011
rect 675382 777063 675434 777069
rect 675382 777005 675434 777011
rect 675394 776630 675422 777005
rect 675778 775483 675806 775995
rect 675764 775474 675820 775483
rect 675764 775409 675820 775418
rect 675490 773707 675518 774155
rect 675476 773698 675532 773707
rect 675476 773633 675532 773642
rect 674132 773106 674188 773115
rect 674132 773041 674188 773050
rect 674422 767517 674474 767523
rect 674420 767482 674422 767491
rect 674474 767482 674476 767491
rect 674420 767417 674476 767426
rect 674614 766925 674666 766931
rect 674612 766890 674614 766899
rect 674666 766890 674668 766899
rect 674612 766825 674668 766834
rect 674422 765889 674474 765895
rect 674420 765854 674422 765863
rect 674474 765854 674476 765863
rect 674420 765789 674476 765798
rect 673844 765114 673900 765123
rect 673844 765049 673900 765058
rect 673844 764226 673900 764235
rect 673844 764161 673900 764170
rect 673858 763305 673886 764161
rect 674420 763560 674476 763569
rect 674420 763495 674422 763504
rect 674474 763495 674476 763504
rect 674422 763463 674474 763469
rect 673846 763299 673898 763305
rect 673846 763241 673898 763247
rect 673844 762746 673900 762755
rect 673844 762681 673900 762690
rect 673858 760419 673886 762681
rect 673846 760413 673898 760419
rect 673846 760355 673898 760361
rect 673364 753274 673420 753283
rect 673364 753209 673420 753218
rect 673268 751646 673324 751655
rect 673268 751581 673324 751590
rect 679796 750166 679852 750175
rect 679796 750101 679852 750110
rect 679810 749583 679838 750101
rect 679796 749574 679852 749583
rect 679796 749509 679852 749518
rect 679810 748875 679838 749509
rect 679798 748869 679850 748875
rect 679798 748811 679850 748817
rect 673846 748795 673898 748801
rect 673846 748737 673898 748743
rect 673858 737479 673886 748737
rect 675394 743219 675422 743330
rect 675380 743210 675436 743219
rect 675380 743145 675436 743154
rect 675094 743023 675146 743029
rect 675094 742965 675146 742971
rect 674710 738065 674762 738071
rect 674710 738007 674762 738013
rect 673846 737473 673898 737479
rect 673846 737415 673898 737421
rect 673366 734809 673418 734815
rect 673366 734751 673418 734757
rect 673174 733625 673226 733631
rect 673174 733567 673226 733573
rect 672982 706837 673034 706843
rect 672982 706779 673034 706785
rect 672982 692481 673034 692487
rect 672982 692423 673034 692429
rect 672790 665249 672842 665255
rect 672790 665191 672842 665197
rect 672994 653785 673022 692423
rect 673078 688633 673130 688639
rect 673078 688575 673130 688581
rect 672982 653779 673034 653785
rect 672982 653721 673034 653727
rect 672598 648081 672650 648087
rect 672598 648023 672650 648029
rect 672502 642309 672554 642315
rect 672502 642251 672554 642257
rect 672406 587475 672458 587481
rect 672406 587417 672458 587423
rect 672406 576079 672458 576085
rect 672406 576021 672458 576027
rect 672310 563499 672362 563505
rect 672310 563441 672362 563447
rect 672118 529533 672170 529539
rect 672118 529475 672170 529481
rect 671830 528941 671882 528947
rect 671830 528883 671882 528889
rect 671638 528053 671690 528059
rect 671638 527995 671690 528001
rect 669718 496529 669770 496535
rect 669718 496471 669770 496477
rect 669622 426229 669674 426235
rect 669622 426171 669674 426177
rect 669622 411873 669674 411879
rect 669622 411815 669674 411821
rect 669526 318929 669578 318935
rect 669526 318871 669578 318877
rect 666934 318337 666986 318343
rect 666934 318279 666986 318285
rect 669634 228951 669662 411815
rect 672418 408401 672446 576021
rect 672514 574383 672542 642251
rect 672502 574377 672554 574383
rect 672502 574319 672554 574325
rect 672502 529977 672554 529983
rect 672502 529919 672554 529925
rect 672406 408395 672458 408401
rect 672406 408337 672458 408343
rect 669718 388859 669770 388865
rect 669718 388801 669770 388807
rect 669622 228945 669674 228951
rect 669622 228887 669674 228893
rect 669730 227915 669758 388801
rect 672514 363335 672542 529919
rect 672610 497349 672638 648023
rect 672790 644603 672842 644609
rect 672790 644545 672842 644551
rect 672694 644085 672746 644091
rect 672694 644027 672746 644033
rect 672706 576011 672734 644027
rect 672694 576005 672746 576011
rect 672694 575947 672746 575953
rect 672802 572015 672830 644545
rect 672886 643419 672938 643425
rect 672886 643361 672938 643367
rect 672898 573125 672926 643361
rect 673090 616383 673118 688575
rect 673186 661375 673214 733567
rect 673268 674094 673324 674103
rect 673268 674029 673324 674038
rect 673172 661366 673228 661375
rect 673172 661301 673228 661310
rect 673282 629851 673310 674029
rect 673378 662263 673406 734751
rect 673858 702699 673886 737415
rect 674518 737325 674570 737331
rect 674518 737267 674570 737273
rect 674530 732077 674558 737267
rect 674614 736659 674666 736665
rect 674614 736601 674666 736607
rect 674518 732071 674570 732077
rect 674518 732013 674570 732019
rect 674518 730517 674570 730523
rect 674518 730459 674570 730465
rect 674230 728667 674282 728673
rect 674230 728609 674282 728615
rect 673942 717049 673994 717055
rect 673940 717014 673942 717023
rect 673994 717014 673996 717023
rect 673940 716949 673996 716958
rect 673846 702693 673898 702699
rect 673846 702635 673898 702641
rect 674038 683675 674090 683681
rect 674038 683617 674090 683623
rect 673750 681381 673802 681387
rect 673750 681323 673802 681329
rect 673762 673363 673790 681323
rect 673846 676793 673898 676799
rect 673846 676735 673898 676741
rect 673858 674843 673886 676735
rect 673844 674834 673900 674843
rect 673844 674769 673900 674778
rect 673748 673354 673804 673363
rect 673748 673289 673804 673298
rect 673364 662254 673420 662263
rect 673364 662189 673420 662198
rect 673366 648303 673418 648309
rect 673366 648245 673418 648251
rect 673268 629842 673324 629851
rect 673268 629777 673324 629786
rect 673270 627805 673322 627811
rect 673270 627747 673322 627753
rect 673076 616374 673132 616383
rect 673076 616309 673132 616318
rect 672982 604125 673034 604131
rect 672982 604067 673034 604073
rect 672886 573119 672938 573125
rect 672886 573061 672938 573067
rect 672790 572009 672842 572015
rect 672790 571951 672842 571957
rect 672994 531167 673022 604067
rect 673078 603311 673130 603317
rect 673078 603253 673130 603259
rect 672982 531161 673034 531167
rect 672982 531103 673034 531109
rect 673090 530099 673118 603253
rect 673174 598427 673226 598433
rect 673174 598369 673226 598375
rect 673076 530090 673132 530099
rect 673076 530025 673132 530034
rect 673186 526251 673214 598369
rect 673282 582343 673310 627747
rect 673268 582334 673324 582343
rect 673268 582269 673324 582278
rect 673282 581931 673310 582269
rect 673270 581925 673322 581931
rect 673270 581867 673322 581873
rect 673378 575239 673406 648245
rect 673762 628371 673790 673289
rect 674050 665255 674078 683617
rect 674242 667813 674270 728609
rect 674422 722525 674474 722531
rect 674420 722490 674422 722499
rect 674474 722490 674476 722499
rect 674420 722425 674476 722434
rect 674422 720897 674474 720903
rect 674420 720862 674422 720871
rect 674474 720862 674476 720871
rect 674420 720797 674476 720806
rect 674422 710537 674474 710543
rect 674420 710502 674422 710511
rect 674474 710502 674476 710511
rect 674420 710437 674476 710446
rect 674422 707429 674474 707435
rect 674420 707394 674422 707403
rect 674474 707394 674476 707403
rect 674420 707329 674476 707338
rect 674326 698993 674378 698999
rect 674326 698935 674378 698941
rect 674338 668627 674366 698935
rect 674422 685525 674474 685531
rect 674422 685467 674474 685473
rect 674324 668618 674380 668627
rect 674324 668553 674380 668562
rect 674228 667804 674284 667813
rect 674228 667739 674284 667748
rect 673846 665249 673898 665255
rect 673846 665191 673898 665197
rect 674038 665249 674090 665255
rect 674038 665191 674090 665197
rect 674326 665249 674378 665255
rect 674326 665191 674378 665197
rect 673858 664483 673886 665191
rect 673844 664474 673900 664483
rect 673844 664409 673900 664418
rect 673846 664361 673898 664367
rect 673846 664303 673898 664309
rect 673858 663891 673886 664303
rect 673844 663882 673900 663891
rect 673844 663817 673900 663826
rect 674230 653779 674282 653785
rect 674230 653721 674282 653727
rect 674242 647125 674270 653721
rect 674230 647119 674282 647125
rect 674230 647061 674282 647067
rect 674132 630730 674188 630739
rect 674132 630665 674134 630674
rect 674186 630665 674188 630674
rect 674134 630633 674186 630639
rect 673844 629102 673900 629111
rect 673844 629037 673900 629046
rect 673748 628362 673804 628371
rect 673748 628297 673804 628306
rect 673762 627959 673790 628297
rect 673750 627953 673802 627959
rect 673750 627895 673802 627901
rect 673858 627885 673886 629037
rect 673846 627879 673898 627885
rect 673846 627821 673898 627827
rect 674242 613381 674270 647061
rect 674338 622747 674366 665191
rect 674434 625929 674462 685467
rect 674530 671143 674558 730459
rect 674626 692339 674654 736601
rect 674722 727975 674750 738007
rect 675106 736665 675134 742965
rect 675778 742479 675806 742664
rect 675764 742470 675820 742479
rect 675764 742405 675820 742414
rect 675778 741739 675806 742035
rect 675764 741730 675820 741739
rect 675764 741665 675820 741674
rect 675476 740398 675532 740407
rect 675476 740333 675532 740342
rect 675490 740222 675518 740333
rect 675490 739371 675518 739630
rect 675476 739362 675532 739371
rect 675476 739297 675532 739306
rect 675394 738631 675422 738999
rect 675380 738622 675436 738631
rect 675380 738557 675436 738566
rect 675394 738071 675422 738372
rect 675382 738065 675434 738071
rect 675382 738007 675434 738013
rect 675490 737479 675518 737780
rect 675478 737473 675530 737479
rect 675478 737415 675530 737421
rect 675394 736665 675422 737159
rect 675094 736659 675146 736665
rect 675094 736601 675146 736607
rect 675382 736659 675434 736665
rect 675382 736601 675434 736607
rect 675490 735481 675518 735856
rect 675094 735475 675146 735481
rect 675094 735417 675146 735423
rect 675478 735475 675530 735481
rect 675478 735417 675530 735423
rect 674708 727966 674764 727975
rect 675106 727933 675134 735417
rect 675394 734815 675422 735338
rect 675382 734809 675434 734815
rect 675382 734751 675434 734757
rect 675394 734445 675422 734672
rect 675382 734439 675434 734445
rect 675382 734381 675434 734387
rect 675490 733631 675518 734006
rect 675478 733625 675530 733631
rect 675478 733567 675530 733573
rect 675490 732373 675518 732822
rect 675478 732367 675530 732373
rect 675478 732309 675530 732315
rect 675382 732071 675434 732077
rect 675382 732013 675434 732019
rect 675394 731638 675422 732013
rect 675490 730523 675518 730972
rect 675478 730517 675530 730523
rect 675478 730459 675530 730465
rect 675490 728673 675518 729155
rect 675478 728667 675530 728673
rect 675478 728609 675530 728615
rect 674708 727901 674764 727910
rect 675094 727927 675146 727933
rect 675094 727869 675146 727875
rect 675574 727927 675626 727933
rect 675574 727869 675626 727875
rect 674710 721933 674762 721939
rect 674708 721898 674710 721907
rect 674762 721898 674764 721907
rect 674708 721833 674764 721842
rect 674710 720305 674762 720311
rect 674708 720270 674710 720279
rect 674762 720270 674764 720279
rect 674708 720205 674764 720214
rect 674708 719086 674764 719095
rect 674708 719021 674710 719030
rect 674762 719021 674764 719030
rect 674710 718989 674762 718995
rect 674710 711573 674762 711579
rect 674708 711538 674710 711547
rect 674762 711538 674764 711547
rect 674708 711473 674764 711482
rect 674710 708465 674762 708471
rect 674708 708430 674710 708439
rect 674762 708430 674764 708439
rect 674708 708365 674764 708374
rect 674710 706837 674762 706843
rect 674708 706802 674710 706811
rect 674762 706802 674764 706811
rect 674708 706737 674764 706746
rect 674710 702693 674762 702699
rect 674710 702635 674762 702641
rect 674722 692487 674750 702635
rect 675586 698999 675614 727869
rect 679796 705174 679852 705183
rect 679796 705109 679852 705118
rect 679810 704591 679838 705109
rect 679796 704582 679852 704591
rect 679796 704517 679852 704526
rect 679810 702773 679838 704517
rect 679798 702767 679850 702773
rect 679798 702709 679850 702715
rect 675574 698993 675626 698999
rect 675574 698935 675626 698941
rect 675490 697931 675518 698338
rect 675476 697922 675532 697931
rect 675476 697857 675532 697866
rect 675778 697339 675806 697672
rect 675764 697330 675820 697339
rect 675764 697265 675820 697274
rect 675764 697182 675820 697191
rect 675764 697117 675820 697126
rect 675778 697035 675806 697117
rect 675682 694823 675710 695195
rect 675668 694814 675724 694823
rect 675668 694749 675724 694758
rect 675490 694379 675518 694638
rect 675476 694370 675532 694379
rect 675476 694305 675532 694314
rect 675490 693491 675518 693972
rect 675476 693482 675532 693491
rect 675476 693417 675532 693426
rect 675394 692931 675422 693380
rect 675382 692925 675434 692931
rect 675382 692867 675434 692873
rect 675490 692487 675518 692788
rect 674710 692481 674762 692487
rect 674710 692423 674762 692429
rect 675478 692481 675530 692487
rect 675478 692423 675530 692429
rect 674614 692333 674666 692339
rect 674614 692275 674666 692281
rect 675382 692333 675434 692339
rect 675382 692275 675434 692281
rect 675394 692173 675422 692275
rect 675394 692159 675792 692173
rect 675408 692145 675806 692159
rect 675778 691715 675806 692145
rect 675764 691706 675820 691715
rect 675764 691641 675820 691650
rect 675490 690711 675518 690864
rect 674806 690705 674858 690711
rect 674806 690647 674858 690653
rect 675478 690705 675530 690711
rect 675478 690647 675530 690653
rect 674710 677533 674762 677539
rect 674708 677498 674710 677507
rect 674762 677498 674764 677507
rect 674708 677433 674764 677442
rect 674708 676758 674764 676767
rect 674708 676693 674710 676702
rect 674762 676693 674764 676702
rect 674710 676661 674762 676667
rect 674818 676300 674846 690647
rect 675394 689823 675422 690346
rect 674902 689817 674954 689823
rect 674902 689759 674954 689765
rect 675382 689817 675434 689823
rect 675382 689759 675434 689765
rect 674914 687571 674942 689759
rect 675394 689199 675422 689680
rect 675380 689190 675436 689199
rect 675380 689125 675436 689134
rect 675490 688639 675518 689014
rect 675478 688633 675530 688639
rect 675478 688575 675530 688581
rect 674900 687562 674956 687571
rect 674900 687497 674956 687506
rect 675490 687381 675518 687830
rect 674902 687375 674954 687381
rect 674902 687317 674954 687323
rect 675478 687375 675530 687381
rect 675478 687317 675530 687323
rect 674914 681979 674942 687317
rect 675394 686271 675422 686646
rect 675382 686265 675434 686271
rect 675382 686207 675434 686213
rect 675490 685531 675518 685980
rect 675478 685525 675530 685531
rect 675478 685467 675530 685473
rect 675490 683681 675518 684130
rect 675478 683675 675530 683681
rect 675478 683617 675530 683623
rect 674902 681973 674954 681979
rect 674902 681915 674954 681921
rect 675478 681973 675530 681979
rect 675478 681915 675530 681921
rect 674722 676272 674846 676300
rect 674722 676059 674750 676272
rect 674710 676053 674762 676059
rect 674710 675995 674762 676001
rect 674998 676053 675050 676059
rect 674998 675995 675050 676001
rect 674710 675905 674762 675911
rect 674708 675870 674710 675879
rect 674762 675870 674764 675879
rect 674708 675805 674764 675814
rect 674708 672318 674764 672327
rect 674708 672253 674764 672262
rect 674516 671134 674572 671143
rect 674516 671069 674572 671078
rect 674614 660957 674666 660963
rect 674614 660899 674666 660905
rect 674518 632541 674570 632547
rect 674516 632506 674518 632515
rect 674570 632506 674572 632515
rect 674516 632441 674572 632450
rect 674518 631801 674570 631807
rect 674516 631766 674518 631775
rect 674570 631766 674572 631775
rect 674516 631701 674572 631710
rect 674420 625920 674476 625929
rect 674420 625855 674476 625864
rect 674626 623783 674654 660899
rect 674722 638171 674750 672253
rect 675010 660963 675038 675995
rect 674998 660957 675050 660963
rect 674998 660899 675050 660905
rect 675490 656819 675518 681915
rect 679700 660034 679756 660043
rect 679700 659969 679756 659978
rect 679714 659303 679742 659969
rect 679700 659294 679756 659303
rect 679700 659229 679756 659238
rect 674902 656813 674954 656819
rect 674902 656755 674954 656761
rect 675478 656813 675530 656819
rect 675478 656755 675530 656761
rect 674804 653670 674860 653679
rect 674804 653605 674860 653614
rect 674818 646459 674846 653605
rect 674806 646453 674858 646459
rect 674806 646395 674858 646401
rect 674818 638245 674846 646395
rect 674806 638239 674858 638245
rect 674806 638181 674858 638187
rect 674710 638165 674762 638171
rect 674710 638107 674762 638113
rect 674914 623815 674942 656755
rect 679714 656745 679742 659229
rect 679702 656739 679754 656745
rect 679702 656681 679754 656687
rect 675394 652643 675422 653124
rect 675380 652634 675436 652643
rect 675380 652569 675436 652578
rect 675490 652199 675518 652458
rect 675476 652190 675532 652199
rect 675476 652125 675532 652134
rect 675490 651459 675518 651835
rect 675476 651450 675532 651459
rect 675476 651385 675532 651394
rect 675778 649831 675806 650016
rect 675764 649822 675820 649831
rect 675764 649757 675820 649766
rect 675490 648943 675518 649424
rect 675476 648934 675532 648943
rect 675476 648869 675532 648878
rect 675394 648309 675422 648799
rect 675382 648303 675434 648309
rect 675382 648245 675434 648251
rect 675394 648013 675422 648166
rect 675382 648007 675434 648013
rect 675382 647949 675434 647955
rect 675394 647125 675422 647603
rect 675382 647119 675434 647125
rect 675382 647061 675434 647067
rect 675394 646459 675422 646982
rect 675382 646453 675434 646459
rect 675382 646395 675434 646401
rect 675778 645391 675806 645650
rect 675764 645382 675820 645391
rect 675764 645317 675820 645326
rect 675490 644609 675518 645132
rect 675478 644603 675530 644609
rect 675478 644545 675530 644551
rect 675490 644091 675518 644466
rect 675478 644085 675530 644091
rect 675478 644027 675530 644033
rect 675394 643425 675422 643831
rect 675382 643419 675434 643425
rect 675382 643361 675434 643367
rect 675490 642315 675518 642616
rect 675478 642309 675530 642315
rect 675478 642251 675530 642257
rect 675490 641131 675518 641432
rect 675478 641125 675530 641131
rect 675478 641067 675530 641073
rect 675394 640359 675422 640795
rect 675380 640350 675436 640359
rect 675380 640285 675436 640294
rect 675490 638583 675518 638955
rect 675476 638574 675532 638583
rect 675476 638509 675532 638518
rect 675574 638239 675626 638245
rect 675574 638181 675626 638187
rect 675382 638165 675434 638171
rect 675382 638107 675434 638113
rect 675394 628075 675422 638107
rect 675380 628066 675436 628075
rect 675380 628001 675436 628010
rect 675394 627811 675422 628001
rect 675382 627805 675434 627811
rect 675382 627747 675434 627753
rect 674902 623809 674954 623815
rect 674612 623774 674668 623783
rect 674902 623751 674954 623757
rect 675382 623809 675434 623815
rect 675382 623751 675434 623757
rect 674612 623709 674668 623718
rect 674324 622738 674380 622747
rect 674324 622673 674380 622682
rect 675394 620083 675422 623751
rect 675380 620074 675436 620083
rect 675380 620009 675436 620018
rect 674422 618037 674474 618043
rect 674420 618002 674422 618011
rect 674474 618002 674476 618011
rect 674420 617937 674476 617946
rect 675586 613455 675614 638181
rect 675764 638130 675820 638139
rect 675764 638065 675820 638074
rect 675778 631035 675806 638065
rect 675764 631026 675820 631035
rect 675764 630961 675820 630970
rect 675764 630878 675820 630887
rect 675764 630813 675820 630822
rect 675778 630443 675806 630813
rect 675764 630434 675820 630443
rect 675764 630369 675820 630378
rect 679700 615042 679756 615051
rect 679700 614977 679756 614986
rect 679714 614459 679742 614977
rect 679700 614450 679756 614459
rect 679700 614385 679756 614394
rect 679714 613529 679742 614385
rect 679702 613523 679754 613529
rect 679702 613465 679754 613471
rect 674998 613449 675050 613455
rect 674998 613391 675050 613397
rect 675574 613449 675626 613455
rect 675574 613391 675626 613397
rect 674230 613375 674282 613381
rect 674230 613317 674282 613323
rect 673750 603089 673802 603095
rect 673750 603031 673802 603037
rect 673558 599611 673610 599617
rect 673558 599553 673610 599559
rect 673364 575230 673420 575239
rect 673364 575165 673420 575174
rect 673570 526991 673598 599553
rect 673762 564171 673790 603031
rect 675010 602503 675038 613391
rect 675094 613375 675146 613381
rect 675094 613317 675146 613323
rect 675106 603095 675134 613317
rect 675394 607799 675422 608132
rect 675380 607790 675436 607799
rect 675380 607725 675436 607734
rect 675490 607207 675518 607466
rect 675476 607198 675532 607207
rect 675476 607133 675532 607142
rect 675682 606467 675710 606835
rect 675668 606458 675724 606467
rect 675668 606393 675724 606402
rect 675394 604839 675422 604995
rect 675380 604830 675436 604839
rect 675380 604765 675436 604774
rect 675490 604131 675518 604432
rect 675478 604125 675530 604131
rect 675478 604067 675530 604073
rect 675394 603317 675422 603799
rect 675382 603311 675434 603317
rect 675382 603253 675434 603259
rect 675094 603089 675146 603095
rect 675094 603031 675146 603037
rect 675382 603089 675434 603095
rect 675382 603031 675434 603037
rect 675394 602582 675422 603031
rect 675490 602947 675518 603174
rect 675478 602941 675530 602947
rect 675478 602883 675530 602889
rect 674998 602497 675050 602503
rect 674998 602439 675050 602445
rect 675382 602497 675434 602503
rect 675382 602439 675434 602445
rect 674422 601979 674474 601985
rect 675394 601959 675422 602439
rect 674422 601921 674474 601927
rect 674434 596879 674462 601921
rect 675490 600251 675518 600658
rect 675476 600242 675532 600251
rect 675476 600177 675532 600186
rect 675394 599617 675422 600140
rect 675382 599611 675434 599617
rect 675382 599553 675434 599559
rect 675394 599321 675422 599474
rect 675382 599315 675434 599321
rect 675382 599257 675434 599263
rect 675490 598433 675518 598808
rect 675478 598427 675530 598433
rect 675478 598369 675530 598375
rect 675490 597175 675518 597624
rect 675478 597169 675530 597175
rect 675478 597111 675530 597117
rect 674422 596873 674474 596879
rect 674422 596815 674474 596821
rect 675382 596873 675434 596879
rect 675382 596815 675434 596821
rect 675394 596440 675422 596815
rect 675490 595325 675518 595774
rect 674902 595319 674954 595325
rect 674902 595261 674954 595267
rect 675478 595319 675530 595325
rect 675478 595261 675530 595267
rect 673846 587475 673898 587481
rect 673846 587417 673898 587423
rect 673858 586339 673886 587417
rect 674612 586774 674668 586783
rect 674612 586709 674668 586718
rect 673844 586330 673900 586339
rect 673844 586265 673900 586274
rect 673846 586217 673898 586223
rect 673846 586159 673898 586165
rect 673858 584711 673886 586159
rect 674422 585477 674474 585483
rect 674420 585442 674422 585451
rect 674474 585442 674476 585451
rect 674420 585377 674476 585386
rect 674626 584817 674654 586709
rect 674614 584811 674666 584817
rect 674614 584753 674666 584759
rect 673844 584702 673900 584711
rect 673844 584637 673900 584646
rect 673844 583814 673900 583823
rect 673844 583749 673900 583758
rect 673858 581857 673886 583749
rect 674614 583405 674666 583411
rect 674612 583370 674614 583379
rect 674666 583370 674668 583379
rect 674612 583305 674668 583314
rect 673846 581851 673898 581857
rect 673846 581793 673898 581799
rect 673846 576005 673898 576011
rect 673846 575947 673898 575953
rect 673858 573611 673886 575947
rect 674422 574377 674474 574383
rect 674420 574342 674422 574351
rect 674474 574342 674476 574351
rect 674420 574277 674476 574286
rect 673844 573602 673900 573611
rect 673844 573537 673900 573546
rect 673846 573119 673898 573125
rect 673846 573061 673898 573067
rect 673858 571243 673886 573061
rect 674422 572897 674474 572903
rect 674420 572862 674422 572871
rect 674474 572862 674476 572871
rect 674420 572797 674476 572806
rect 674422 572009 674474 572015
rect 674420 571974 674422 571983
rect 674474 571974 674476 571983
rect 674420 571909 674476 571918
rect 673844 571234 673900 571243
rect 673844 571169 673900 571178
rect 674914 568727 674942 595261
rect 675778 593443 675806 593955
rect 675764 593434 675820 593443
rect 675764 593369 675820 593378
rect 679796 570198 679852 570207
rect 679796 570133 679852 570142
rect 679810 569319 679838 570133
rect 679796 569310 679852 569319
rect 679796 569245 679852 569254
rect 674900 568718 674956 568727
rect 674900 568653 674956 568662
rect 679810 567427 679838 569245
rect 679798 567421 679850 567427
rect 679798 567363 679850 567369
rect 673750 564165 673802 564171
rect 673750 564107 673802 564113
rect 675094 564165 675146 564171
rect 675094 564107 675146 564113
rect 674998 563499 675050 563505
rect 674998 563441 675050 563447
rect 674710 559577 674762 559583
rect 674710 559519 674762 559525
rect 674230 555285 674282 555291
rect 674230 555227 674282 555233
rect 673750 553213 673802 553219
rect 673750 553155 673802 553161
rect 673556 526982 673612 526991
rect 673556 526917 673612 526926
rect 673172 526242 673228 526251
rect 673172 526177 673228 526186
rect 672598 497343 672650 497349
rect 672598 497285 672650 497291
rect 673762 482295 673790 553155
rect 674038 546405 674090 546411
rect 674038 546347 674090 546353
rect 673940 541486 673996 541495
rect 673940 541421 673996 541430
rect 673954 539825 673982 541421
rect 673942 539819 673994 539825
rect 673942 539761 673994 539767
rect 674050 529983 674078 546347
rect 674242 539992 674270 555227
rect 674422 553805 674474 553811
rect 674422 553747 674474 553753
rect 674326 551955 674378 551961
rect 674326 551897 674378 551903
rect 674338 546411 674366 551897
rect 674326 546405 674378 546411
rect 674326 546347 674378 546353
rect 674324 542078 674380 542087
rect 674324 542013 674380 542022
rect 674338 541527 674366 542013
rect 674326 541521 674378 541527
rect 674434 541495 674462 553747
rect 674518 548255 674570 548261
rect 674518 548197 674570 548203
rect 674326 541463 674378 541469
rect 674420 541486 674476 541495
rect 674420 541421 674476 541430
rect 674242 539964 674366 539992
rect 674230 539819 674282 539825
rect 674230 539761 674282 539767
rect 674038 529977 674090 529983
rect 674038 529919 674090 529925
rect 674242 484663 674270 539761
rect 674338 489399 674366 539964
rect 674530 539400 674558 548197
rect 674612 541486 674668 541495
rect 674612 541421 674614 541430
rect 674666 541421 674668 541430
rect 674614 541389 674666 541395
rect 674614 540781 674666 540787
rect 674612 540746 674614 540755
rect 674666 540746 674668 540755
rect 674612 540681 674668 540690
rect 674614 539893 674666 539899
rect 674612 539858 674614 539867
rect 674666 539858 674668 539867
rect 674612 539793 674668 539802
rect 674530 539372 674654 539400
rect 674518 539301 674570 539307
rect 674518 539243 674570 539249
rect 674422 529977 674474 529983
rect 674422 529919 674474 529925
rect 674434 497497 674462 529919
rect 674422 497491 674474 497497
rect 674422 497433 674474 497439
rect 674422 497343 674474 497349
rect 674420 497308 674422 497317
rect 674474 497308 674476 497317
rect 674420 497243 674476 497252
rect 674422 496529 674474 496535
rect 674420 496494 674422 496503
rect 674474 496494 674476 496503
rect 674420 496429 674476 496438
rect 674530 491915 674558 539243
rect 674516 491906 674572 491915
rect 674516 491841 674572 491850
rect 674324 489390 674380 489399
rect 674324 489325 674380 489334
rect 674626 488807 674654 539372
rect 674722 497960 674750 559519
rect 675010 557752 675038 563441
rect 675106 557881 675134 564107
rect 675490 562511 675518 562918
rect 675476 562502 675532 562511
rect 675476 562437 675532 562446
rect 675490 562067 675518 562252
rect 675476 562058 675532 562067
rect 675476 561993 675532 562002
rect 675476 561762 675532 561771
rect 675476 561697 675532 561706
rect 675490 561660 675518 561697
rect 675394 559583 675422 559810
rect 675382 559577 675434 559583
rect 675382 559519 675434 559525
rect 675490 558811 675518 559218
rect 675476 558802 675532 558811
rect 675476 558737 675532 558746
rect 675394 558219 675422 558626
rect 675380 558210 675436 558219
rect 675380 558145 675436 558154
rect 675094 557875 675146 557881
rect 675094 557817 675146 557823
rect 675382 557875 675434 557881
rect 675382 557817 675434 557823
rect 675010 557724 675134 557752
rect 675106 557141 675134 557724
rect 675394 557403 675422 557817
rect 675778 557627 675806 557960
rect 675764 557618 675820 557627
rect 675764 557553 675820 557562
rect 675094 557135 675146 557141
rect 675094 557077 675146 557083
rect 675478 557135 675530 557141
rect 675478 557077 675530 557083
rect 675490 556776 675518 557077
rect 674998 555877 675050 555883
rect 674998 555819 675050 555825
rect 675010 551665 675038 555819
rect 675490 555291 675518 555444
rect 675478 555285 675530 555291
rect 675478 555227 675530 555233
rect 675394 554519 675422 554926
rect 675380 554510 675436 554519
rect 675380 554445 675436 554454
rect 675490 553811 675518 554260
rect 675478 553805 675530 553811
rect 675478 553747 675530 553753
rect 675394 553219 675422 553631
rect 675382 553213 675434 553219
rect 675382 553155 675434 553161
rect 675490 551961 675518 552410
rect 675478 551955 675530 551961
rect 675478 551897 675530 551903
rect 674998 551659 675050 551665
rect 674998 551601 675050 551607
rect 675382 551659 675434 551665
rect 675382 551601 675434 551607
rect 675394 551226 675422 551601
rect 675490 550111 675518 550595
rect 674998 550105 675050 550111
rect 674998 550047 675050 550053
rect 675478 550105 675530 550111
rect 675478 550047 675530 550053
rect 675010 541176 675038 550047
rect 675490 548261 675518 548755
rect 675478 548255 675530 548261
rect 675478 548197 675530 548203
rect 675010 541148 675134 541176
rect 675106 539307 675134 541148
rect 675094 539301 675146 539307
rect 675094 539243 675146 539249
rect 676724 538674 676780 538683
rect 676724 538609 676780 538618
rect 676532 537638 676588 537647
rect 676532 537573 676588 537582
rect 676546 535607 676574 537573
rect 676628 537046 676684 537055
rect 676628 536981 676684 536990
rect 676642 535681 676670 536981
rect 676630 535675 676682 535681
rect 676630 535617 676682 535623
rect 676534 535601 676586 535607
rect 676534 535543 676586 535549
rect 674806 531161 674858 531167
rect 674804 531126 674806 531135
rect 674858 531126 674860 531135
rect 674804 531061 674860 531070
rect 674806 529533 674858 529539
rect 674804 529498 674806 529507
rect 674858 529498 674860 529507
rect 674804 529433 674860 529442
rect 674806 528941 674858 528947
rect 674804 528906 674806 528915
rect 674858 528906 674860 528915
rect 674804 528841 674860 528850
rect 674806 528053 674858 528059
rect 674804 528018 674806 528027
rect 674858 528018 674860 528027
rect 674804 527953 674860 527962
rect 674722 497932 675038 497960
rect 674708 497826 674764 497835
rect 674708 497761 674764 497770
rect 674722 495573 674750 497761
rect 674902 497491 674954 497497
rect 674902 497433 674954 497439
rect 674710 495567 674762 495573
rect 674710 495509 674762 495515
rect 674612 488798 674668 488807
rect 674612 488733 674668 488742
rect 674914 485551 674942 497433
rect 675010 490287 675038 497932
rect 676546 493987 676574 535543
rect 676532 493978 676588 493987
rect 676532 493913 676588 493922
rect 674996 490278 675052 490287
rect 674996 490213 675052 490222
rect 674900 485542 674956 485551
rect 674900 485477 674956 485486
rect 674228 484654 674284 484663
rect 674228 484589 674284 484598
rect 673748 482286 673804 482295
rect 673748 482221 673804 482230
rect 676546 412143 676574 493913
rect 676642 493099 676670 535617
rect 676738 495911 676766 538609
rect 679796 524762 679852 524771
rect 679796 524697 679852 524706
rect 679810 524179 679838 524697
rect 679796 524170 679852 524179
rect 679796 524105 679852 524114
rect 679810 521325 679838 524105
rect 679798 521319 679850 521325
rect 679798 521261 679850 521267
rect 676724 495902 676780 495911
rect 676724 495837 676780 495846
rect 676724 494570 676780 494579
rect 676724 494505 676780 494514
rect 676628 493090 676684 493099
rect 676628 493025 676684 493034
rect 676532 412134 676588 412143
rect 676532 412069 676588 412078
rect 676642 411995 676670 493025
rect 676628 411986 676684 411995
rect 676628 411921 676684 411930
rect 674708 409322 674764 409331
rect 674708 409257 674764 409266
rect 674422 409209 674474 409215
rect 674422 409151 674474 409157
rect 674434 409109 674462 409151
rect 674722 409141 674750 409257
rect 674710 409135 674762 409141
rect 674420 409100 674476 409109
rect 674710 409077 674762 409083
rect 674420 409035 674476 409044
rect 674708 408434 674764 408443
rect 674708 408369 674710 408378
rect 674762 408369 674764 408378
rect 674710 408337 674762 408343
rect 676738 407703 676766 494505
rect 679796 480806 679852 480815
rect 679796 480741 679852 480750
rect 679810 480075 679838 480741
rect 679796 480066 679852 480075
rect 679796 480001 679852 480010
rect 679810 478183 679838 480001
rect 679798 478177 679850 478183
rect 679798 478119 679850 478125
rect 676724 407694 676780 407703
rect 676724 407629 676780 407638
rect 673844 406658 673900 406667
rect 673844 406593 673900 406602
rect 672502 363329 672554 363335
rect 672502 363271 672554 363277
rect 673858 362267 673886 406593
rect 674036 404290 674092 404299
rect 674036 404225 674092 404234
rect 673940 401922 673996 401931
rect 673940 401857 673996 401866
rect 673954 383167 673982 401857
rect 674050 384869 674078 404225
rect 675380 402070 675436 402079
rect 675380 402005 675436 402014
rect 675188 399406 675244 399415
rect 675188 399341 675244 399350
rect 674612 398518 674668 398527
rect 674612 398453 674668 398462
rect 674324 397926 674380 397935
rect 674324 397861 674380 397870
rect 674132 397186 674188 397195
rect 674132 397121 674188 397130
rect 674038 384863 674090 384869
rect 674038 384805 674090 384811
rect 673942 383161 673994 383167
rect 673942 383103 673994 383109
rect 674146 375767 674174 397121
rect 674338 385165 674366 397861
rect 674326 385159 674378 385165
rect 674326 385101 674378 385107
rect 674626 382501 674654 398453
rect 674900 396150 674956 396159
rect 674900 396085 674956 396094
rect 674708 393782 674764 393791
rect 674708 393717 674764 393726
rect 674614 382495 674666 382501
rect 674614 382437 674666 382443
rect 674722 376877 674750 393717
rect 674914 377617 674942 396085
rect 675092 395410 675148 395419
rect 675092 395345 675148 395354
rect 674996 394522 675052 394531
rect 674996 394457 675052 394466
rect 675010 378209 675038 394457
rect 675106 381336 675134 395345
rect 675202 385461 675230 399341
rect 675394 386423 675422 402005
rect 679700 392598 679756 392607
rect 679700 392533 679756 392542
rect 679714 392163 679742 392533
rect 679700 392154 679756 392163
rect 679700 392089 679756 392098
rect 679714 391751 679742 392089
rect 679702 391745 679754 391751
rect 679702 391687 679754 391693
rect 675382 386417 675434 386423
rect 675382 386359 675434 386365
rect 675382 386195 675434 386201
rect 675382 386137 675434 386143
rect 675394 385723 675422 386137
rect 675190 385455 675242 385461
rect 675190 385397 675242 385403
rect 675478 385455 675530 385461
rect 675478 385397 675530 385403
rect 675190 385159 675242 385165
rect 675190 385101 675242 385107
rect 675202 381410 675230 385101
rect 675490 385096 675518 385397
rect 675382 384863 675434 384869
rect 675382 384805 675434 384811
rect 675394 384430 675422 384805
rect 675286 383161 675338 383167
rect 675286 383103 675338 383109
rect 675298 382668 675326 383103
rect 675298 382640 675422 382668
rect 675394 382580 675422 382640
rect 675478 382495 675530 382501
rect 675478 382437 675530 382443
rect 675490 382062 675518 382437
rect 675202 381382 675408 381410
rect 675106 381308 675422 381336
rect 675394 380730 675422 381308
rect 675106 380198 675408 380226
rect 675106 379116 675134 380198
rect 675298 379532 675408 379560
rect 675106 379088 675230 379116
rect 675094 379017 675146 379023
rect 675094 378959 675146 378965
rect 674998 378203 675050 378209
rect 674998 378145 675050 378151
rect 674902 377611 674954 377617
rect 674902 377553 674954 377559
rect 674710 376871 674762 376877
rect 674710 376813 674762 376819
rect 674134 375761 674186 375767
rect 674134 375703 674186 375709
rect 675106 374107 675134 378959
rect 675202 374551 675230 379088
rect 675298 379023 675326 379532
rect 675286 379017 675338 379023
rect 675286 378959 675338 378965
rect 675476 378834 675532 378843
rect 675476 378769 675532 378778
rect 675490 378288 675518 378769
rect 675382 378203 675434 378209
rect 675382 378145 675434 378151
rect 675394 377696 675422 378145
rect 675382 377611 675434 377617
rect 675382 377553 675434 377559
rect 675394 377075 675422 377553
rect 675478 376871 675530 376877
rect 675478 376813 675530 376819
rect 675490 376438 675518 376813
rect 675478 375761 675530 375767
rect 675478 375703 675530 375709
rect 675490 375254 675518 375703
rect 675188 374542 675244 374551
rect 675188 374477 675244 374486
rect 675092 374098 675148 374107
rect 675092 374033 675148 374042
rect 675476 373950 675532 373959
rect 675476 373885 675532 373894
rect 675490 373404 675518 373885
rect 675380 372026 675436 372035
rect 675380 371961 675436 371970
rect 675394 371554 675422 371961
rect 674710 364957 674762 364963
rect 674708 364922 674710 364931
rect 674762 364922 674764 364931
rect 674708 364857 674764 364866
rect 674422 363921 674474 363927
rect 674420 363886 674422 363895
rect 674474 363886 674476 363895
rect 674420 363821 674476 363830
rect 674710 363329 674762 363335
rect 674708 363294 674710 363303
rect 674762 363294 674764 363303
rect 674708 363229 674764 363238
rect 673844 362258 673900 362267
rect 673844 362193 673900 362202
rect 673940 359150 673996 359159
rect 673940 359085 673996 359094
rect 673954 339581 673982 359085
rect 677108 358114 677164 358123
rect 677108 358049 677164 358058
rect 674612 357226 674668 357235
rect 674612 357161 674668 357170
rect 674324 352786 674380 352795
rect 674324 352721 674380 352730
rect 674228 351306 674284 351315
rect 674228 351241 674284 351250
rect 674036 349530 674092 349539
rect 674036 349465 674092 349474
rect 673942 339575 673994 339581
rect 673942 339517 673994 339523
rect 674050 332773 674078 349465
rect 674132 348790 674188 348799
rect 674132 348725 674188 348734
rect 674038 332767 674090 332773
rect 674038 332709 674090 332715
rect 674146 331589 674174 348725
rect 674242 332403 674270 351241
rect 674338 336621 674366 352721
rect 674626 340987 674654 357161
rect 675188 356486 675244 356495
rect 675188 356421 675244 356430
rect 675092 353378 675148 353387
rect 675092 353313 675148 353322
rect 674804 350270 674860 350279
rect 674804 350205 674860 350214
rect 674710 344459 674762 344465
rect 674710 344401 674762 344407
rect 674614 340981 674666 340987
rect 674614 340923 674666 340929
rect 674326 336615 674378 336621
rect 674326 336557 674378 336563
rect 674230 332397 674282 332403
rect 674230 332339 674282 332345
rect 674134 331583 674186 331589
rect 674134 331525 674186 331531
rect 674722 330553 674750 344401
rect 674818 335569 674846 350205
rect 675106 336862 675134 353313
rect 675202 337409 675230 356421
rect 676916 355746 676972 355755
rect 676916 355681 676972 355690
rect 675284 354118 675340 354127
rect 675284 354053 675340 354062
rect 675298 339896 675326 354053
rect 676820 351750 676876 351759
rect 676820 351685 676876 351694
rect 676834 344465 676862 351685
rect 676930 345395 676958 355681
rect 677012 355006 677068 355015
rect 677012 354941 677068 354950
rect 676916 345386 676972 345395
rect 676916 345321 676972 345330
rect 677026 345247 677054 354941
rect 677122 345543 677150 358049
rect 679796 347458 679852 347467
rect 679796 347393 679852 347402
rect 679810 346727 679838 347393
rect 679796 346718 679852 346727
rect 679796 346653 679852 346662
rect 679810 345649 679838 346653
rect 679798 345643 679850 345649
rect 679798 345585 679850 345591
rect 677108 345534 677164 345543
rect 677108 345469 677164 345478
rect 677012 345238 677068 345247
rect 677012 345173 677068 345182
rect 676822 344459 676874 344465
rect 676822 344401 676874 344407
rect 675478 340981 675530 340987
rect 675478 340923 675530 340929
rect 675490 340548 675518 340923
rect 675298 339868 675408 339896
rect 675382 339575 675434 339581
rect 675382 339517 675434 339523
rect 675394 339216 675422 339517
rect 675202 337381 675408 337409
rect 675106 336834 675408 336862
rect 675382 336615 675434 336621
rect 675382 336557 675434 336563
rect 675394 336182 675422 336557
rect 674818 335541 675408 335569
rect 675476 335174 675532 335183
rect 675476 335109 675532 335118
rect 675490 335012 675518 335109
rect 675202 334998 675518 335012
rect 675202 334984 675504 334998
rect 674710 330547 674762 330553
rect 674710 330489 674762 330495
rect 675202 329559 675230 334984
rect 675490 333851 675518 334332
rect 675476 333842 675532 333851
rect 675476 333777 675532 333786
rect 675764 333546 675820 333555
rect 675764 333481 675820 333490
rect 675778 333074 675806 333481
rect 675382 332767 675434 332773
rect 675382 332709 675434 332715
rect 675394 332519 675422 332709
rect 675478 332397 675530 332403
rect 675478 332339 675530 332345
rect 675490 331890 675518 332339
rect 675382 331583 675434 331589
rect 675382 331525 675434 331531
rect 675394 331224 675422 331525
rect 675478 330547 675530 330553
rect 675478 330489 675530 330495
rect 675490 330040 675518 330489
rect 675188 329550 675244 329559
rect 675188 329485 675244 329494
rect 675778 328079 675806 328190
rect 675764 328070 675820 328079
rect 675764 328005 675820 328014
rect 675764 326886 675820 326895
rect 675764 326821 675820 326830
rect 675778 326340 675806 326821
rect 674422 319743 674474 319749
rect 674420 319708 674422 319717
rect 674474 319708 674476 319717
rect 674420 319643 674476 319652
rect 674422 318929 674474 318935
rect 674420 318894 674422 318903
rect 674474 318894 674476 318903
rect 674420 318829 674476 318838
rect 674710 318337 674762 318343
rect 674708 318302 674710 318311
rect 674762 318302 674764 318311
rect 674708 318237 674764 318246
rect 674036 314158 674092 314167
rect 674036 314093 674092 314102
rect 673940 311642 673996 311651
rect 673940 311577 673996 311586
rect 673954 292961 673982 311577
rect 674050 294811 674078 314093
rect 675092 312234 675148 312243
rect 675092 312169 675148 312178
rect 674900 309126 674956 309135
rect 674900 309061 674956 309070
rect 674228 308534 674284 308543
rect 674228 308469 674284 308478
rect 674132 303798 674188 303807
rect 674132 303733 674188 303742
rect 674038 294805 674090 294811
rect 674038 294747 674090 294753
rect 673942 292955 673994 292961
rect 673942 292897 673994 292903
rect 674146 286597 674174 303733
rect 674242 294293 674270 308469
rect 674612 307498 674668 307507
rect 674612 307433 674668 307442
rect 674324 305426 674380 305435
rect 674324 305361 674380 305370
rect 674230 294287 674282 294293
rect 674230 294229 674282 294235
rect 674338 291111 674366 305361
rect 674420 304612 674476 304621
rect 674420 304547 674476 304556
rect 674326 291105 674378 291111
rect 674326 291047 674378 291053
rect 674434 287781 674462 304547
rect 674626 291777 674654 307433
rect 674710 299541 674762 299547
rect 674710 299483 674762 299489
rect 674614 291771 674666 291777
rect 674614 291713 674666 291719
rect 674422 287775 674474 287781
rect 674422 287717 674474 287723
rect 674722 287411 674750 299483
rect 674806 299467 674858 299473
rect 674806 299409 674858 299415
rect 674818 288595 674846 299409
rect 674914 294904 674942 309061
rect 675106 295537 675134 312169
rect 676916 310754 676972 310763
rect 676916 310689 676972 310698
rect 676820 306018 676876 306027
rect 676820 305953 676876 305962
rect 676834 299547 676862 305953
rect 676822 299541 676874 299547
rect 676822 299483 676874 299489
rect 676930 299473 676958 310689
rect 677108 310014 677164 310023
rect 677108 309949 677164 309958
rect 677012 306758 677068 306767
rect 677012 306693 677068 306702
rect 677026 299515 677054 306693
rect 677012 299506 677068 299515
rect 676918 299467 676970 299473
rect 677012 299441 677068 299450
rect 676918 299409 676970 299415
rect 677122 299367 677150 309949
rect 679796 302466 679852 302475
rect 679796 302401 679852 302410
rect 679810 301735 679838 302401
rect 679796 301726 679852 301735
rect 679796 301661 679852 301670
rect 679810 299621 679838 301661
rect 679798 299615 679850 299621
rect 679798 299557 679850 299563
rect 677108 299358 677164 299367
rect 677108 299293 677164 299302
rect 675106 295509 675408 295537
rect 674914 294876 675408 294904
rect 675190 294805 675242 294811
rect 675190 294747 675242 294753
rect 675094 294287 675146 294293
rect 675094 294229 675146 294235
rect 675202 294238 675230 294747
rect 675106 291870 675134 294229
rect 675202 294210 675408 294238
rect 675382 292955 675434 292961
rect 675382 292897 675434 292903
rect 675394 292374 675422 292897
rect 675106 291842 675408 291870
rect 675094 291771 675146 291777
rect 675094 291713 675146 291719
rect 675106 291204 675134 291713
rect 675106 291176 675408 291204
rect 675094 291105 675146 291111
rect 675094 291047 675146 291053
rect 675106 290569 675134 291047
rect 675106 290541 675408 290569
rect 675490 289747 675518 290006
rect 675476 289738 675532 289747
rect 675476 289673 675532 289682
rect 675380 289590 675436 289599
rect 675380 289525 675436 289534
rect 675394 289354 675422 289525
rect 675394 289340 675504 289354
rect 675408 289326 675518 289340
rect 675490 288836 675518 289326
rect 675202 288808 675518 288836
rect 674806 288589 674858 288595
rect 674806 288531 674858 288537
rect 674710 287405 674762 287411
rect 674710 287347 674762 287353
rect 674134 286591 674186 286597
rect 674134 286533 674186 286539
rect 675202 285011 675230 288808
rect 675478 288589 675530 288595
rect 675478 288531 675530 288537
rect 675490 288082 675518 288531
rect 675382 287775 675434 287781
rect 675382 287717 675434 287723
rect 675394 287519 675422 287717
rect 675478 287405 675530 287411
rect 675478 287347 675530 287353
rect 675490 286898 675518 287347
rect 675382 286591 675434 286597
rect 675382 286533 675434 286539
rect 675394 286232 675422 286533
rect 675188 285002 675244 285011
rect 675188 284937 675244 284946
rect 675778 284863 675806 285048
rect 675764 284854 675820 284863
rect 675764 284789 675820 284798
rect 675380 283670 675436 283679
rect 675380 283605 675436 283614
rect 675394 283198 675422 283605
rect 675764 281894 675820 281903
rect 675764 281829 675820 281838
rect 675778 281348 675806 281829
rect 674710 274973 674762 274979
rect 674708 274938 674710 274947
rect 674762 274938 674764 274947
rect 674708 274873 674764 274882
rect 674710 274085 674762 274091
rect 674708 274050 674710 274059
rect 674762 274050 674764 274059
rect 674708 273985 674764 273994
rect 674710 273345 674762 273351
rect 674708 273310 674710 273319
rect 674762 273310 674764 273319
rect 674708 273245 674764 273254
rect 674132 269166 674188 269175
rect 674132 269101 674188 269110
rect 673940 266650 673996 266659
rect 673940 266585 673996 266594
rect 673954 247969 673982 266585
rect 674036 263542 674092 263551
rect 674036 263477 674092 263486
rect 673942 247963 673994 247969
rect 673942 247905 673994 247911
rect 674050 247303 674078 263477
rect 674146 249597 674174 269101
rect 674516 267242 674572 267251
rect 674516 267177 674572 267186
rect 674324 262802 674380 262811
rect 674324 262737 674380 262746
rect 674228 258806 674284 258815
rect 674228 258741 674284 258750
rect 674134 249591 674186 249597
rect 674134 249533 674186 249539
rect 674038 247297 674090 247303
rect 674038 247239 674090 247245
rect 673364 244746 673420 244755
rect 673364 244681 673420 244690
rect 673378 242091 673406 244681
rect 673844 244598 673900 244607
rect 673844 244533 673900 244542
rect 673858 242239 673886 244533
rect 673844 242230 673900 242239
rect 673844 242165 673900 242174
rect 673364 242082 673420 242091
rect 673364 242017 673420 242026
rect 669718 227909 669770 227915
rect 669718 227851 669770 227857
rect 673378 225843 673406 242017
rect 673366 225837 673418 225843
rect 673366 225779 673418 225785
rect 673858 224775 673886 242165
rect 674242 241605 674270 258741
rect 674338 246785 674366 262737
rect 674530 251003 674558 267177
rect 678164 265022 678220 265031
rect 678164 264957 678220 264966
rect 674612 264134 674668 264143
rect 674612 264069 674668 264078
rect 674518 250997 674570 251003
rect 674518 250939 674570 250945
rect 674626 250411 674654 264069
rect 676916 261766 676972 261775
rect 676916 261701 676972 261710
rect 676820 261026 676876 261035
rect 676820 260961 676876 260970
rect 675284 260138 675340 260147
rect 675284 260073 675340 260082
rect 675188 259398 675244 259407
rect 675188 259333 675244 259342
rect 674998 251663 675050 251669
rect 674998 251605 675050 251611
rect 674614 250405 674666 250411
rect 674614 250347 674666 250353
rect 674326 246779 674378 246785
rect 674326 246721 674378 246727
rect 674804 245930 674860 245939
rect 674804 245865 674860 245874
rect 674818 244343 674846 245865
rect 674900 245190 674956 245199
rect 674900 245125 674956 245134
rect 674914 244903 674942 245125
rect 674900 244894 674956 244903
rect 674900 244829 674956 244838
rect 674806 244337 674858 244343
rect 674806 244279 674858 244285
rect 674230 241599 674282 241605
rect 674230 241541 674282 241547
rect 674818 238983 674846 244279
rect 674914 241943 674942 244829
rect 674900 241934 674956 241943
rect 674900 241869 674956 241878
rect 675010 240569 675038 251605
rect 675094 251589 675146 251595
rect 675094 251531 675146 251537
rect 675106 242419 675134 251531
rect 675202 243011 675230 259333
rect 675298 246064 675326 260073
rect 676834 251595 676862 260961
rect 676930 251669 676958 261701
rect 678178 253487 678206 264957
rect 679796 257474 679852 257483
rect 679796 257409 679852 257418
rect 679810 256891 679838 257409
rect 679796 256882 679852 256891
rect 679796 256817 679852 256826
rect 679810 256405 679838 256817
rect 679798 256399 679850 256405
rect 679798 256341 679850 256347
rect 678164 253478 678220 253487
rect 678164 253413 678220 253422
rect 676918 251663 676970 251669
rect 676918 251605 676970 251611
rect 676822 251589 676874 251595
rect 676822 251531 676874 251537
rect 675382 250997 675434 251003
rect 675382 250939 675434 250945
rect 675394 250523 675422 250939
rect 675478 250405 675530 250411
rect 675478 250347 675530 250353
rect 675490 249898 675518 250347
rect 675382 249591 675434 249597
rect 675382 249533 675434 249539
rect 675394 249232 675422 249533
rect 675382 247963 675434 247969
rect 675382 247905 675434 247911
rect 675394 247382 675422 247905
rect 675478 247297 675530 247303
rect 675478 247239 675530 247245
rect 675490 246864 675518 247239
rect 675382 246779 675434 246785
rect 675382 246721 675434 246727
rect 675394 246198 675422 246721
rect 675298 246036 675422 246064
rect 675394 245532 675422 246036
rect 675476 245190 675532 245199
rect 675476 245125 675532 245134
rect 675490 245014 675518 245125
rect 675298 244343 675408 244362
rect 675286 244337 675408 244343
rect 675338 244334 675408 244337
rect 675286 244279 675338 244285
rect 675476 243562 675532 243571
rect 675476 243497 675532 243506
rect 675490 243090 675518 243497
rect 675190 243005 675242 243011
rect 675190 242947 675242 242953
rect 675382 243005 675434 243011
rect 675382 242947 675434 242953
rect 675394 242498 675422 242947
rect 675094 242413 675146 242419
rect 675094 242355 675146 242361
rect 675382 242413 675434 242419
rect 675382 242355 675434 242361
rect 675394 241875 675422 242355
rect 675478 241599 675530 241605
rect 675478 241541 675530 241547
rect 675490 241240 675518 241541
rect 674998 240563 675050 240569
rect 674998 240505 675050 240511
rect 675478 240563 675530 240569
rect 675478 240505 675530 240511
rect 675490 240056 675518 240505
rect 674804 238974 674860 238983
rect 674804 238909 674860 238918
rect 675476 238678 675532 238687
rect 675476 238613 675532 238622
rect 675490 238206 675518 238613
rect 675764 236902 675820 236911
rect 675764 236837 675820 236846
rect 675778 236356 675806 236837
rect 674422 229537 674474 229543
rect 674420 229502 674422 229511
rect 674474 229502 674476 229511
rect 674420 229437 674476 229446
rect 674710 228945 674762 228951
rect 674708 228910 674710 228919
rect 674762 228910 674764 228919
rect 674708 228845 674764 228854
rect 674422 227909 674474 227915
rect 674420 227874 674422 227883
rect 674474 227874 674476 227883
rect 674420 227809 674476 227818
rect 674710 225837 674762 225843
rect 674708 225802 674710 225811
rect 679798 225837 679850 225843
rect 674762 225802 674764 225811
rect 679798 225779 679850 225785
rect 674708 225737 674764 225746
rect 673844 224766 673900 224775
rect 673844 224701 673846 224710
rect 673898 224701 673900 224710
rect 673846 224669 673898 224675
rect 673858 224641 673886 224669
rect 673940 223878 673996 223887
rect 673940 223813 673996 223822
rect 673954 204457 673982 223813
rect 674420 222250 674476 222259
rect 674420 222185 674476 222194
rect 674036 217514 674092 217523
rect 674036 217449 674092 217458
rect 673942 204451 673994 204457
rect 673942 204393 673994 204399
rect 674050 201349 674078 217449
rect 674434 205789 674462 222185
rect 674996 221214 675052 221223
rect 674996 221149 675052 221158
rect 674900 214702 674956 214711
rect 674900 214637 674956 214646
rect 674804 214258 674860 214267
rect 674804 214193 674860 214202
rect 674708 213370 674764 213379
rect 674708 213305 674764 213314
rect 674614 207411 674666 207417
rect 674614 207353 674666 207359
rect 674422 205783 674474 205789
rect 674422 205725 674474 205731
rect 674038 201343 674090 201349
rect 674038 201285 674090 201291
rect 674626 197057 674654 207353
rect 674614 197051 674666 197057
rect 674614 196993 674666 196999
rect 674722 196613 674750 213305
rect 674818 197649 674846 214193
rect 674914 200905 674942 214637
rect 675010 202237 675038 221149
rect 677012 220622 677068 220631
rect 677012 220557 677068 220566
rect 675188 218994 675244 219003
rect 675188 218929 675244 218938
rect 675092 217810 675148 217819
rect 675092 217745 675148 217754
rect 674998 202231 675050 202237
rect 674998 202173 675050 202179
rect 675106 202089 675134 217745
rect 675202 205197 675230 218929
rect 676916 216478 676972 216487
rect 676916 216413 676972 216422
rect 676820 215886 676876 215895
rect 676820 215821 676876 215830
rect 676834 207417 676862 215821
rect 676930 207459 676958 216413
rect 677026 207755 677054 220557
rect 677108 219734 677164 219743
rect 677108 219669 677164 219678
rect 677012 207746 677068 207755
rect 677012 207681 677068 207690
rect 677122 207607 677150 219669
rect 679810 212301 679838 225779
rect 679990 224727 680042 224733
rect 679990 224669 680042 224675
rect 679798 212295 679850 212301
rect 679798 212237 679850 212243
rect 679796 212186 679852 212195
rect 679796 212121 679852 212130
rect 679810 211455 679838 212121
rect 679796 211446 679852 211455
rect 679796 211381 679852 211390
rect 679810 210303 679838 211381
rect 679798 210297 679850 210303
rect 679798 210239 679850 210245
rect 680002 210123 680030 224669
rect 680086 212295 680138 212301
rect 680086 212237 680138 212243
rect 680098 210271 680126 212237
rect 680084 210262 680140 210271
rect 680084 210197 680140 210206
rect 679988 210114 680044 210123
rect 679988 210049 680044 210058
rect 677108 207598 677164 207607
rect 677108 207533 677164 207542
rect 676916 207450 676972 207459
rect 676822 207411 676874 207417
rect 676916 207385 676972 207394
rect 676822 207353 676874 207359
rect 675478 205783 675530 205789
rect 675478 205725 675530 205731
rect 675490 205350 675518 205725
rect 675190 205191 675242 205197
rect 675190 205133 675242 205139
rect 675478 205191 675530 205197
rect 675478 205133 675530 205139
rect 675490 204684 675518 205133
rect 675382 204451 675434 204457
rect 675382 204393 675434 204399
rect 675394 204018 675422 204393
rect 675298 202237 675422 202256
rect 675286 202231 675422 202237
rect 675338 202228 675422 202231
rect 675286 202173 675338 202179
rect 675394 202168 675422 202228
rect 675094 202083 675146 202089
rect 675094 202025 675146 202031
rect 675286 202083 675338 202089
rect 675286 202025 675338 202031
rect 675298 201664 675326 202025
rect 675298 201636 675408 201664
rect 675382 201343 675434 201349
rect 675382 201285 675434 201291
rect 675394 200984 675422 201285
rect 674902 200899 674954 200905
rect 674902 200841 674954 200847
rect 675382 200899 675434 200905
rect 675382 200841 675434 200847
rect 675394 200355 675422 200841
rect 675394 199319 675422 199800
rect 675380 199310 675436 199319
rect 675380 199245 675436 199254
rect 675490 198727 675518 199134
rect 675476 198718 675532 198727
rect 675476 198653 675532 198662
rect 675764 198422 675820 198431
rect 675764 198357 675820 198366
rect 675778 197876 675806 198357
rect 674806 197643 674858 197649
rect 674806 197585 674858 197591
rect 675382 197643 675434 197649
rect 675382 197585 675434 197591
rect 675394 197319 675422 197585
rect 675478 197051 675530 197057
rect 675478 196993 675530 196999
rect 675490 196692 675518 196993
rect 674710 196607 674762 196613
rect 674710 196549 674762 196555
rect 675382 196607 675434 196613
rect 675382 196549 675434 196555
rect 675394 196026 675422 196549
rect 675764 195314 675820 195323
rect 675764 195249 675820 195258
rect 675778 194842 675806 195249
rect 675380 193538 675436 193547
rect 675380 193473 675436 193482
rect 675394 192992 675422 193473
rect 675764 191614 675820 191623
rect 675764 191549 675820 191558
rect 675778 191142 675806 191549
rect 674420 184510 674476 184519
rect 674420 184445 674476 184454
rect 674434 184403 674462 184445
rect 674422 184397 674474 184403
rect 674422 184339 674474 184345
rect 674710 183953 674762 183959
rect 674708 183918 674710 183927
rect 674762 183918 674764 183927
rect 674708 183853 674764 183862
rect 666742 182917 666794 182923
rect 674422 182917 674474 182923
rect 666742 182859 666794 182865
rect 674420 182882 674422 182891
rect 674474 182882 674476 182891
rect 674420 182817 674476 182826
rect 679700 179922 679756 179931
rect 679700 179857 679756 179866
rect 674900 177110 674956 177119
rect 674900 177045 674956 177054
rect 674804 173114 674860 173123
rect 674804 173049 674860 173058
rect 674516 172374 674572 172383
rect 674516 172309 674572 172318
rect 674228 169414 674284 169423
rect 674228 169349 674284 169358
rect 674132 168526 674188 168535
rect 674132 168461 674188 168470
rect 674146 151473 674174 168461
rect 674242 152657 674270 169349
rect 674530 157763 674558 172309
rect 674708 167342 674764 167351
rect 674708 167277 674764 167286
rect 674722 167235 674750 167277
rect 674710 167229 674762 167235
rect 674710 167171 674762 167177
rect 674612 166602 674668 166611
rect 674612 166537 674668 166546
rect 674626 164275 674654 166537
rect 674708 165714 674764 165723
rect 674708 165649 674764 165658
rect 674614 164269 674666 164275
rect 674614 164211 674666 164217
rect 674722 164201 674750 165649
rect 674710 164195 674762 164201
rect 674710 164137 674762 164143
rect 674818 163776 674846 173049
rect 674626 163748 674846 163776
rect 674518 157757 674570 157763
rect 674518 157699 674570 157705
rect 674626 156949 674654 163748
rect 674710 163677 674762 163683
rect 674710 163619 674762 163625
rect 674614 156943 674666 156949
rect 674614 156885 674666 156891
rect 674230 152651 674282 152657
rect 674230 152593 674282 152599
rect 674134 151467 674186 151473
rect 674134 151409 674186 151415
rect 674722 150363 674750 163619
rect 674806 163307 674858 163313
rect 674806 163249 674858 163255
rect 674818 152213 674846 163249
rect 674914 160797 674942 177045
rect 677012 176222 677068 176231
rect 677012 176157 677068 176166
rect 676916 175630 676972 175639
rect 676916 175565 676972 175574
rect 674996 174002 675052 174011
rect 674996 173937 675052 173946
rect 674902 160791 674954 160797
rect 674902 160733 674954 160739
rect 675010 160057 675038 173937
rect 676820 170894 676876 170903
rect 676820 170829 676876 170838
rect 675092 170006 675148 170015
rect 675092 169941 675148 169950
rect 674998 160051 675050 160057
rect 674998 159993 675050 159999
rect 675106 155369 675134 169941
rect 675764 166454 675820 166463
rect 675764 166389 675820 166398
rect 675778 165575 675806 166389
rect 675764 165566 675820 165575
rect 675764 165501 675820 165510
rect 676834 163313 676862 170829
rect 676822 163307 676874 163313
rect 676822 163249 676874 163255
rect 676930 162911 676958 175565
rect 676916 162902 676972 162911
rect 676916 162837 676972 162846
rect 677026 161431 677054 176157
rect 677204 174742 677260 174751
rect 677204 174677 677260 174686
rect 677108 171486 677164 171495
rect 677108 171421 677164 171430
rect 677122 163683 677150 171421
rect 677218 164095 677246 174677
rect 679714 166611 679742 179857
rect 679796 179478 679852 179487
rect 679796 179413 679852 179422
rect 679700 166602 679756 166611
rect 679700 166537 679756 166546
rect 679810 166463 679838 179413
rect 679796 166454 679852 166463
rect 679796 166389 679852 166398
rect 677204 164086 677260 164095
rect 677204 164021 677260 164030
rect 677110 163677 677162 163683
rect 677110 163619 677162 163625
rect 677012 161422 677068 161431
rect 677012 161357 677068 161366
rect 675382 160791 675434 160797
rect 675382 160733 675434 160739
rect 675394 160323 675422 160733
rect 675478 160051 675530 160057
rect 675478 159993 675530 159999
rect 675490 159692 675518 159993
rect 675380 159350 675436 159359
rect 675380 159285 675436 159294
rect 675394 159026 675422 159285
rect 675190 157757 675242 157763
rect 675190 157699 675242 157705
rect 675764 157722 675820 157731
rect 675202 156006 675230 157699
rect 675764 157657 675820 157666
rect 675778 157176 675806 157657
rect 675478 156943 675530 156949
rect 675478 156885 675530 156891
rect 675490 156658 675518 156885
rect 675202 155978 675408 156006
rect 675106 155341 675408 155369
rect 675394 154623 675422 154808
rect 675380 154614 675436 154623
rect 675380 154549 675436 154558
rect 675380 154318 675436 154327
rect 675298 154276 675380 154304
rect 675298 154156 675326 154276
rect 675380 154253 675436 154262
rect 675202 154128 675326 154156
rect 675394 154142 675422 154253
rect 674806 152207 674858 152213
rect 674806 152149 674858 152155
rect 674710 150357 674762 150363
rect 674710 150299 674762 150305
rect 675202 148407 675230 154128
rect 675764 153430 675820 153439
rect 675764 153365 675820 153374
rect 675778 152884 675806 153365
rect 675382 152651 675434 152657
rect 675382 152593 675434 152599
rect 675394 152292 675422 152593
rect 675478 152207 675530 152213
rect 675478 152149 675530 152155
rect 675490 151700 675518 152149
rect 675382 151467 675434 151473
rect 675382 151409 675434 151415
rect 675394 151034 675422 151409
rect 675478 150357 675530 150363
rect 675478 150299 675530 150305
rect 675490 149850 675518 150299
rect 675476 148546 675532 148555
rect 675476 148481 675532 148490
rect 675188 148398 675244 148407
rect 675188 148333 675244 148342
rect 675490 148000 675518 148481
rect 675764 146622 675820 146631
rect 675764 146557 675820 146566
rect 675778 146150 675806 146557
rect 674708 139074 674764 139083
rect 674708 139009 674764 139018
rect 674722 138597 674750 139009
rect 674710 138591 674762 138597
rect 674710 138533 674762 138539
rect 674420 138482 674476 138491
rect 674420 138417 674422 138426
rect 674474 138417 674476 138426
rect 674422 138385 674474 138391
rect 674612 137298 674668 137307
rect 674612 137233 674668 137242
rect 674626 135637 674654 137233
rect 674708 135670 674764 135679
rect 655414 135631 655466 135637
rect 655414 135573 655466 135579
rect 674614 135631 674666 135637
rect 674708 135605 674764 135614
rect 674614 135573 674666 135579
rect 674722 135415 674750 135605
rect 646486 135409 646538 135415
rect 646486 135351 646538 135357
rect 674710 135409 674762 135415
rect 674710 135351 674762 135357
rect 646498 120435 646526 135351
rect 673556 134930 673612 134939
rect 673486 134888 673556 134916
rect 673556 134865 673612 134874
rect 675476 131822 675532 131831
rect 675476 131757 675532 131766
rect 675188 131082 675244 131091
rect 675188 131017 675244 131026
rect 674804 128714 674860 128723
rect 674804 128649 674860 128658
rect 674516 124866 674572 124875
rect 674516 124801 674572 124810
rect 674324 124274 674380 124283
rect 674324 124209 674380 124218
rect 674132 123386 674188 123395
rect 674132 123321 674188 123330
rect 647732 121462 647788 121471
rect 647732 121397 647788 121406
rect 647746 121207 647774 121397
rect 647830 121275 647882 121281
rect 647830 121217 647882 121223
rect 647734 121201 647786 121207
rect 647842 121175 647870 121217
rect 647734 121143 647786 121149
rect 647828 121166 647884 121175
rect 647828 121101 647884 121110
rect 647926 121127 647978 121133
rect 647926 121069 647978 121075
rect 647938 120879 647966 121069
rect 647924 120870 647980 120879
rect 647924 120805 647980 120814
rect 646484 120426 646540 120435
rect 646484 120361 646540 120370
rect 674146 106185 674174 123321
rect 674338 107369 674366 124209
rect 674422 121201 674474 121207
rect 674422 121143 674474 121149
rect 674434 121101 674462 121143
rect 674420 121092 674476 121101
rect 674420 121027 674476 121036
rect 674530 110995 674558 124801
rect 674708 122350 674764 122359
rect 674708 122285 674764 122294
rect 674612 121314 674668 121323
rect 674722 121281 674750 122285
rect 674612 121249 674668 121258
rect 674710 121275 674762 121281
rect 674626 121133 674654 121249
rect 674710 121217 674762 121223
rect 674614 121127 674666 121133
rect 674614 121069 674666 121075
rect 674818 121004 674846 128649
rect 675092 127974 675148 127983
rect 675092 127909 675148 127918
rect 674900 127086 674956 127095
rect 674900 127021 674956 127030
rect 674626 120976 674846 121004
rect 674626 114843 674654 120976
rect 674806 118093 674858 118099
rect 674806 118035 674858 118041
rect 674710 118019 674762 118025
rect 674710 117961 674762 117967
rect 674614 114837 674666 114843
rect 674614 114779 674666 114785
rect 674518 110989 674570 110995
rect 674518 110931 674570 110937
rect 674326 107363 674378 107369
rect 674326 107305 674378 107311
rect 674134 106179 674186 106185
rect 674134 106121 674186 106127
rect 674722 105223 674750 117961
rect 674818 106999 674846 118035
rect 674914 111088 674942 127021
rect 675106 111458 675134 127909
rect 675202 112009 675230 131017
rect 675490 115805 675518 131757
rect 677012 130342 677068 130351
rect 677012 130277 677068 130286
rect 676916 126346 676972 126355
rect 676916 126281 676972 126290
rect 676820 125606 676876 125615
rect 676820 125541 676876 125550
rect 676834 118099 676862 125541
rect 676822 118093 676874 118099
rect 676822 118035 676874 118041
rect 676930 118025 676958 126281
rect 677026 120435 677054 130277
rect 677108 129602 677164 129611
rect 677108 129537 677164 129546
rect 677012 120426 677068 120435
rect 677012 120361 677068 120370
rect 677122 118067 677150 129537
rect 677108 118058 677164 118067
rect 676918 118019 676970 118025
rect 677108 117993 677164 118002
rect 676918 117961 676970 117967
rect 675478 115799 675530 115805
rect 675478 115741 675530 115747
rect 675478 115577 675530 115583
rect 675478 115519 675530 115525
rect 675490 115232 675518 115519
rect 675404 115204 675518 115232
rect 675404 115130 675432 115204
rect 675382 114837 675434 114843
rect 675382 114779 675434 114785
rect 675394 114478 675422 114779
rect 675380 114210 675436 114219
rect 675380 114145 675436 114154
rect 675394 113812 675422 114145
rect 675202 111981 675408 112009
rect 675106 111430 675408 111458
rect 674914 111060 675422 111088
rect 675094 110989 675146 110995
rect 675094 110931 675146 110937
rect 675106 110169 675134 110931
rect 675394 110778 675422 111060
rect 675106 110141 675408 110169
rect 675380 110066 675436 110075
rect 675380 110001 675436 110010
rect 675394 109594 675422 110001
rect 675092 109326 675148 109335
rect 675092 109261 675148 109270
rect 675106 108973 675134 109261
rect 675106 108945 675408 108973
rect 674806 106993 674858 106999
rect 674806 106935 674858 106941
rect 675106 106523 675134 108945
rect 675764 108142 675820 108151
rect 675764 108077 675820 108086
rect 675778 107670 675806 108077
rect 675382 107363 675434 107369
rect 675382 107305 675434 107311
rect 675394 107119 675422 107305
rect 675478 106993 675530 106999
rect 675478 106935 675530 106941
rect 675092 106514 675148 106523
rect 675490 106486 675518 106935
rect 675092 106449 675148 106458
rect 675382 106179 675434 106185
rect 675382 106121 675434 106127
rect 675394 105820 675422 106121
rect 674710 105217 674762 105223
rect 668180 105182 668236 105191
rect 674710 105159 674762 105165
rect 675382 105217 675434 105223
rect 675382 105159 675434 105165
rect 668180 105117 668236 105126
rect 665204 104590 665260 104599
rect 647926 104551 647978 104557
rect 665204 104525 665206 104534
rect 647926 104493 647978 104499
rect 665258 104525 665260 104534
rect 665206 104493 665258 104499
rect 647938 104303 647966 104493
rect 647924 104294 647980 104303
rect 647924 104229 647980 104238
rect 668194 99377 668222 105117
rect 675394 104636 675422 105159
rect 675380 103258 675436 103267
rect 675380 103193 675436 103202
rect 675394 102786 675422 103193
rect 675764 101482 675820 101491
rect 675764 101417 675820 101426
rect 675778 100936 675806 101417
rect 668182 99371 668234 99377
rect 668182 99313 668234 99319
rect 647350 92785 647402 92791
rect 647350 92727 647402 92733
rect 660694 92785 660746 92791
rect 660694 92727 660746 92733
rect 646678 92711 646730 92717
rect 646678 92653 646730 92659
rect 646198 92267 646250 92273
rect 646198 92209 646250 92215
rect 646210 85803 646238 92209
rect 646582 92193 646634 92199
rect 646582 92135 646634 92141
rect 646196 85794 646252 85803
rect 646196 85729 646252 85738
rect 645908 84166 645964 84175
rect 645908 84101 645964 84110
rect 645922 81839 645950 84101
rect 645910 81833 645962 81839
rect 645910 81775 645962 81781
rect 646486 76949 646538 76955
rect 646484 76914 646486 76923
rect 646538 76914 646540 76923
rect 646484 76849 646540 76858
rect 646486 76801 646538 76807
rect 646486 76743 646538 76749
rect 646498 76035 646526 76743
rect 646484 76026 646540 76035
rect 646484 75961 646540 75970
rect 646102 75839 646154 75845
rect 646102 75781 646154 75787
rect 646114 75295 646142 75781
rect 646486 75469 646538 75475
rect 646484 75434 646486 75443
rect 646538 75434 646540 75443
rect 646484 75369 646540 75378
rect 646100 75286 646156 75295
rect 646594 75272 646622 92135
rect 646100 75221 646156 75230
rect 646498 75244 646622 75272
rect 646100 72918 646156 72927
rect 646100 72853 646156 72862
rect 646114 72293 646142 72853
rect 646102 72287 646154 72293
rect 646102 72229 646154 72235
rect 646498 72187 646526 75244
rect 646690 72631 646718 92653
rect 647254 92489 647306 92495
rect 647254 92431 647306 92437
rect 646868 88162 646924 88171
rect 646868 88097 646924 88106
rect 646882 88055 646910 88097
rect 646870 88049 646922 88055
rect 646870 87991 646922 87997
rect 646870 85163 646922 85169
rect 646870 85105 646922 85111
rect 646882 85063 646910 85105
rect 646868 85054 646924 85063
rect 646868 84989 646924 84998
rect 647266 83879 647294 92431
rect 647252 83870 647308 83879
rect 647252 83805 647308 83814
rect 647362 80919 647390 92727
rect 659830 92711 659882 92717
rect 659830 92653 659882 92659
rect 647542 92637 647594 92643
rect 647542 92579 647594 92585
rect 647444 87422 647500 87431
rect 647444 87357 647500 87366
rect 647348 80910 647404 80919
rect 647348 80845 647404 80854
rect 647458 77769 647486 87357
rect 647554 82251 647582 92579
rect 659734 92489 659786 92495
rect 659734 92431 659786 92437
rect 647830 92415 647882 92421
rect 647830 92357 647882 92363
rect 647734 92341 647786 92347
rect 647734 92283 647786 92289
rect 647636 89050 647692 89059
rect 647636 88985 647692 88994
rect 647540 82242 647596 82251
rect 647540 82177 647596 82186
rect 647650 81691 647678 88985
rect 647746 85507 647774 92283
rect 647842 86247 647870 92357
rect 658870 92193 658922 92199
rect 658870 92135 658922 92141
rect 650902 88049 650954 88055
rect 650902 87991 650954 87997
rect 647924 87718 647980 87727
rect 647924 87653 647980 87662
rect 647938 87093 647966 87653
rect 647926 87087 647978 87093
rect 647926 87029 647978 87035
rect 647924 86534 647980 86543
rect 647924 86469 647926 86478
rect 647978 86469 647980 86478
rect 647926 86437 647978 86443
rect 647828 86238 647884 86247
rect 647828 86173 647884 86182
rect 647732 85498 647788 85507
rect 647732 85433 647788 85442
rect 650914 85359 650942 87991
rect 658882 87986 658910 92135
rect 659746 87852 659774 92431
rect 659842 88000 659870 92653
rect 659842 87972 660144 88000
rect 660706 87986 660734 92727
rect 661750 92637 661802 92643
rect 661750 92579 661802 92585
rect 661174 92267 661226 92273
rect 661174 92209 661226 92215
rect 661186 88000 661214 92209
rect 661762 88000 661790 92579
rect 663094 92415 663146 92421
rect 663094 92357 663146 92363
rect 662518 92341 662570 92347
rect 662518 92283 662570 92289
rect 661186 87972 661440 88000
rect 661762 87972 662016 88000
rect 662530 87986 662558 92283
rect 663106 87986 663134 92357
rect 659616 87824 659774 87852
rect 658006 87309 658058 87315
rect 656866 87232 657792 87260
rect 658058 87257 658320 87260
rect 658006 87251 658320 87257
rect 658018 87232 658320 87251
rect 650996 86978 651052 86987
rect 650996 86913 651052 86922
rect 650900 85350 650956 85359
rect 650900 85285 650956 85294
rect 651010 85169 651038 86913
rect 651094 86495 651146 86501
rect 651094 86437 651146 86443
rect 650998 85163 651050 85169
rect 650998 85105 651050 85111
rect 650996 84314 651052 84323
rect 650996 84249 651052 84258
rect 647926 83461 647978 83467
rect 647924 83426 647926 83435
rect 647978 83426 647980 83435
rect 647924 83361 647980 83370
rect 650900 82686 650956 82695
rect 650900 82621 650956 82630
rect 647924 82538 647980 82547
rect 647924 82473 647980 82482
rect 647938 81913 647966 82473
rect 647926 81907 647978 81913
rect 647926 81849 647978 81855
rect 647638 81685 647690 81691
rect 647638 81627 647690 81633
rect 647924 81354 647980 81363
rect 647924 81289 647926 81298
rect 647978 81289 647980 81298
rect 647926 81257 647978 81263
rect 647828 80466 647884 80475
rect 647828 80401 647884 80410
rect 647734 79317 647786 79323
rect 647734 79259 647786 79265
rect 647746 78995 647774 79259
rect 647732 78986 647788 78995
rect 647732 78921 647788 78930
rect 647842 78879 647870 80401
rect 647926 80205 647978 80211
rect 647924 80170 647926 80179
rect 647978 80170 647980 80179
rect 647924 80105 647980 80114
rect 647924 79282 647980 79291
rect 647924 79217 647980 79226
rect 647830 78873 647882 78879
rect 647830 78815 647882 78821
rect 647938 78361 647966 79217
rect 647926 78355 647978 78361
rect 647926 78297 647978 78303
rect 647446 77763 647498 77769
rect 647446 77705 647498 77711
rect 647926 77689 647978 77695
rect 647924 77654 647926 77663
rect 647978 77654 647980 77663
rect 647924 77589 647980 77598
rect 647926 77319 647978 77325
rect 647926 77261 647978 77267
rect 647938 77071 647966 77261
rect 647924 77062 647980 77071
rect 647924 76997 647980 77006
rect 650914 76807 650942 82621
rect 651010 77695 651038 84249
rect 651106 83435 651134 86437
rect 651188 86238 651244 86247
rect 651188 86173 651244 86182
rect 651092 83426 651148 83435
rect 651092 83361 651148 83370
rect 651202 79693 651230 86173
rect 651190 79687 651242 79693
rect 651190 79629 651242 79635
rect 650998 77689 651050 77695
rect 650998 77631 651050 77637
rect 650902 76801 650954 76807
rect 650902 76743 650954 76749
rect 656866 75475 656894 87232
rect 657046 87161 657098 87167
rect 657046 87103 657098 87109
rect 657058 83467 657086 87103
rect 663286 87087 663338 87093
rect 663286 87029 663338 87035
rect 663298 85211 663326 87029
rect 663380 85646 663436 85655
rect 663380 85581 663436 85590
rect 663284 85202 663340 85211
rect 663284 85137 663340 85146
rect 657046 83461 657098 83467
rect 657046 83403 657098 83409
rect 663394 82968 663422 85581
rect 663476 84758 663532 84767
rect 663476 84693 663532 84702
rect 663202 82940 663422 82968
rect 661078 81685 661130 81691
rect 661130 81633 661440 81636
rect 661078 81627 661440 81633
rect 661090 81608 661440 81627
rect 657538 81321 657792 81340
rect 657526 81315 657792 81321
rect 657578 81312 657792 81315
rect 657526 81257 657578 81263
rect 662900 81206 662956 81215
rect 662900 81141 662956 81150
rect 656962 81016 657216 81044
rect 656962 80211 656990 81016
rect 656950 80205 657002 80211
rect 656950 80147 657002 80153
rect 658306 76955 658334 81030
rect 658882 79323 658910 81030
rect 659602 80748 659630 81030
rect 659554 80729 659630 80748
rect 659446 80723 659498 80729
rect 659446 80665 659498 80671
rect 659542 80723 659630 80729
rect 659594 80720 659630 80723
rect 659542 80665 659594 80671
rect 658870 79317 658922 79323
rect 658870 79259 658922 79265
rect 659458 77769 659486 80665
rect 659446 77763 659498 77769
rect 659446 77705 659498 77711
rect 658294 76949 658346 76955
rect 658294 76891 658346 76897
rect 656854 75469 656906 75475
rect 656854 75411 656906 75417
rect 647252 74398 647308 74407
rect 647252 74333 647308 74342
rect 646868 73806 646924 73815
rect 646868 73741 646924 73750
rect 646676 72622 646732 72631
rect 646676 72557 646732 72566
rect 646882 72515 646910 73741
rect 647266 72589 647294 74333
rect 647254 72583 647306 72589
rect 647254 72525 647306 72531
rect 660130 72515 660158 81030
rect 660706 78879 660734 81030
rect 661762 81016 662016 81044
rect 660694 78873 660746 78879
rect 660694 78815 660746 78821
rect 661762 75845 661790 81016
rect 662530 78361 662558 81030
rect 662518 78355 662570 78361
rect 662518 78297 662570 78303
rect 662914 77325 662942 81141
rect 662902 77319 662954 77325
rect 662902 77261 662954 77267
rect 661750 75839 661802 75845
rect 661750 75781 661802 75787
rect 663202 72589 663230 82940
rect 663380 82834 663436 82843
rect 663380 82769 663436 82778
rect 663284 82094 663340 82103
rect 663284 82029 663340 82038
rect 663298 81913 663326 82029
rect 663286 81907 663338 81913
rect 663286 81849 663338 81855
rect 663394 81839 663422 82769
rect 663382 81833 663434 81839
rect 663382 81775 663434 81781
rect 663490 80156 663518 84693
rect 663394 80128 663518 80156
rect 663190 72583 663242 72589
rect 663190 72525 663242 72531
rect 646870 72509 646922 72515
rect 646870 72451 646922 72457
rect 660118 72509 660170 72515
rect 660118 72451 660170 72457
rect 663394 72293 663422 80128
rect 663382 72287 663434 72293
rect 663382 72229 663434 72235
rect 646484 72178 646540 72187
rect 646484 72113 646540 72122
rect 645718 51789 645770 51795
rect 645718 51731 645770 51737
rect 645622 46461 645674 46467
rect 645622 46403 645674 46409
rect 640724 40654 640780 40663
rect 640724 40589 640780 40598
rect 454964 40358 455020 40367
rect 454964 40293 455020 40302
rect 136532 40210 136588 40219
rect 136532 40145 136588 40154
<< via2 >>
rect 87860 995790 87916 995846
rect 92564 995790 92620 995846
rect 85940 995642 85996 995698
rect 92660 995642 92716 995698
rect 41780 968706 41836 968762
rect 41780 967078 41836 967134
rect 41780 965006 41836 965062
rect 41780 963970 41836 964026
rect 41780 963230 41836 963286
rect 42164 962786 42220 962842
rect 42068 962194 42124 962250
rect 42164 962046 42220 962102
rect 42452 962046 42508 962102
rect 42164 959530 42220 959586
rect 41780 959086 41836 959142
rect 41972 958346 42028 958402
rect 42164 957754 42220 957810
rect 41780 956570 41836 956626
rect 42452 949318 42508 949374
rect 42356 948447 42412 948486
rect 42356 948430 42358 948447
rect 42358 948430 42410 948447
rect 42410 948430 42412 948447
rect 42644 947877 42646 947894
rect 42646 947877 42698 947894
rect 42698 947877 42700 947894
rect 42644 947838 42700 947877
rect 40628 946506 40684 946562
rect 40244 945026 40300 945082
rect 37364 942806 37420 942862
rect 40436 944878 40492 944934
rect 40244 819966 40300 820022
rect 42836 939106 42892 939162
rect 42356 932446 42412 932502
rect 42356 930983 42412 931022
rect 42356 930966 42358 930983
rect 42358 930966 42410 930983
rect 42410 930966 42412 930983
rect 42164 823853 42166 823870
rect 42166 823853 42218 823870
rect 42218 823853 42220 823870
rect 42164 823814 42220 823853
rect 42164 823113 42166 823130
rect 42166 823113 42218 823130
rect 42218 823113 42220 823130
rect 42164 823074 42220 823113
rect 42164 822225 42166 822242
rect 42166 822225 42218 822242
rect 42218 822225 42220 822242
rect 42164 822186 42220 822225
rect 43220 821150 43276 821206
rect 40628 820706 40684 820762
rect 40436 819522 40492 819578
rect 37268 819078 37324 819134
rect 41684 817894 41740 817950
rect 40148 816710 40204 816766
rect 37364 812714 37420 812770
rect 40244 815822 40300 815878
rect 37364 802206 37420 802262
rect 37268 802058 37324 802114
rect 41492 811086 41548 811142
rect 40244 801910 40300 801966
rect 41588 809162 41644 809218
rect 42836 815674 42892 815730
rect 41876 813602 41932 813658
rect 41780 809606 41836 809662
rect 41684 800430 41740 800486
rect 41780 800282 41836 800338
rect 41972 812270 42028 812326
rect 42068 808274 42124 808330
rect 42068 800282 42124 800338
rect 43028 814934 43084 814990
rect 43028 810346 43084 810402
rect 42836 806942 42892 806998
rect 42836 805479 42892 805518
rect 42836 805462 42838 805479
rect 42838 805462 42890 805479
rect 42890 805462 42892 805479
rect 42452 802206 42508 802262
rect 42452 799690 42508 799746
rect 43124 807682 43180 807738
rect 43028 798358 43084 798414
rect 41876 794214 41932 794270
rect 42068 793770 42124 793826
rect 42452 792438 42508 792494
rect 42068 791106 42124 791162
rect 42164 790958 42220 791014
rect 43028 792290 43084 792346
rect 42836 791846 42892 791902
rect 42740 790514 42796 790570
rect 42164 788590 42220 788646
rect 42932 791698 42988 791754
rect 42740 780467 42796 780506
rect 42740 780450 42742 780467
rect 42742 780450 42794 780467
rect 42794 780450 42796 780467
rect 42740 779675 42742 779692
rect 42742 779675 42794 779692
rect 42794 779675 42796 779692
rect 42740 779636 42796 779675
rect 42740 778861 42742 778878
rect 42742 778861 42794 778878
rect 42794 778861 42796 778878
rect 42740 778822 42796 778861
rect 43316 777934 43372 777990
rect 43220 777194 43276 777250
rect 42932 774826 42988 774882
rect 38996 773494 39052 773550
rect 38804 772606 38860 772662
rect 37364 769498 37420 769554
rect 41492 771126 41548 771182
rect 41396 769054 41452 769110
rect 38804 760174 38860 760230
rect 37364 758694 37420 758750
rect 41876 770386 41932 770442
rect 41588 767870 41644 767926
rect 41780 765946 41836 766002
rect 41684 765206 41740 765262
rect 41588 757362 41644 757418
rect 41780 757066 41836 757122
rect 42068 767278 42124 767334
rect 41972 766390 42028 766446
rect 41972 758398 42028 758454
rect 43028 772458 43084 772514
rect 42164 763430 42220 763486
rect 42164 761967 42220 762006
rect 42164 761950 42166 761967
rect 42166 761950 42218 761967
rect 42218 761950 42220 761967
rect 43028 760470 43084 760526
rect 42068 757066 42124 757122
rect 42068 753070 42124 753126
rect 42068 751738 42124 751794
rect 42068 750998 42124 751054
rect 41780 748630 41836 748686
rect 41780 747446 41836 747502
rect 41876 747298 41932 747354
rect 43220 751738 43276 751794
rect 43028 747150 43084 747206
rect 42932 746706 42988 746762
rect 42452 745966 42508 746022
rect 42836 737251 42892 737290
rect 42836 737234 42838 737251
rect 42838 737234 42890 737251
rect 42890 737234 42892 737251
rect 42164 736681 42166 736698
rect 42166 736681 42218 736698
rect 42218 736681 42220 736698
rect 42164 736642 42220 736681
rect 42836 735645 42838 735662
rect 42838 735645 42890 735662
rect 42890 735645 42892 735662
rect 42836 735606 42892 735645
rect 43220 734866 43276 734922
rect 43124 731610 43180 731666
rect 40244 730278 40300 730334
rect 41684 728798 41740 728854
rect 41588 725838 41644 725894
rect 41492 723174 41548 723230
rect 41396 722730 41452 722786
rect 41492 714294 41548 714350
rect 41396 714146 41452 714202
rect 41780 727910 41836 727966
rect 41684 714146 41740 714202
rect 41876 727170 41932 727226
rect 41780 713850 41836 713906
rect 42164 724654 42220 724710
rect 41972 724062 42028 724118
rect 42068 721990 42124 722046
rect 42452 720362 42508 720418
rect 42452 718751 42508 718790
rect 42452 718734 42454 718751
rect 42454 718734 42506 718751
rect 42506 718734 42508 718751
rect 42164 713850 42220 713906
rect 43124 711334 43180 711390
rect 43028 711038 43084 711094
rect 42068 708522 42124 708578
rect 41876 707930 41932 707986
rect 42740 707930 42796 707986
rect 41780 706746 41836 706802
rect 42452 705414 42508 705470
rect 42068 704674 42124 704730
rect 41780 704082 41836 704138
rect 43124 709706 43180 709762
rect 43028 702750 43084 702806
rect 42836 694035 42892 694074
rect 42836 694018 42838 694035
rect 42838 694018 42890 694035
rect 42890 694018 42892 694035
rect 42452 693426 42508 693482
rect 42452 692725 42454 692742
rect 42454 692725 42506 692742
rect 42506 692725 42508 692742
rect 42452 692686 42508 692725
rect 43316 733978 43372 734034
rect 43412 711482 43468 711538
rect 43508 691650 43564 691706
rect 43220 690762 43276 690818
rect 41684 688246 41740 688302
rect 40148 687062 40204 687118
rect 37364 683214 37420 683270
rect 37364 672558 37420 672614
rect 40244 686322 40300 686378
rect 40916 684842 40972 684898
rect 40244 673890 40300 673946
rect 41300 681438 41356 681494
rect 41300 670930 41356 670986
rect 41780 685582 41836 685638
rect 41972 683954 42028 684010
rect 41876 679514 41932 679570
rect 42068 682622 42124 682678
rect 43028 681290 43084 681346
rect 42164 678774 42220 678830
rect 42452 676702 42508 676758
rect 42452 675666 42508 675722
rect 41972 670782 42028 670838
rect 42164 670930 42220 670986
rect 42164 670821 42166 670838
rect 42166 670821 42218 670838
rect 42218 670821 42220 670838
rect 42164 670782 42220 670821
rect 42068 670634 42124 670690
rect 42164 670338 42220 670394
rect 43124 678182 43180 678238
rect 43124 670930 43180 670986
rect 42164 665306 42220 665362
rect 42452 662790 42508 662846
rect 42164 661458 42220 661514
rect 42164 660718 42220 660774
rect 41780 660274 41836 660330
rect 41876 659090 41932 659146
rect 42836 663382 42892 663438
rect 43124 662346 43180 662402
rect 41780 656574 41836 656630
rect 42452 651098 42508 651154
rect 42452 649783 42508 649822
rect 42452 649766 42454 649783
rect 42454 649766 42506 649783
rect 42506 649766 42508 649783
rect 42452 649509 42454 649526
rect 42454 649509 42506 649526
rect 42506 649509 42508 649526
rect 42452 649470 42508 649509
rect 43220 648434 43276 648490
rect 43124 645326 43180 645382
rect 39860 643846 39916 643902
rect 37364 639998 37420 640054
rect 37364 628158 37420 628214
rect 39956 643106 40012 643162
rect 41492 642366 41548 642422
rect 41300 639406 41356 639462
rect 39956 627862 40012 627918
rect 41684 641626 41740 641682
rect 41588 636298 41644 636354
rect 41300 627714 41356 627770
rect 41588 627714 41644 627770
rect 41876 640738 41932 640794
rect 41972 637630 42028 637686
rect 42068 636742 42124 636798
rect 42164 635558 42220 635614
rect 43028 634966 43084 635022
rect 42452 633486 42508 633542
rect 42452 632302 42508 632358
rect 42164 627566 42220 627622
rect 42068 627418 42124 627474
rect 42068 621646 42124 621702
rect 41972 620758 42028 620814
rect 41780 618242 41836 618298
rect 41972 618094 42028 618150
rect 41780 617798 41836 617854
rect 41780 616466 41836 616522
rect 41780 613358 41836 613414
rect 41780 612766 41836 612822
rect 42740 607699 42742 607716
rect 42742 607699 42794 607716
rect 42794 607699 42796 607716
rect 42740 607660 42796 607699
rect 42740 606863 42796 606902
rect 42740 606846 42742 606863
rect 42742 606846 42794 606863
rect 42794 606846 42796 606863
rect 42164 606254 42220 606310
rect 43892 680550 43948 680606
rect 43508 647546 43564 647602
rect 43604 646954 43660 647010
rect 43316 625050 43372 625106
rect 43508 605218 43564 605274
rect 43220 604626 43276 604682
rect 43412 602850 43468 602906
rect 41588 601814 41644 601870
rect 40052 600630 40108 600686
rect 41396 598410 41452 598466
rect 41492 596190 41548 596246
rect 41876 599150 41932 599206
rect 41780 595154 41836 595210
rect 41588 584794 41644 584850
rect 41492 584646 41548 584702
rect 41396 584498 41452 584554
rect 41972 597522 42028 597578
rect 41876 584350 41932 584406
rect 42068 593082 42124 593138
rect 42164 592342 42220 592398
rect 42068 584202 42124 584258
rect 42836 591750 42892 591806
rect 42740 590418 42796 590474
rect 42740 589382 42796 589438
rect 42740 584646 42796 584702
rect 42836 583758 42892 583814
rect 41972 581982 42028 582038
rect 42932 581390 42988 581446
rect 41780 580206 41836 580262
rect 42164 578874 42220 578930
rect 42932 578282 42988 578338
rect 41780 576950 41836 577006
rect 42452 576358 42508 576414
rect 41780 575914 41836 575970
rect 41780 575026 41836 575082
rect 42164 574582 42220 574638
rect 42452 573102 42508 573158
rect 43028 577542 43084 577598
rect 34484 564666 34540 564722
rect 42164 563499 42220 563538
rect 42164 563482 42166 563499
rect 42166 563482 42218 563499
rect 42218 563482 42220 563499
rect 43124 573990 43180 574046
rect 42836 562816 42892 562872
rect 43220 562002 43276 562058
rect 42932 558894 42988 558950
rect 40244 557414 40300 557470
rect 41396 555934 41452 555990
rect 41684 555934 41740 555990
rect 41396 552974 41452 553030
rect 41588 551938 41644 551994
rect 41012 544094 41068 544150
rect 42164 555194 42220 555250
rect 41972 554306 42028 554362
rect 41780 552974 41836 553030
rect 41492 541282 41548 541338
rect 41684 541282 41740 541338
rect 41876 540986 41932 541042
rect 42068 550014 42124 550070
rect 42452 551346 42508 551402
rect 42452 551198 42508 551254
rect 42452 541134 42508 541190
rect 42932 549274 42988 549330
rect 43028 548534 43084 548590
rect 42164 540986 42220 541042
rect 41876 538914 41932 538970
rect 42068 536990 42124 537046
rect 42164 535214 42220 535270
rect 41972 533734 42028 533790
rect 42164 532698 42220 532754
rect 41780 531810 41836 531866
rect 42932 534474 42988 534530
rect 42452 531366 42508 531422
rect 42932 530034 42988 530090
rect 41780 526482 41836 526538
rect 41588 524114 41644 524170
rect 41588 503986 41644 504042
rect 41780 490962 41836 491018
rect 41780 481046 41836 481102
rect 42164 510054 42220 510110
rect 42164 503986 42220 504042
rect 42260 437129 42262 437146
rect 42262 437129 42314 437146
rect 42314 437129 42316 437146
rect 42260 437090 42316 437129
rect 42260 436241 42262 436258
rect 42262 436241 42314 436258
rect 42314 436241 42316 436258
rect 42260 436202 42316 436241
rect 41876 435462 41932 435518
rect 43796 646066 43852 646122
rect 43604 603738 43660 603794
rect 43508 561558 43564 561614
rect 43796 602850 43852 602906
rect 43604 560522 43660 560578
rect 43412 559782 43468 559838
rect 43316 547646 43372 547702
rect 43316 546166 43372 546222
rect 43316 434426 43372 434482
rect 43220 433538 43276 433594
rect 41972 429838 42028 429894
rect 41780 426878 41836 426934
rect 37364 423622 37420 423678
rect 37268 421994 37324 422050
rect 40148 423178 40204 423234
rect 40244 421254 40300 421310
rect 43604 432946 43660 433002
rect 43412 432058 43468 432114
rect 42548 424362 42604 424418
rect 42356 419922 42412 419978
rect 42356 418459 42412 418498
rect 42356 418442 42358 418459
rect 42358 418442 42410 418459
rect 42410 418442 42412 418459
rect 43124 420958 43180 421014
rect 42068 406306 42124 406362
rect 42164 405122 42220 405178
rect 41780 403642 41836 403698
rect 42260 403198 42316 403254
rect 43508 403198 43564 403254
rect 43700 403198 43756 403254
rect 41780 402606 41836 402662
rect 41780 401866 41836 401922
rect 41780 400090 41836 400146
rect 41780 399498 41836 399554
rect 41780 398758 41836 398814
rect 42356 393913 42358 393930
rect 42358 393913 42410 393930
rect 42410 393913 42412 393930
rect 42356 393874 42412 393913
rect 42644 392877 42646 392894
rect 42646 392877 42698 392894
rect 42698 392877 42700 392894
rect 42644 392838 42700 392877
rect 42356 392285 42358 392302
rect 42358 392285 42410 392302
rect 42410 392285 42412 392302
rect 42356 392246 42412 392285
rect 43220 391210 43276 391266
rect 41972 386622 42028 386678
rect 37268 381146 37324 381202
rect 40148 380406 40204 380462
rect 40052 379962 40108 380018
rect 37364 378778 37420 378834
rect 40244 378038 40300 378094
rect 38324 370490 38380 370546
rect 42356 383514 42412 383570
rect 42260 376558 42316 376614
rect 42260 375243 42316 375282
rect 42260 375226 42262 375243
rect 42262 375226 42314 375243
rect 42314 375226 42316 375243
rect 43124 377742 43180 377798
rect 42068 362794 42124 362850
rect 41876 361906 41932 361962
rect 41780 360574 41836 360630
rect 42260 360130 42316 360186
rect 41780 359390 41836 359446
rect 41780 358650 41836 358706
rect 41780 356874 41836 356930
rect 41780 356430 41836 356486
rect 41780 355542 41836 355598
rect 42356 350697 42358 350714
rect 42358 350697 42410 350714
rect 42410 350697 42412 350714
rect 42356 350658 42412 350697
rect 42356 349957 42358 349974
rect 42358 349957 42410 349974
rect 42410 349957 42412 349974
rect 42356 349918 42412 349957
rect 42356 349069 42358 349086
rect 42358 349069 42410 349086
rect 42410 349069 42412 349086
rect 42356 349030 42412 349069
rect 43508 390914 43564 390970
rect 43220 347698 43276 347754
rect 43220 347550 43276 347606
rect 41876 343554 41932 343610
rect 41780 340298 41836 340354
rect 37364 339854 37420 339910
rect 37172 337338 37228 337394
rect 39956 337930 40012 337986
rect 37364 336450 37420 336506
rect 37364 335562 37420 335618
rect 40052 337190 40108 337246
rect 40244 334822 40300 334878
rect 42548 334378 42604 334434
rect 42260 333490 42316 333546
rect 42260 332027 42316 332066
rect 42260 332010 42262 332027
rect 42262 332010 42314 332027
rect 42314 332010 42316 332027
rect 42068 319726 42124 319782
rect 41876 318690 41932 318746
rect 41780 317802 41836 317858
rect 41780 316026 41836 316082
rect 41780 315434 41836 315490
rect 41876 313658 41932 313714
rect 41780 313214 41836 313270
rect 41780 312326 41836 312382
rect 42356 307481 42358 307498
rect 42358 307481 42410 307498
rect 42410 307481 42412 307498
rect 42356 307442 42412 307481
rect 42356 306741 42358 306758
rect 42358 306741 42410 306758
rect 42410 306741 42412 306758
rect 42356 306702 42412 306741
rect 42356 305370 42412 305426
rect 43220 304038 43276 304094
rect 43220 303890 43276 303946
rect 41876 300338 41932 300394
rect 37364 296638 37420 296694
rect 37268 293974 37324 294030
rect 40052 294714 40108 294770
rect 37364 292346 37420 292402
rect 40148 293974 40204 294030
rect 40244 291606 40300 291662
rect 40532 284058 40588 284114
rect 42260 297230 42316 297286
rect 42452 292346 42508 292402
rect 42260 288794 42316 288850
rect 42260 283318 42316 283374
rect 42932 291310 42988 291366
rect 42452 282430 42508 282486
rect 41780 279766 41836 279822
rect 41780 276510 41836 276566
rect 41972 275474 42028 275530
rect 41780 274882 41836 274938
rect 42164 274142 42220 274198
rect 42260 273698 42316 273754
rect 41780 272958 41836 273014
rect 41780 272218 41836 272274
rect 41780 270590 41836 270646
rect 42548 270442 42604 270498
rect 41780 269998 41836 270054
rect 41780 269110 41836 269166
rect 42260 264265 42262 264282
rect 42262 264265 42314 264282
rect 42314 264265 42316 264282
rect 42260 264226 42316 264265
rect 42644 263229 42646 263246
rect 42646 263229 42698 263246
rect 42698 263229 42700 263246
rect 42644 263190 42700 263229
rect 42644 262450 42700 262506
rect 41300 259490 41356 259546
rect 40244 251498 40300 251554
rect 37364 250758 37420 250814
rect 40052 250758 40108 250814
rect 40148 248390 40204 248446
rect 42068 257122 42124 257178
rect 41780 254310 41836 254366
rect 40244 242026 40300 242082
rect 43508 261562 43564 261618
rect 43220 260822 43276 260878
rect 43412 259342 43468 259398
rect 42548 249130 42604 249186
rect 42164 247058 42220 247114
rect 42356 246762 42412 246818
rect 43028 247502 43084 247558
rect 42356 245578 42412 245634
rect 42356 239362 42412 239418
rect 42452 238918 42508 238974
rect 41780 233294 41836 233350
rect 41972 231666 42028 231722
rect 41972 230926 42028 230982
rect 41780 230334 41836 230390
rect 41780 229742 41836 229798
rect 41780 229002 41836 229058
rect 41780 227226 41836 227282
rect 41780 226634 41836 226690
rect 42068 226190 42124 226246
rect 42356 221049 42358 221066
rect 42358 221049 42410 221066
rect 42410 221049 42412 221066
rect 42356 221010 42412 221049
rect 42356 220309 42358 220326
rect 42358 220309 42410 220326
rect 42410 220309 42412 220326
rect 42356 220270 42412 220309
rect 42356 219421 42358 219438
rect 42358 219421 42410 219438
rect 42410 219421 42412 219438
rect 42356 219382 42412 219421
rect 43220 217606 43276 217662
rect 43316 216866 43372 216922
rect 47444 946210 47500 946266
rect 43412 216126 43468 216182
rect 41972 213906 42028 213962
rect 40244 210798 40300 210854
rect 40052 207098 40108 207154
rect 37364 206062 37420 206118
rect 40148 205174 40204 205230
rect 40916 198701 40918 198718
rect 40918 198701 40970 198718
rect 40970 198701 40972 198718
rect 40916 198662 40972 198701
rect 42068 209170 42124 209226
rect 42836 208874 42892 208930
rect 42356 207838 42412 207894
rect 42356 204325 42358 204342
rect 42358 204325 42410 204342
rect 42410 204325 42412 204342
rect 42356 204286 42412 204325
rect 42356 202806 42412 202862
rect 42164 197478 42220 197534
rect 43124 204878 43180 204934
rect 42356 195110 42412 195166
rect 41780 190966 41836 191022
rect 41780 190078 41836 190134
rect 41972 189042 42028 189098
rect 41780 188302 41836 188358
rect 41780 185934 41836 185990
rect 47732 946062 47788 946118
rect 59444 975366 59500 975422
rect 47924 944730 47980 944786
rect 62036 992090 62092 992146
rect 80756 995198 80812 995254
rect 80180 993718 80236 993774
rect 86516 995494 86572 995550
rect 85364 995346 85420 995402
rect 84500 993866 84556 993922
rect 83444 993570 83500 993626
rect 92852 993570 92908 993626
rect 62036 962194 62092 962250
rect 61844 962046 61900 962102
rect 59540 960862 59596 960918
rect 57812 946654 57868 946710
rect 59540 932298 59596 932354
rect 59540 917794 59596 917850
rect 59540 903438 59596 903494
rect 59540 889082 59596 889138
rect 59540 874726 59596 874782
rect 58580 860370 58636 860426
rect 59540 846014 59596 846070
rect 59540 831658 59596 831714
rect 59540 817302 59596 817358
rect 59540 802798 59596 802854
rect 59540 788590 59596 788646
rect 59540 774086 59596 774142
rect 59540 759730 59596 759786
rect 59540 745522 59596 745578
rect 59540 731018 59596 731074
rect 59540 716662 59596 716718
rect 59540 702306 59596 702362
rect 59540 687950 59596 688006
rect 59540 673594 59596 673650
rect 59540 659238 59596 659294
rect 59252 644882 59308 644938
rect 53780 589382 53836 589438
rect 59540 630526 59596 630582
rect 59540 616170 59596 616226
rect 59540 601853 59542 601870
rect 59542 601853 59594 601870
rect 59594 601853 59596 601870
rect 59540 601814 59596 601853
rect 58196 587475 58252 587514
rect 58196 587458 58198 587475
rect 58198 587458 58250 587475
rect 58250 587458 58252 587475
rect 59540 572954 59596 573010
rect 59444 558894 59500 558950
rect 59540 544390 59596 544446
rect 59540 530034 59596 530090
rect 59540 515678 59596 515734
rect 59540 501191 59596 501230
rect 59540 501174 59542 501191
rect 59542 501174 59594 501191
rect 59594 501174 59596 501191
rect 58580 486818 58636 486874
rect 59540 472462 59596 472518
rect 59540 458106 59596 458162
rect 59540 443750 59596 443806
rect 59540 429394 59596 429450
rect 58388 415038 58444 415094
rect 57620 400682 57676 400738
rect 59252 386326 59308 386382
rect 59540 371822 59596 371878
rect 60212 357614 60268 357670
rect 58388 343110 58444 343166
rect 57812 328754 57868 328810
rect 58004 314546 58060 314602
rect 59444 300042 59500 300098
rect 58100 285834 58156 285890
rect 65108 246466 65164 246522
rect 115700 1005597 115702 1005614
rect 115702 1005597 115754 1005614
rect 115754 1005597 115756 1005614
rect 115700 1005558 115756 1005597
rect 102164 1005427 102220 1005466
rect 312788 1005449 312790 1005466
rect 312790 1005449 312842 1005466
rect 312842 1005449 312844 1005466
rect 102164 1005410 102166 1005427
rect 102166 1005410 102218 1005427
rect 102218 1005410 102220 1005427
rect 101492 1005301 101494 1005318
rect 101494 1005301 101546 1005318
rect 101546 1005301 101548 1005318
rect 101492 1005262 101548 1005301
rect 114164 1005279 114220 1005318
rect 114164 1005262 114166 1005279
rect 114166 1005262 114218 1005279
rect 114218 1005262 114220 1005279
rect 105428 1005153 105430 1005170
rect 105430 1005153 105482 1005170
rect 105482 1005153 105484 1005170
rect 105428 1005114 105484 1005153
rect 108884 1003673 108886 1003690
rect 108886 1003673 108938 1003690
rect 108938 1003673 108940 1003690
rect 108884 1003634 108940 1003673
rect 102836 1002467 102892 1002506
rect 102836 1002450 102838 1002467
rect 102838 1002450 102890 1002467
rect 102890 1002450 102892 1002467
rect 94964 995642 95020 995698
rect 100532 1002319 100588 1002358
rect 103796 1002341 103798 1002358
rect 103798 1002341 103850 1002358
rect 103850 1002341 103852 1002358
rect 100532 1002302 100534 1002319
rect 100534 1002302 100586 1002319
rect 100586 1002302 100588 1002319
rect 103796 1002302 103852 1002341
rect 104468 1002319 104524 1002358
rect 104468 1002302 104470 1002319
rect 104470 1002302 104522 1002319
rect 104522 1002302 104524 1002319
rect 99764 995198 99820 995254
rect 106964 995938 107020 995994
rect 113300 995938 113356 995994
rect 113396 995807 113452 995846
rect 113396 995790 113398 995807
rect 113398 995790 113450 995807
rect 113450 995790 113452 995807
rect 115220 995494 115276 995550
rect 108212 995346 108268 995402
rect 106484 993718 106540 993774
rect 109844 995198 109900 995254
rect 115316 995346 115372 995402
rect 209012 1005153 209014 1005170
rect 209014 1005153 209066 1005170
rect 209066 1005153 209068 1005170
rect 151220 1002467 151276 1002506
rect 151220 1002450 151222 1002467
rect 151222 1002450 151274 1002467
rect 151274 1002450 151276 1002467
rect 157940 1002489 157942 1002506
rect 157942 1002489 157994 1002506
rect 157994 1002489 157996 1002506
rect 157940 1002450 157996 1002489
rect 136724 995790 136780 995846
rect 137972 995790 138028 995846
rect 137588 995642 137644 995698
rect 139220 995642 139276 995698
rect 129716 993866 129772 993922
rect 137396 995494 137452 995550
rect 150356 1002341 150358 1002358
rect 150358 1002341 150410 1002358
rect 150410 1002341 150412 1002358
rect 150356 1002302 150412 1002341
rect 144020 995938 144076 995994
rect 143924 995790 143980 995846
rect 140372 995346 140428 995402
rect 141140 995346 141196 995402
rect 160244 1000839 160300 1000878
rect 160244 1000822 160246 1000839
rect 160246 1000822 160298 1000839
rect 160298 1000822 160300 1000839
rect 156884 999381 156886 999398
rect 156886 999381 156938 999398
rect 156938 999381 156940 999398
rect 156884 999342 156940 999381
rect 162260 996103 162316 996142
rect 162260 996086 162262 996103
rect 162262 996086 162314 996103
rect 162314 996086 162316 996103
rect 163124 996125 163126 996142
rect 163126 996125 163178 996142
rect 163178 996125 163180 996142
rect 163124 996086 163180 996125
rect 164084 996086 164140 996142
rect 145268 995938 145324 995994
rect 149108 995938 149164 995994
rect 149492 995938 149548 995994
rect 151988 995955 152044 995994
rect 151988 995938 151990 995955
rect 151990 995938 152042 995955
rect 152042 995938 152044 995955
rect 152852 995938 152908 995994
rect 155348 995938 155404 995994
rect 164180 995977 164182 995994
rect 164182 995977 164234 995994
rect 164234 995977 164236 995994
rect 164180 995938 164236 995977
rect 154292 995807 154348 995846
rect 154292 995790 154294 995807
rect 154294 995790 154346 995807
rect 154346 995790 154348 995807
rect 156308 995790 156364 995846
rect 165620 995807 165676 995846
rect 165620 995790 165622 995807
rect 165622 995790 165674 995807
rect 165674 995790 165676 995807
rect 166196 995790 166252 995846
rect 159572 995642 159628 995698
rect 152852 995494 152908 995550
rect 158804 995494 158860 995550
rect 158996 995494 159052 995550
rect 158996 993866 159052 993922
rect 161204 995215 161260 995254
rect 161204 995198 161206 995215
rect 161206 995198 161258 995215
rect 161258 995198 161260 995215
rect 185108 995790 185164 995846
rect 188756 995790 188812 995846
rect 195188 995790 195244 995846
rect 170324 995642 170380 995698
rect 178484 995642 178540 995698
rect 185204 995642 185260 995698
rect 166964 995198 167020 995254
rect 167156 995050 167212 995106
rect 181460 995050 181516 995106
rect 184340 995494 184396 995550
rect 183764 995198 183820 995254
rect 182996 994162 183052 994218
rect 195092 995642 195148 995698
rect 185396 994014 185452 994070
rect 189428 995494 189484 995550
rect 191540 993866 191596 993922
rect 209012 1005114 209068 1005153
rect 208340 1001009 208342 1001026
rect 208342 1001009 208394 1001026
rect 208394 1001009 208396 1001026
rect 208340 1000970 208396 1001009
rect 211700 1000839 211756 1000878
rect 211700 1000822 211702 1000839
rect 211702 1000822 211754 1000839
rect 211754 1000822 211756 1000839
rect 256436 999507 256492 999546
rect 256436 999490 256438 999507
rect 256438 999490 256490 999507
rect 256490 999490 256492 999507
rect 204212 996547 204268 996586
rect 204212 996530 204214 996547
rect 204214 996530 204266 996547
rect 204266 996530 204268 996547
rect 213332 996103 213388 996142
rect 213332 996086 213334 996103
rect 213334 996086 213386 996103
rect 213386 996086 213388 996103
rect 214100 996125 214102 996142
rect 214102 996125 214154 996142
rect 214154 996125 214156 996142
rect 214100 996086 214156 996125
rect 215636 996103 215692 996142
rect 215636 996086 215638 996103
rect 215638 996086 215690 996103
rect 215690 996086 215692 996103
rect 198644 995955 198700 995994
rect 198644 995938 198646 995955
rect 198646 995938 198698 995955
rect 198698 995938 198700 995955
rect 203444 995955 203500 995994
rect 203444 995938 203446 995955
rect 203446 995938 203498 995955
rect 203498 995938 203500 995955
rect 205652 995938 205708 995994
rect 206516 995938 206572 995994
rect 201716 995790 201772 995846
rect 202868 995790 202924 995846
rect 204980 995807 205036 995846
rect 204980 995790 204982 995807
rect 204982 995790 205034 995807
rect 205034 995790 205036 995807
rect 201524 995050 201580 995106
rect 201716 995494 201772 995550
rect 205652 995346 205708 995402
rect 206996 995659 207052 995698
rect 206996 995642 206998 995659
rect 206998 995642 207050 995659
rect 207050 995642 207052 995659
rect 210260 995346 210316 995402
rect 211028 995346 211084 995402
rect 212660 995346 212716 995402
rect 201716 995237 201718 995254
rect 201718 995237 201770 995254
rect 201770 995237 201772 995254
rect 201716 995198 201772 995237
rect 210260 994162 210316 994218
rect 215444 995977 215446 995994
rect 215446 995977 215498 995994
rect 215498 995977 215500 995994
rect 215444 995938 215500 995977
rect 217076 995955 217132 995994
rect 217076 995938 217078 995955
rect 217078 995938 217130 995955
rect 217130 995938 217132 995955
rect 221780 995938 221836 995994
rect 241844 995790 241900 995846
rect 243860 995790 243916 995846
rect 259508 999381 259510 999398
rect 259510 999381 259562 999398
rect 259562 999381 259564 999398
rect 259508 999342 259564 999381
rect 263060 996547 263116 996586
rect 263060 996530 263062 996547
rect 263062 996530 263114 996547
rect 263114 996530 263116 996547
rect 246932 995938 246988 995994
rect 247508 995938 247564 995994
rect 222932 995642 222988 995698
rect 240788 995642 240844 995698
rect 227348 995050 227404 995106
rect 227540 995050 227596 995106
rect 232148 994310 232204 994366
rect 234356 994162 234412 994218
rect 235796 994458 235852 994514
rect 236756 994014 236812 994070
rect 239540 995494 239596 995550
rect 240212 995346 240268 995402
rect 242324 994606 242380 994662
rect 242324 994310 242380 994366
rect 242516 994310 242572 994366
rect 247412 995050 247468 995106
rect 244820 994310 244876 994366
rect 242516 994014 242572 994070
rect 243188 994014 243244 994070
rect 250100 995346 250156 995402
rect 265940 996125 265942 996142
rect 265942 996125 265994 996142
rect 265994 996125 265996 996142
rect 265940 996086 265996 996125
rect 266996 996103 267052 996142
rect 266996 996086 266998 996103
rect 266998 996086 267050 996103
rect 267050 996086 267052 996103
rect 258836 995955 258892 995994
rect 258836 995938 258838 995955
rect 258838 995938 258890 995955
rect 258890 995938 258892 995955
rect 264692 995977 264694 995994
rect 264694 995977 264746 995994
rect 264746 995977 264748 995994
rect 264692 995938 264748 995977
rect 251252 995790 251308 995846
rect 254804 995807 254860 995846
rect 254804 995790 254806 995807
rect 254806 995790 254858 995807
rect 254858 995790 254860 995807
rect 255572 995829 255574 995846
rect 255574 995829 255626 995846
rect 255626 995829 255628 995846
rect 255572 995790 255628 995829
rect 257492 995790 257548 995846
rect 258260 995790 258316 995846
rect 260756 995790 260812 995846
rect 268244 995807 268300 995846
rect 268244 995790 268246 995807
rect 268246 995790 268298 995807
rect 268298 995790 268300 995807
rect 250484 994606 250540 994662
rect 247604 994458 247660 994514
rect 254708 995346 254764 995402
rect 259124 995050 259180 995106
rect 254708 994162 254764 994218
rect 268436 995790 268492 995846
rect 262388 995642 262444 995698
rect 262196 995050 262252 995106
rect 262196 994754 262252 994810
rect 264020 995346 264076 995402
rect 273620 995790 273676 995846
rect 270740 995642 270796 995698
rect 283124 995790 283180 995846
rect 294836 995790 294892 995846
rect 286292 995642 286348 995698
rect 292532 995494 292588 995550
rect 298388 995938 298444 995994
rect 298292 995790 298348 995846
rect 312788 1005410 312844 1005449
rect 313844 1005427 313900 1005466
rect 313844 1005410 313846 1005427
rect 313846 1005410 313898 1005427
rect 313898 1005410 313900 1005427
rect 321044 1005410 321100 1005466
rect 321428 1005410 321484 1005466
rect 325460 1005410 325516 1005466
rect 365108 1005449 365110 1005466
rect 365110 1005449 365162 1005466
rect 365162 1005449 365164 1005466
rect 365108 1005410 365164 1005449
rect 298484 995642 298540 995698
rect 308756 1005279 308812 1005318
rect 308756 1005262 308758 1005279
rect 308758 1005262 308810 1005279
rect 308810 1005262 308812 1005279
rect 309620 1005301 309622 1005318
rect 309622 1005301 309674 1005318
rect 309674 1005301 309676 1005318
rect 309620 1005262 309676 1005301
rect 318644 1005279 318700 1005318
rect 318644 1005262 318646 1005279
rect 318646 1005262 318698 1005279
rect 318698 1005262 318700 1005279
rect 358676 1005301 358678 1005318
rect 358678 1005301 358730 1005318
rect 358730 1005301 358732 1005318
rect 358676 1005262 358732 1005301
rect 359924 1005279 359980 1005318
rect 359924 1005262 359926 1005279
rect 359926 1005262 359978 1005279
rect 359978 1005262 359980 1005279
rect 310292 1005153 310294 1005170
rect 310294 1005153 310346 1005170
rect 310346 1005153 310348 1005170
rect 310292 1005114 310348 1005153
rect 308084 1002598 308140 1002654
rect 314708 999507 314764 999546
rect 314708 999490 314710 999507
rect 314710 999490 314762 999507
rect 314762 999490 314764 999507
rect 315476 999529 315478 999546
rect 315478 999529 315530 999546
rect 315530 999529 315532 999546
rect 315476 999490 315532 999529
rect 311444 999381 311446 999398
rect 311446 999381 311498 999398
rect 311498 999381 311500 999398
rect 311444 999342 311500 999381
rect 299156 995642 299212 995698
rect 296660 994162 296716 994218
rect 317108 996103 317164 996142
rect 317108 996086 317110 996103
rect 317110 996086 317162 996103
rect 317162 996086 317164 996103
rect 318644 996125 318646 996142
rect 318646 996125 318698 996142
rect 318698 996125 318700 996142
rect 318644 996086 318700 996125
rect 305588 995938 305644 995994
rect 316340 995977 316342 995994
rect 316342 995977 316394 995994
rect 316394 995977 316396 995994
rect 316340 995938 316396 995977
rect 357044 1005153 357046 1005170
rect 357046 1005153 357098 1005170
rect 357098 1005153 357100 1005170
rect 328244 995938 328300 995994
rect 306452 995790 306508 995846
rect 307412 995790 307468 995846
rect 311924 995790 311980 995846
rect 325268 995642 325324 995698
rect 316724 995198 316780 995254
rect 316724 995050 316780 995106
rect 357044 1005114 357100 1005153
rect 364244 1005131 364300 1005170
rect 364244 1005114 364246 1005131
rect 364246 1005114 364298 1005131
rect 364298 1005114 364300 1005131
rect 357620 1003821 357622 1003838
rect 357622 1003821 357674 1003838
rect 357674 1003821 357676 1003838
rect 357620 1003782 357676 1003821
rect 359060 1003799 359116 1003838
rect 359060 1003782 359062 1003799
rect 359062 1003782 359114 1003799
rect 359114 1003782 359116 1003799
rect 355988 1003673 355990 1003690
rect 355990 1003673 356042 1003690
rect 356042 1003673 356044 1003690
rect 355988 1003634 356044 1003673
rect 360692 1000839 360748 1000878
rect 360692 1000822 360694 1000839
rect 360694 1000822 360746 1000839
rect 360746 1000822 360748 1000839
rect 361556 1000861 361558 1000878
rect 361558 1000861 361610 1000878
rect 361610 1000861 361612 1000878
rect 361556 1000822 361612 1000861
rect 367892 997901 367894 997918
rect 367894 997901 367946 997918
rect 367946 997901 367948 997918
rect 367892 997862 367948 997901
rect 369044 997731 369100 997770
rect 369044 997714 369046 997731
rect 369046 997714 369098 997731
rect 369098 997714 369100 997731
rect 362324 995938 362380 995994
rect 367124 995977 367126 995994
rect 367126 995977 367178 995994
rect 367178 995977 367180 995994
rect 367124 995938 367180 995977
rect 348692 995790 348748 995846
rect 339764 995198 339820 995254
rect 339764 994902 339820 994958
rect 365876 995790 365932 995846
rect 366644 995807 366700 995846
rect 366644 995790 366646 995807
rect 366646 995790 366698 995807
rect 366698 995790 366700 995807
rect 377300 995938 377356 995994
rect 379316 995938 379372 995994
rect 371828 995807 371884 995846
rect 371828 995790 371830 995807
rect 371830 995790 371882 995807
rect 371882 995790 371884 995807
rect 368660 995642 368716 995698
rect 374420 995642 374476 995698
rect 362804 995198 362860 995254
rect 368468 995198 368524 995254
rect 362804 995050 362860 995106
rect 368468 994754 368524 994810
rect 374516 995494 374572 995550
rect 380276 995494 380332 995550
rect 430868 1005427 430924 1005466
rect 430868 1005410 430870 1005427
rect 430870 1005410 430922 1005427
rect 430922 1005410 430924 1005427
rect 433172 1005449 433174 1005466
rect 433174 1005449 433226 1005466
rect 433226 1005449 433228 1005466
rect 433172 1005410 433228 1005449
rect 425300 1005279 425356 1005318
rect 425300 1005262 425302 1005279
rect 425302 1005262 425354 1005279
rect 425354 1005262 425356 1005279
rect 431540 1005301 431542 1005318
rect 431542 1005301 431594 1005318
rect 431594 1005301 431596 1005318
rect 431540 1005262 431596 1005301
rect 427604 1005153 427606 1005170
rect 427606 1005153 427658 1005170
rect 427658 1005153 427660 1005170
rect 427604 1005114 427660 1005153
rect 435572 1005131 435628 1005170
rect 435572 1005114 435574 1005131
rect 435574 1005114 435626 1005131
rect 435626 1005114 435628 1005131
rect 428084 1003947 428140 1003986
rect 428084 1003930 428086 1003947
rect 428086 1003930 428138 1003947
rect 428138 1003930 428140 1003947
rect 423380 1003799 423436 1003838
rect 423380 1003782 423382 1003799
rect 423382 1003782 423434 1003799
rect 423434 1003782 423436 1003799
rect 426452 1003821 426454 1003838
rect 426454 1003821 426506 1003838
rect 426506 1003821 426508 1003838
rect 426452 1003782 426508 1003821
rect 425780 1003673 425782 1003690
rect 425782 1003673 425834 1003690
rect 425834 1003673 425836 1003690
rect 425780 1003634 425836 1003673
rect 434036 1001135 434092 1001174
rect 434036 1001118 434038 1001135
rect 434038 1001118 434090 1001135
rect 434090 1001118 434092 1001135
rect 381716 995642 381772 995698
rect 377396 995346 377452 995402
rect 432500 1000987 432556 1001026
rect 432500 1000970 432502 1000987
rect 432502 1000970 432554 1000987
rect 432554 1000970 432556 1000987
rect 424148 1000839 424204 1000878
rect 424148 1000822 424150 1000839
rect 424150 1000822 424202 1000839
rect 424202 1000822 424204 1000839
rect 428948 1000861 428950 1000878
rect 428950 1000861 429002 1000878
rect 429002 1000861 429004 1000878
rect 428948 1000822 429004 1000861
rect 399860 996086 399916 996142
rect 385844 995790 385900 995846
rect 389108 995790 389164 995846
rect 393716 995790 393772 995846
rect 389396 995642 389452 995698
rect 386324 995494 386380 995550
rect 386324 995198 386380 995254
rect 383252 995050 383308 995106
rect 391796 995494 391852 995550
rect 396692 995346 396748 995402
rect 393044 995050 393100 995106
rect 390836 994162 390892 994218
rect 422516 995790 422572 995846
rect 399860 994754 399916 994810
rect 436340 996234 436396 996290
rect 436436 996125 436438 996142
rect 436438 996125 436490 996142
rect 436490 996125 436492 996142
rect 436436 996086 436492 996125
rect 554516 1005427 554572 1005466
rect 554516 1005410 554518 1005427
rect 554518 1005410 554570 1005427
rect 554570 1005410 554572 1005427
rect 429716 995938 429772 995994
rect 434132 995977 434134 995994
rect 434134 995977 434186 995994
rect 434186 995977 434188 995994
rect 434132 995938 434188 995977
rect 446228 995938 446284 995994
rect 438740 995807 438796 995846
rect 438740 995790 438742 995807
rect 438742 995790 438794 995807
rect 438794 995790 438796 995807
rect 440756 995642 440812 995698
rect 443540 995237 443542 995254
rect 443542 995237 443594 995254
rect 443594 995237 443596 995254
rect 443540 995198 443596 995237
rect 500660 1005279 500716 1005318
rect 556916 1005301 556918 1005318
rect 556918 1005301 556970 1005318
rect 556970 1005301 556972 1005318
rect 500660 1005262 500662 1005279
rect 500662 1005262 500714 1005279
rect 500714 1005262 500716 1005279
rect 556916 1005262 556972 1005301
rect 498164 1005114 498220 1005170
rect 501140 1005153 501142 1005170
rect 501142 1005153 501194 1005170
rect 501194 1005153 501196 1005170
rect 501140 1005114 501196 1005153
rect 467060 995642 467116 995698
rect 463604 995346 463660 995402
rect 471860 995938 471916 995994
rect 472244 995790 472300 995846
rect 488852 999342 488908 999398
rect 477044 995790 477100 995846
rect 485780 995790 485836 995846
rect 480980 995642 481036 995698
rect 472148 995494 472204 995550
rect 497588 999359 497644 999398
rect 497588 999342 497590 999359
rect 497590 999342 497642 999359
rect 497642 999342 497644 999359
rect 478388 995494 478444 995550
rect 471764 995346 471820 995402
rect 479924 995494 479980 995550
rect 482036 995346 482092 995402
rect 479828 994162 479884 994218
rect 488852 995494 488908 995550
rect 503444 1002489 503446 1002506
rect 503446 1002489 503498 1002506
rect 503498 1002489 503500 1002506
rect 503444 1002450 503500 1002489
rect 505076 1002319 505132 1002358
rect 505076 1002302 505078 1002319
rect 505078 1002302 505130 1002319
rect 505130 1002302 505132 1002319
rect 509396 1000691 509452 1000730
rect 509396 1000674 509398 1000691
rect 509398 1000674 509450 1000691
rect 509450 1000674 509452 1000691
rect 503060 999951 503116 999990
rect 503060 999934 503062 999951
rect 503062 999934 503114 999951
rect 503114 999934 503116 999951
rect 509876 999803 509932 999842
rect 509876 999786 509878 999803
rect 509878 999786 509930 999803
rect 509930 999786 509932 999803
rect 506228 999677 506230 999694
rect 506230 999677 506282 999694
rect 506282 999677 506284 999694
rect 506228 999638 506284 999677
rect 507764 999655 507820 999694
rect 507764 999638 507766 999655
rect 507766 999638 507818 999655
rect 507818 999638 507820 999655
rect 502388 999529 502390 999546
rect 502390 999529 502442 999546
rect 502442 999529 502444 999546
rect 502388 999490 502444 999529
rect 508628 999507 508684 999546
rect 508628 999490 508630 999507
rect 508630 999490 508682 999507
rect 508682 999490 508684 999507
rect 553748 1005153 553750 1005170
rect 553750 1005153 553802 1005170
rect 553802 1005153 553804 1005170
rect 553748 1005114 553804 1005153
rect 562484 1005153 562486 1005170
rect 562486 1005153 562538 1005170
rect 562538 1005153 562540 1005170
rect 562484 1005114 562540 1005153
rect 554900 1003821 554902 1003838
rect 554902 1003821 554954 1003838
rect 554954 1003821 554956 1003838
rect 554900 1003782 554956 1003821
rect 511124 996103 511180 996142
rect 511124 996086 511126 996103
rect 511126 996086 511178 996103
rect 511178 996086 511180 996103
rect 513428 996125 513430 996142
rect 513430 996125 513482 996142
rect 513482 996125 513484 996142
rect 513428 996086 513484 996125
rect 511892 995977 511894 995994
rect 511894 995977 511946 995994
rect 511946 995977 511948 995994
rect 511892 995938 511948 995977
rect 513332 995977 513334 995994
rect 513334 995977 513386 995994
rect 513386 995977 513388 995994
rect 513332 995938 513388 995977
rect 504692 995807 504748 995846
rect 504692 995790 504694 995807
rect 504694 995790 504746 995807
rect 504746 995790 504748 995807
rect 555668 1003673 555670 1003690
rect 555670 1003673 555722 1003690
rect 555722 1003673 555724 1003690
rect 555668 1003634 555724 1003673
rect 516692 1000230 516748 1000286
rect 516884 999786 516940 999842
rect 516788 999677 516790 999694
rect 516790 999677 516842 999694
rect 516842 999677 516844 999694
rect 516788 999638 516844 999677
rect 516788 999529 516790 999546
rect 516790 999529 516842 999546
rect 516842 999529 516844 999546
rect 516788 999490 516844 999529
rect 516692 999342 516748 999398
rect 517172 996086 517228 996142
rect 518516 995642 518572 995698
rect 518708 995642 518764 995698
rect 506612 995198 506668 995254
rect 509684 995050 509740 995106
rect 509876 994754 509932 994810
rect 518708 995494 518764 995550
rect 559124 1002489 559126 1002506
rect 559126 1002489 559178 1002506
rect 559178 1002489 559180 1002506
rect 559124 1002450 559180 1002489
rect 560564 1002467 560620 1002506
rect 560564 1002450 560566 1002467
rect 560566 1002450 560618 1002467
rect 560618 1002450 560620 1002467
rect 560084 1002341 560086 1002358
rect 560086 1002341 560138 1002358
rect 560138 1002341 560140 1002358
rect 560084 1002302 560140 1002341
rect 561524 1002319 561580 1002358
rect 564788 1002341 564790 1002358
rect 564790 1002341 564842 1002358
rect 564842 1002341 564844 1002358
rect 561524 1002302 561526 1002319
rect 561526 1002302 561578 1002319
rect 561578 1002302 561580 1002319
rect 523508 999786 523564 999842
rect 521396 995938 521452 995994
rect 519284 994902 519340 994958
rect 521588 995938 521644 995994
rect 521492 995494 521548 995550
rect 564788 1002302 564844 1002341
rect 523796 1000230 523852 1000286
rect 523700 999490 523756 999546
rect 523892 999638 523948 999694
rect 524084 999342 524140 999398
rect 523988 995790 524044 995846
rect 527924 995790 527980 995846
rect 532244 995790 532300 995846
rect 535316 995790 535372 995846
rect 552980 999381 552982 999398
rect 552982 999381 553034 999398
rect 553034 999381 553036 999398
rect 552980 999342 553036 999381
rect 557300 997879 557356 997918
rect 557300 997862 557302 997879
rect 557302 997862 557354 997879
rect 557354 997862 557356 997879
rect 558164 995790 558220 995846
rect 529076 995642 529132 995698
rect 534068 995642 534124 995698
rect 544244 995642 544300 995698
rect 526100 995346 526156 995402
rect 526484 995346 526540 995402
rect 530708 995346 530764 995402
rect 521684 995198 521740 995254
rect 526484 994902 526540 994958
rect 536852 995346 536908 995402
rect 537140 995198 537196 995254
rect 536852 994162 536908 994218
rect 562868 995938 562924 995994
rect 564788 995977 564790 995994
rect 564790 995977 564842 995994
rect 564842 995977 564844 995994
rect 564788 995938 564844 995977
rect 567092 995955 567148 995994
rect 567092 995938 567094 995955
rect 567094 995938 567146 995955
rect 567146 995938 567148 995955
rect 563732 995790 563788 995846
rect 566324 995807 566380 995846
rect 566324 995790 566326 995807
rect 566326 995790 566378 995807
rect 566378 995790 566380 995807
rect 561620 995346 561676 995402
rect 561428 994310 561484 994366
rect 570452 995050 570508 995106
rect 572852 994754 572908 994810
rect 573044 996382 573100 996438
rect 573140 995790 573196 995846
rect 572948 994458 573004 994514
rect 604820 996399 604876 996438
rect 604820 996382 604822 996399
rect 604822 996382 604874 996399
rect 604874 996382 604876 996399
rect 624884 995938 624940 995994
rect 634100 995790 634156 995846
rect 635828 995642 635884 995698
rect 581684 995385 581686 995402
rect 581686 995385 581738 995402
rect 581738 995385 581740 995402
rect 581684 995346 581740 995385
rect 584756 995198 584812 995254
rect 604724 995198 604780 995254
rect 575444 994902 575500 994958
rect 575348 994606 575404 994662
rect 629972 995050 630028 995106
rect 630932 994902 630988 994958
rect 631796 994754 631852 994810
rect 632372 994162 632428 994218
rect 634868 994310 634924 994366
rect 637364 994606 637420 994662
rect 638516 994606 638572 994662
rect 639188 994458 639244 994514
rect 640532 993866 640588 993922
rect 640916 994014 640972 994070
rect 641108 995050 641164 995106
rect 649844 994606 649900 994662
rect 82868 278434 82924 278490
rect 65204 245874 65260 245930
rect 71732 272810 71788 272866
rect 70580 272366 70636 272422
rect 69428 272218 69484 272274
rect 76532 272514 76588 272570
rect 74132 272070 74188 272126
rect 72980 266890 73036 266946
rect 78932 272662 78988 272718
rect 77780 269554 77836 269610
rect 83636 273254 83692 273310
rect 81332 272958 81388 273014
rect 86036 273106 86092 273162
rect 85268 269571 85324 269610
rect 85268 269554 85270 269571
rect 85270 269554 85322 269571
rect 85322 269554 85324 269571
rect 88436 273402 88492 273458
rect 90836 271626 90892 271682
rect 91988 271478 92044 271534
rect 87188 271330 87244 271386
rect 86516 269406 86572 269462
rect 90644 246614 90700 246670
rect 93236 271922 93292 271978
rect 96788 271774 96844 271830
rect 95636 271182 95692 271238
rect 100532 246614 100588 246670
rect 113492 276658 113548 276714
rect 116564 273550 116620 273606
rect 116564 271626 116620 271682
rect 116948 267778 117004 267834
rect 120500 276806 120556 276862
rect 118100 269850 118156 269906
rect 118100 269406 118156 269462
rect 121748 271626 121804 271682
rect 132500 266742 132556 266798
rect 140948 247502 141004 247558
rect 141140 269702 141196 269758
rect 141140 269554 141196 269610
rect 146900 273550 146956 273606
rect 143924 247650 143980 247706
rect 146708 247354 146764 247410
rect 146900 271626 146956 271682
rect 147092 271626 147148 271682
rect 146900 270738 146956 270794
rect 149588 247058 149644 247114
rect 146324 240546 146380 240602
rect 145556 236846 145612 236902
rect 144404 232110 144460 232166
rect 144020 226634 144076 226690
rect 144020 225006 144076 225062
rect 144116 223674 144172 223730
rect 144020 222934 144076 222990
rect 146420 235070 146476 235126
rect 144020 220122 144076 220178
rect 145364 218938 145420 218994
rect 144020 218198 144076 218254
rect 144116 215238 144172 215294
rect 144020 214498 144076 214554
rect 144116 209762 144172 209818
rect 144020 207433 144022 207450
rect 144022 207433 144074 207450
rect 144074 207433 144076 207450
rect 144020 207394 144076 207433
rect 144020 205618 144076 205674
rect 144020 203398 144076 203454
rect 144596 202066 144652 202122
rect 144116 201326 144172 201382
rect 144020 198958 144076 199014
rect 144020 197774 144076 197830
rect 144404 196590 144460 196646
rect 144308 194814 144364 194870
rect 144020 192890 144076 192946
rect 41780 184158 41836 184214
rect 41780 183566 41836 183622
rect 41780 182826 41836 182882
rect 144020 166546 144076 166602
rect 144020 162846 144076 162902
rect 144116 159886 144172 159942
rect 144020 159294 144076 159350
rect 144212 158110 144268 158166
rect 144116 156334 144172 156390
rect 144020 155759 144076 155798
rect 144020 155742 144022 155759
rect 144022 155742 144074 155759
rect 144074 155742 144076 155759
rect 144116 154410 144172 154466
rect 144020 152930 144076 152986
rect 144116 151598 144172 151654
rect 144020 150858 144076 150914
rect 143924 141238 143980 141294
rect 143828 138295 143884 138334
rect 143828 138278 143830 138295
rect 143830 138278 143882 138295
rect 143882 138278 143884 138295
rect 39860 125293 39862 125310
rect 39862 125293 39914 125310
rect 39914 125293 39916 125310
rect 39860 125254 39916 125293
rect 144212 147010 144268 147066
rect 144212 145974 144268 146030
rect 144212 144198 144268 144254
rect 144212 143162 144268 143218
rect 144212 142422 144268 142478
rect 144212 134726 144268 134782
rect 144212 133986 144268 134042
rect 144212 129990 144268 130046
rect 144116 104682 144172 104738
rect 144116 102758 144172 102814
rect 144020 101591 144076 101630
rect 144020 101574 144022 101591
rect 144022 101574 144074 101591
rect 144074 101574 144076 101591
rect 144116 99058 144172 99114
rect 144020 98061 144022 98078
rect 144022 98061 144074 98078
rect 144074 98061 144076 98078
rect 144020 98022 144076 98061
rect 144116 96246 144172 96302
rect 144020 95506 144076 95562
rect 144116 94322 144172 94378
rect 144020 92694 144076 92750
rect 144116 91362 144172 91418
rect 144020 89586 144076 89642
rect 144116 87810 144172 87866
rect 144020 75082 144076 75138
rect 144116 74934 144172 74990
rect 144116 72714 144172 72770
rect 144020 70938 144076 70994
rect 144020 69754 144076 69810
rect 144116 67386 144172 67442
rect 144020 62798 144076 62854
rect 144020 59581 144022 59598
rect 144022 59581 144074 59598
rect 144074 59581 144076 59598
rect 144020 59542 144076 59581
rect 144020 58654 144076 58710
rect 144020 57065 144022 57082
rect 144022 57065 144074 57082
rect 144074 57065 144076 57082
rect 144020 57026 144076 57065
rect 144020 56138 144076 56194
rect 144020 54675 144076 54714
rect 144020 54658 144022 54675
rect 144022 54658 144074 54675
rect 144074 54658 144076 54675
rect 144020 53770 144076 53826
rect 144500 185194 144556 185250
rect 144500 164770 144556 164826
rect 144500 147898 144556 147954
rect 144500 139462 144556 139518
rect 144500 132802 144556 132858
rect 144500 131026 144556 131082
rect 144692 180458 144748 180514
rect 145268 179718 145324 179774
rect 145268 176018 145324 176074
rect 145172 174390 145228 174446
rect 144884 172022 144940 172078
rect 144692 163586 144748 163642
rect 144788 161366 144844 161422
rect 144308 115042 144364 115098
rect 144596 115042 144652 115098
rect 144404 113118 144460 113174
rect 144404 111194 144460 111250
rect 144404 108234 144460 108290
rect 144308 105866 144364 105922
rect 144308 103646 144364 103702
rect 144308 99798 144364 99854
rect 144308 90770 144364 90826
rect 144692 106458 144748 106514
rect 144788 103942 144844 103998
rect 144404 80706 144460 80762
rect 144308 78634 144364 78690
rect 144308 77450 144364 77506
rect 144308 64574 144364 64630
rect 144596 83518 144652 83574
rect 144788 66202 144844 66258
rect 145076 170098 145132 170154
rect 144980 168322 145036 168378
rect 144980 65462 145036 65518
rect 144980 64574 145036 64630
rect 145460 216422 145516 216478
rect 145556 211686 145612 211742
rect 146708 238622 146764 238678
rect 146804 236271 146860 236310
rect 146804 236254 146806 236271
rect 146806 236254 146858 236271
rect 146858 236254 146860 236271
rect 146804 233590 146860 233646
rect 146804 231370 146860 231426
rect 146708 230186 146764 230242
rect 146804 229002 146860 229058
rect 146804 227670 146860 227726
rect 146420 213331 146476 213370
rect 146420 213314 146422 213331
rect 146422 213314 146474 213331
rect 146474 213314 146476 213331
rect 145748 210502 145804 210558
rect 145652 207986 145708 208042
rect 145844 205026 145900 205082
rect 146228 199550 146284 199606
rect 145940 193630 145996 193686
rect 146036 191706 146092 191762
rect 146228 190078 146284 190134
rect 146132 189338 146188 189394
rect 146036 73898 146092 73954
rect 146420 188154 146476 188210
rect 146420 186378 146476 186434
rect 146324 127474 146380 127530
rect 146324 125106 146380 125162
rect 146324 119038 146380 119094
rect 146324 84110 146380 84166
rect 146324 69014 146380 69070
rect 146612 183270 146668 183326
rect 146516 126734 146572 126790
rect 146516 115190 146572 115246
rect 146516 87070 146572 87126
rect 146804 184454 146860 184510
rect 146804 181790 146860 181846
rect 146804 178573 146806 178590
rect 146806 178573 146858 178590
rect 146858 178573 146860 178590
rect 146804 178534 146860 178573
rect 146804 176758 146860 176814
rect 146804 173354 146860 173410
rect 146804 171299 146860 171338
rect 146804 171282 146806 171299
rect 146806 171282 146858 171299
rect 146858 171282 146860 171299
rect 146804 167582 146860 167638
rect 146900 137538 146956 137594
rect 146900 136058 146956 136114
rect 146804 134430 146860 134486
rect 146804 132506 146860 132562
rect 146708 129250 146764 129306
rect 146708 124366 146764 124422
rect 146708 122590 146764 122646
rect 146708 120814 146764 120870
rect 146708 118446 146764 118502
rect 146708 116670 146764 116726
rect 146708 114154 146764 114210
rect 146708 112395 146764 112434
rect 146708 112378 146710 112395
rect 146710 112378 146762 112395
rect 146762 112378 146764 112395
rect 146708 109714 146764 109770
rect 146708 107494 146764 107550
rect 146708 85886 146764 85942
rect 146708 82334 146764 82390
rect 146708 79374 146764 79430
rect 146516 75674 146572 75730
rect 146516 74934 146572 74990
rect 146900 121406 146956 121462
rect 146900 115930 146956 115986
rect 147092 126899 147148 126938
rect 147092 126882 147094 126899
rect 147094 126882 147146 126899
rect 147146 126882 147148 126899
rect 146804 66350 146860 66406
rect 146900 62354 146956 62410
rect 146900 60726 146956 60782
rect 149108 149674 149164 149730
rect 155348 246910 155404 246966
rect 156884 273402 156940 273458
rect 156980 273254 157036 273310
rect 157172 273254 157228 273310
rect 156692 272662 156748 272718
rect 156884 272662 156940 272718
rect 156692 271034 156748 271090
rect 157172 271626 157228 271682
rect 156980 270886 157036 270942
rect 156884 247650 156940 247706
rect 156884 247206 156940 247262
rect 161108 247650 161164 247706
rect 158324 245282 158380 245338
rect 163988 245874 164044 245930
rect 157940 242322 157996 242378
rect 161204 242322 161260 242378
rect 161204 242026 161260 242082
rect 162740 237586 162796 237642
rect 161300 52159 161356 52198
rect 161300 52142 161302 52159
rect 161302 52142 161354 52159
rect 161354 52142 161356 52159
rect 166772 271626 166828 271682
rect 166772 270738 166828 270794
rect 166868 246022 166924 246078
rect 168596 245321 168598 245338
rect 168598 245321 168650 245338
rect 168650 245321 168652 245338
rect 168596 245282 168652 245321
rect 165524 48146 165580 48202
rect 171668 247206 171724 247262
rect 171764 246170 171820 246226
rect 172724 245726 172780 245782
rect 177044 273402 177100 273458
rect 177428 273254 177484 273310
rect 177044 272662 177100 272718
rect 177236 272662 177292 272718
rect 175508 245578 175564 245634
rect 171764 245282 171820 245338
rect 171668 245134 171724 245190
rect 171284 48590 171340 48646
rect 177716 273254 177772 273310
rect 177236 271034 177292 271090
rect 177428 271034 177484 271090
rect 177716 270886 177772 270942
rect 177044 246614 177100 246670
rect 177044 245874 177100 245930
rect 178388 245726 178444 245782
rect 174164 48442 174220 48498
rect 178580 270146 178636 270202
rect 178580 269702 178636 269758
rect 181364 245578 181420 245634
rect 181268 245430 181324 245486
rect 177044 48294 177100 48350
rect 168404 47850 168460 47906
rect 186836 245430 186892 245486
rect 187028 245430 187084 245486
rect 187028 244986 187084 245042
rect 187220 273550 187276 273606
rect 187220 271626 187276 271682
rect 188372 267482 188428 267538
rect 194516 273402 194572 273458
rect 187892 247058 187948 247114
rect 187700 246910 187756 246966
rect 187604 246762 187660 246818
rect 187988 246614 188044 246670
rect 187988 245282 188044 245338
rect 187700 245134 187756 245190
rect 188180 247206 188236 247262
rect 197588 273254 197644 273310
rect 197204 272662 197260 272718
rect 197204 271034 197260 271090
rect 197588 270886 197644 270942
rect 194516 270738 194572 270794
rect 195860 270146 195916 270202
rect 195956 269998 196012 270054
rect 207284 273550 207340 273606
rect 207284 271626 207340 271682
rect 201524 246949 201526 246966
rect 201526 246949 201578 246966
rect 201578 246949 201580 246966
rect 201524 246910 201580 246949
rect 202100 246466 202156 246522
rect 202196 245282 202252 245338
rect 202100 244690 202156 244746
rect 198932 239954 198988 240010
rect 204500 227670 204556 227726
rect 181364 52159 181420 52198
rect 181364 52142 181366 52159
rect 181366 52142 181418 52159
rect 181418 52142 181420 52159
rect 204884 232110 204940 232166
rect 204788 231518 204844 231574
rect 204692 230926 204748 230982
rect 205172 228262 205228 228318
rect 204884 226634 204940 226690
rect 204500 223970 204556 224026
rect 204596 222786 204652 222842
rect 204500 221158 204556 221214
rect 204596 219382 204652 219438
rect 204500 218494 204556 218550
rect 204596 217902 204652 217958
rect 204692 217754 204748 217810
rect 204788 215830 204844 215886
rect 204500 215238 204556 215294
rect 204980 221010 205036 221066
rect 204884 212870 204940 212926
rect 205268 226042 205324 226098
rect 205556 232258 205612 232314
rect 205460 225598 205516 225654
rect 205460 223378 205516 223434
rect 205364 220122 205420 220178
rect 205364 216866 205420 216922
rect 205652 227226 205708 227282
rect 205748 224414 205804 224470
rect 206996 266594 207052 266650
rect 211508 261848 211564 261904
rect 207284 255346 207340 255402
rect 205940 230482 205996 230538
rect 206132 229298 206188 229354
rect 204884 210206 204940 210262
rect 205076 210206 205132 210262
rect 206132 214646 206188 214702
rect 206420 221750 206476 221806
rect 206324 214498 206380 214554
rect 206516 213610 206572 213666
rect 206900 249870 206956 249926
rect 206804 229890 206860 229946
rect 206708 216274 206764 216330
rect 206612 213018 206668 213074
rect 206228 211982 206284 212038
rect 210548 245430 210604 245486
rect 207284 243358 207340 243414
rect 208724 239954 208780 240010
rect 208724 239066 208780 239122
rect 209876 239066 209932 239122
rect 209780 236698 209836 236754
rect 209684 236550 209740 236606
rect 207380 232110 207436 232166
rect 207092 229890 207148 229946
rect 206996 225006 207052 225062
rect 206900 222342 206956 222398
rect 206900 219530 206956 219586
rect 206804 211390 206860 211446
rect 205652 202658 205708 202714
rect 204500 102018 204556 102074
rect 204500 100390 204556 100446
rect 204596 100242 204652 100298
rect 204788 99354 204844 99410
rect 204692 98614 204748 98670
rect 204500 97765 204502 97782
rect 204502 97765 204554 97782
rect 204554 97765 204556 97782
rect 204500 97726 204556 97765
rect 204500 97134 204556 97190
rect 204500 94635 204556 94674
rect 204500 94618 204502 94635
rect 204502 94618 204554 94635
rect 204554 94618 204556 94635
rect 204596 93730 204652 93786
rect 204596 91954 204652 92010
rect 204500 91214 204556 91270
rect 204692 90622 204748 90678
rect 204596 90030 204652 90086
rect 204788 89586 204844 89642
rect 206708 101574 206764 101630
rect 206228 100982 206284 101038
rect 206900 98762 206956 98818
rect 206132 96986 206188 97042
rect 205268 96098 205324 96154
rect 206516 95506 206572 95562
rect 205748 94470 205804 94526
rect 205844 93878 205900 93934
rect 206900 92842 206956 92898
rect 206324 92250 206380 92306
rect 204500 88402 204556 88458
rect 204596 87958 204652 88014
rect 204788 88994 204844 89050
rect 204692 86774 204748 86830
rect 204500 86330 204556 86386
rect 204500 85738 204556 85794
rect 204596 84702 204652 84758
rect 204692 83518 204748 83574
rect 204500 83074 204556 83130
rect 204500 81890 204556 81946
rect 204500 80114 204556 80170
rect 204596 79226 204652 79282
rect 205268 87366 205324 87422
rect 205556 85146 205612 85202
rect 206612 84110 206668 84166
rect 205748 82482 205804 82538
rect 206708 81446 206764 81502
rect 206228 80854 206284 80910
rect 205268 80262 205324 80318
rect 204692 78634 204748 78690
rect 204788 77598 204844 77654
rect 204596 77006 204652 77062
rect 204500 75970 204556 76026
rect 204692 75230 204748 75286
rect 204500 74342 204556 74398
rect 204596 73602 204652 73658
rect 204692 72122 204748 72178
rect 204500 71695 204556 71734
rect 204500 71678 204502 71695
rect 204502 71678 204554 71695
rect 204554 71678 204556 71695
rect 204596 71086 204652 71142
rect 204980 69458 205036 69514
rect 205940 76858 205996 76914
rect 206516 75378 206572 75434
rect 205748 73750 205804 73806
rect 206804 72714 206860 72770
rect 205460 70494 205516 70550
rect 206804 69902 206860 69958
rect 204500 68866 204556 68922
rect 206420 68274 206476 68330
rect 204596 67830 204652 67886
rect 204116 67238 204172 67294
rect 206516 66646 206572 66702
rect 204500 66202 204556 66258
rect 206324 65610 206380 65666
rect 205460 65018 205516 65074
rect 204500 64574 204556 64630
rect 204596 63982 204652 64038
rect 204500 63407 204556 63446
rect 204500 63390 204502 63407
rect 204502 63390 204554 63407
rect 204554 63390 204556 63407
rect 204596 62946 204652 63002
rect 204692 62354 204748 62410
rect 204500 60726 204556 60782
rect 204884 61762 204940 61818
rect 204788 61318 204844 61374
rect 204500 60134 204556 60190
rect 206804 59986 206860 60042
rect 204596 59098 204652 59154
rect 206900 55842 206956 55898
rect 207956 230926 208012 230982
rect 207188 210206 207244 210262
rect 207284 190078 207340 190134
rect 207284 57618 207340 57674
rect 207092 53178 207148 53234
rect 209588 231518 209644 231574
rect 209396 230482 209452 230538
rect 209300 202658 209356 202714
rect 209204 57174 209260 57230
rect 209300 56582 209356 56638
rect 211412 246318 211468 246374
rect 211316 246170 211372 246226
rect 211124 246022 211180 246078
rect 211028 245874 211084 245930
rect 210740 245578 210796 245634
rect 211220 244690 211276 244746
rect 210932 236254 210988 236310
rect 210164 234774 210220 234830
rect 209972 55990 210028 56046
rect 209972 54732 210028 54788
rect 210164 228854 210220 228910
rect 210164 172614 210220 172670
rect 210164 152634 210220 152690
rect 210164 119038 210220 119094
rect 210164 94174 210220 94230
rect 210164 78116 210220 78172
rect 210260 54954 210316 55010
rect 211412 244690 211468 244746
rect 212564 273402 212620 273458
rect 211796 271330 211852 271386
rect 211604 246614 211660 246670
rect 211988 271182 212044 271238
rect 213044 272810 213100 272866
rect 212564 270738 212620 270794
rect 212756 270738 212812 270794
rect 216020 269889 216022 269906
rect 216022 269889 216074 269906
rect 216074 269889 216076 269906
rect 216020 269850 216076 269889
rect 217364 273254 217420 273310
rect 217364 270886 217420 270942
rect 227540 271626 227596 271682
rect 227540 271034 227596 271090
rect 237620 273402 237676 273458
rect 237524 272810 237580 272866
rect 237524 271330 237580 271386
rect 237716 273254 237772 273310
rect 237716 271330 237772 271386
rect 237620 271182 237676 271238
rect 243284 269889 243286 269906
rect 243286 269889 243338 269906
rect 243338 269889 243340 269906
rect 243284 269850 243340 269889
rect 247604 271626 247660 271682
rect 247604 271034 247660 271090
rect 248180 273550 248236 273606
rect 248180 272662 248236 272718
rect 249812 273994 249868 274050
rect 249140 273846 249196 273902
rect 250676 274142 250732 274198
rect 250580 273254 250636 273310
rect 250580 271330 250636 271386
rect 251828 274290 251884 274346
rect 252404 274438 252460 274494
rect 252020 268814 252076 268870
rect 253940 274586 253996 274642
rect 253364 269850 253420 269906
rect 253364 269702 253420 269758
rect 253364 269110 253420 269166
rect 252884 268962 252940 269018
rect 255092 273698 255148 273754
rect 254612 270294 254668 270350
rect 256436 270590 256492 270646
rect 256340 269406 256396 269462
rect 256148 267630 256204 267686
rect 256340 267334 256396 267390
rect 256820 267186 256876 267242
rect 257204 267038 257260 267094
rect 257684 273402 257740 273458
rect 257684 271182 257740 271238
rect 257876 270442 257932 270498
rect 258548 268518 258604 268574
rect 258356 267926 258412 267982
rect 259412 274734 259468 274790
rect 258932 268074 258988 268130
rect 260084 272810 260140 272866
rect 262676 276362 262732 276418
rect 262004 274882 262060 274938
rect 261140 271034 261196 271090
rect 260564 269554 260620 269610
rect 260660 268222 260716 268278
rect 261620 269258 261676 269314
rect 262868 276066 262924 276122
rect 263636 275918 263692 275974
rect 263732 275770 263788 275826
rect 264404 275622 264460 275678
rect 265460 275474 265516 275530
rect 264884 270886 264940 270942
rect 265076 268370 265132 268426
rect 265940 275178 265996 275234
rect 267668 275365 267670 275382
rect 267670 275365 267722 275382
rect 267722 275365 267724 275382
rect 267668 275326 267724 275365
rect 267860 275326 267916 275382
rect 266900 275030 266956 275086
rect 268148 275622 268204 275678
rect 268820 275474 268876 275530
rect 267860 271626 267916 271682
rect 267860 271330 267916 271386
rect 268148 269406 268204 269462
rect 267572 267334 267628 267390
rect 267764 267669 267766 267686
rect 267766 267669 267818 267686
rect 267818 267669 267820 267686
rect 267764 267630 267820 267669
rect 267860 267521 267862 267538
rect 267862 267521 267914 267538
rect 267914 267521 267916 267538
rect 267860 267482 267916 267521
rect 268052 267482 268108 267538
rect 269204 268666 269260 268722
rect 270644 271478 270700 271534
rect 276308 270590 276364 270646
rect 276596 270146 276652 270202
rect 276308 269850 276364 269906
rect 276500 269850 276556 269906
rect 287636 266759 287692 266798
rect 287636 266742 287638 266759
rect 287638 266742 287690 266759
rect 287690 266742 287692 266759
rect 287636 266594 287692 266650
rect 287924 266742 287980 266798
rect 287924 266594 287980 266650
rect 296564 270146 296620 270202
rect 296564 269850 296620 269906
rect 304532 278434 304588 278490
rect 299636 276214 299692 276270
rect 299492 269850 299548 269906
rect 299732 269702 299788 269758
rect 302420 271626 302476 271682
rect 303380 276510 303436 276566
rect 305204 278286 305260 278342
rect 305588 278138 305644 278194
rect 306356 277990 306412 278046
rect 307028 277842 307084 277898
rect 307796 277694 307852 277750
rect 309524 277546 309580 277602
rect 310388 277398 310444 277454
rect 311540 277250 311596 277306
rect 311636 277102 311692 277158
rect 313172 276954 313228 277010
rect 312116 270590 312172 270646
rect 312884 269998 312940 270054
rect 315764 271478 315820 271534
rect 317492 269998 317548 270054
rect 317492 269850 317548 269906
rect 318164 269406 318220 269462
rect 320180 276362 320236 276418
rect 319124 270146 319180 270202
rect 318740 269998 318796 270054
rect 322484 276214 322540 276270
rect 322676 276214 322732 276270
rect 322484 271330 322540 271386
rect 322580 271182 322636 271238
rect 320564 270590 320620 270646
rect 322484 270590 322540 270646
rect 320852 269406 320908 269462
rect 324404 271626 324460 271682
rect 323252 271330 323308 271386
rect 323252 269998 323308 270054
rect 323156 269702 323212 269758
rect 322772 268666 322828 268722
rect 323444 269998 323500 270054
rect 324404 269406 324460 269462
rect 324980 271478 325036 271534
rect 325364 271478 325420 271534
rect 325460 271034 325516 271090
rect 325652 271073 325654 271090
rect 325654 271073 325706 271090
rect 325706 271073 325708 271090
rect 324692 269850 324748 269906
rect 325652 271034 325708 271073
rect 325460 269406 325516 269462
rect 324596 268666 324652 268722
rect 327092 269850 327148 269906
rect 328820 271626 328876 271682
rect 329012 271626 329068 271682
rect 327956 271182 328012 271238
rect 328148 271182 328204 271238
rect 328052 270590 328108 270646
rect 328628 271034 328684 271090
rect 328820 271034 328876 271090
rect 328628 270590 328684 270646
rect 329012 269998 329068 270054
rect 328436 269850 328492 269906
rect 328820 269406 328876 269462
rect 329012 269406 329068 269462
rect 328628 268666 328684 268722
rect 328820 268666 328876 268722
rect 328436 267778 328492 267834
rect 328052 267038 328108 267094
rect 328340 267038 328396 267094
rect 328436 266890 328492 266946
rect 328628 266890 328684 266946
rect 328532 266594 328588 266650
rect 329300 266594 329356 266650
rect 325460 264929 325516 264985
rect 330836 271182 330892 271238
rect 336596 269702 336652 269758
rect 336980 271330 337036 271386
rect 336980 270146 337036 270202
rect 372884 278582 372940 278638
rect 339764 271182 339820 271238
rect 342452 271034 342508 271090
rect 342548 269850 342604 269906
rect 347828 266890 347884 266946
rect 347732 266594 347788 266650
rect 348788 267778 348844 267834
rect 348980 267778 349036 267834
rect 348500 266890 348556 266946
rect 348788 266890 348844 266946
rect 348692 266742 348748 266798
rect 349076 266594 349132 266650
rect 349364 267038 349420 267094
rect 349844 266594 349900 266650
rect 351284 270886 351340 270942
rect 355220 270738 355276 270794
rect 356948 270886 357004 270942
rect 356948 268074 357004 268130
rect 357812 267778 357868 267834
rect 363764 271330 363820 271386
rect 368180 271034 368236 271090
rect 368180 268074 368236 268130
rect 370004 274882 370060 274938
rect 368468 274734 368524 274790
rect 369140 273441 369142 273458
rect 369142 273441 369194 273458
rect 369194 273441 369196 273458
rect 369140 273402 369196 273441
rect 368660 272662 368716 272718
rect 368852 272662 368908 272718
rect 368372 270738 368428 270794
rect 368756 270738 368812 270794
rect 368948 270738 369004 270794
rect 368564 269702 368620 269758
rect 368756 269702 368812 269758
rect 368372 268222 368428 268278
rect 368756 268074 368812 268130
rect 369236 268222 369292 268278
rect 368756 267038 368812 267094
rect 368468 266890 368524 266946
rect 368372 266594 368428 266650
rect 365012 264929 365068 264985
rect 368660 266890 368716 266946
rect 370388 274734 370444 274790
rect 370964 271478 371020 271534
rect 370580 271330 370636 271386
rect 369812 271034 369868 271090
rect 369812 270442 369868 270498
rect 370004 270442 370060 270498
rect 370580 268518 370636 268574
rect 370772 268518 370828 268574
rect 371444 271478 371500 271534
rect 372404 274586 372460 274642
rect 371444 270886 371500 270942
rect 371444 268518 371500 268574
rect 372692 267778 372748 267834
rect 373172 270738 373228 270794
rect 374324 278582 374380 278638
rect 373556 270738 373612 270794
rect 375188 276806 375244 276862
rect 375380 276806 375436 276862
rect 375284 276658 375340 276714
rect 375476 276658 375532 276714
rect 374996 272218 375052 272274
rect 374516 271922 374572 271978
rect 374132 267186 374188 267242
rect 374420 267225 374422 267242
rect 374422 267225 374474 267242
rect 374474 267225 374476 267242
rect 374420 267186 374476 267225
rect 374612 267186 374668 267242
rect 376340 273106 376396 273162
rect 376532 273106 376588 273162
rect 376628 270886 376684 270942
rect 377108 267926 377164 267982
rect 376820 267778 376876 267834
rect 376820 267482 376876 267538
rect 395060 278582 395116 278638
rect 378836 274882 378892 274938
rect 377972 273550 378028 273606
rect 378164 273550 378220 273606
rect 377396 267926 377452 267982
rect 379700 273550 379756 273606
rect 379028 273254 379084 273310
rect 378932 272958 378988 273014
rect 379220 273402 379276 273458
rect 379412 273402 379468 273458
rect 379316 273106 379372 273162
rect 379220 272958 379276 273014
rect 379316 272218 379372 272274
rect 379316 271626 379372 271682
rect 378740 267482 378796 267538
rect 379796 272218 379852 272274
rect 380180 272218 380236 272274
rect 380180 269702 380236 269758
rect 380564 269702 380620 269758
rect 381236 273698 381292 273754
rect 381812 273402 381868 273458
rect 381620 272366 381676 272422
rect 381812 272366 381868 272422
rect 381812 272070 381868 272126
rect 383348 273698 383404 273754
rect 383540 273698 383596 273754
rect 383252 273550 383308 273606
rect 383156 273402 383212 273458
rect 383540 272514 383596 272570
rect 383348 272070 383404 272126
rect 383444 271922 383500 271978
rect 383156 269850 383212 269906
rect 384404 273106 384460 273162
rect 384788 273106 384844 273162
rect 383924 272514 383980 272570
rect 383636 271922 383692 271978
rect 383924 270738 383980 270794
rect 384884 272070 384940 272126
rect 386132 272366 386188 272422
rect 385556 271922 385612 271978
rect 386036 270886 386092 270942
rect 387092 272514 387148 272570
rect 386612 272366 386668 272422
rect 388052 271626 388108 271682
rect 387572 270738 387628 270794
rect 387764 270755 387820 270794
rect 387764 270738 387766 270755
rect 387766 270738 387818 270755
rect 387818 270738 387820 270755
rect 388724 276658 388780 276714
rect 389012 272514 389068 272570
rect 389204 271774 389260 271830
rect 388628 271626 388684 271682
rect 388916 271665 388918 271682
rect 388918 271665 388970 271682
rect 388970 271665 388972 271682
rect 388916 271626 388972 271665
rect 388724 270442 388780 270498
rect 388916 270442 388972 270498
rect 389012 268074 389068 268130
rect 388916 267482 388972 267538
rect 388820 266890 388876 266946
rect 388628 266594 388684 266650
rect 389684 273698 389740 273754
rect 389684 273106 389740 273162
rect 389972 272531 390028 272570
rect 389972 272514 389974 272531
rect 389974 272514 390026 272531
rect 390026 272514 390028 272531
rect 389396 268370 389452 268426
rect 390836 271626 390892 271682
rect 391412 271774 391468 271830
rect 391028 267778 391084 267834
rect 393716 276806 393772 276862
rect 474740 278434 474796 278490
rect 481844 278286 481900 278342
rect 485396 278138 485452 278194
rect 488948 277990 489004 278046
rect 393908 268518 393964 268574
rect 394100 268518 394156 268574
rect 393716 268074 393772 268130
rect 393908 268074 393964 268130
rect 394676 273106 394732 273162
rect 394580 270738 394636 270794
rect 395348 272958 395404 273014
rect 395828 270738 395884 270794
rect 396884 267926 396940 267982
rect 396596 267334 396652 267390
rect 396788 267351 396844 267390
rect 396788 267334 396790 267351
rect 396790 267334 396842 267351
rect 396842 267334 396844 267351
rect 397172 267334 397228 267390
rect 398900 269702 398956 269758
rect 398900 268518 398956 268574
rect 399284 266594 399340 266650
rect 399476 266594 399532 266650
rect 400532 268370 400588 268426
rect 400532 267926 400588 267982
rect 400148 266594 400204 266650
rect 400436 266594 400492 266650
rect 401108 268370 401164 268426
rect 401204 266594 401260 266650
rect 401588 270886 401644 270942
rect 403124 269850 403180 269906
rect 402452 266594 402508 266650
rect 403220 266594 403276 266650
rect 403892 266594 403948 266650
rect 404756 266594 404812 266650
rect 405236 266594 405292 266650
rect 406100 269702 406156 269758
rect 406196 266594 406252 266650
rect 406580 266594 406636 266650
rect 409172 274586 409228 274642
rect 409172 273698 409228 273754
rect 406868 266611 406924 266650
rect 406868 266594 406870 266611
rect 406870 266594 406922 266611
rect 406922 266594 406924 266611
rect 407156 266594 407212 266650
rect 407348 266594 407404 266650
rect 408596 267778 408652 267834
rect 408788 267778 408844 267834
rect 408500 266907 408556 266946
rect 408500 266890 408502 266907
rect 408502 266890 408554 266907
rect 408554 266890 408556 266907
rect 408692 267482 408748 267538
rect 408884 267482 408940 267538
rect 408788 266890 408844 266946
rect 408788 266594 408844 266650
rect 409076 266611 409132 266650
rect 409076 266594 409078 266611
rect 409078 266594 409130 266611
rect 409130 266594 409132 266611
rect 409460 266594 409516 266650
rect 409652 266594 409708 266650
rect 413780 266298 413836 266354
rect 414740 269850 414796 269906
rect 427604 269889 427606 269906
rect 427606 269889 427658 269906
rect 427658 269889 427660 269906
rect 427604 269850 427660 269889
rect 419156 266890 419212 266946
rect 419348 266890 419404 266946
rect 419156 266594 419212 266650
rect 419348 266298 419404 266354
rect 413684 266150 413740 266206
rect 429140 276066 429196 276122
rect 429044 274586 429100 274642
rect 428948 273698 429004 273754
rect 429236 274625 429238 274642
rect 429238 274625 429290 274642
rect 429290 274625 429292 274642
rect 429236 274586 429292 274625
rect 429140 273698 429196 273754
rect 429140 270442 429196 270498
rect 429140 268370 429196 268426
rect 434804 269702 434860 269758
rect 437588 269889 437590 269906
rect 437590 269889 437642 269906
rect 437642 269889 437644 269906
rect 437588 269850 437644 269889
rect 439124 266742 439180 266798
rect 439028 266298 439084 266354
rect 413396 265854 413452 265910
rect 413204 265706 413260 265762
rect 439220 266594 439276 266650
rect 439124 266002 439180 266058
rect 439316 266150 439372 266206
rect 439220 265854 439276 265910
rect 439028 265558 439084 265614
rect 449204 276066 449260 276122
rect 449108 274625 449110 274642
rect 449110 274625 449162 274642
rect 449162 274625 449164 274642
rect 449108 274586 449164 274625
rect 449204 273698 449260 273754
rect 449204 270442 449260 270498
rect 449204 268370 449260 268426
rect 457940 269702 457996 269758
rect 458612 269702 458668 269758
rect 459284 266742 459340 266798
rect 458132 266298 458188 266354
rect 459380 266594 459436 266650
rect 459284 266002 459340 266058
rect 459380 265854 459436 265910
rect 459572 265854 459628 265910
rect 458132 265558 458188 265614
rect 467828 276510 467884 276566
rect 469460 276066 469516 276122
rect 469556 274586 469612 274642
rect 469460 273698 469516 273754
rect 469460 270442 469516 270498
rect 469364 269850 469420 269906
rect 469556 269850 469612 269906
rect 469460 269702 469516 269758
rect 477428 273846 477484 273902
rect 477620 273846 477676 273902
rect 484436 273994 484492 274050
rect 483860 269702 483916 269758
rect 483860 269554 483916 269610
rect 484148 269554 484204 269610
rect 489524 276066 489580 276122
rect 489428 274586 489484 274642
rect 489428 273846 489484 273902
rect 489524 273698 489580 273754
rect 491636 274142 491692 274198
rect 489524 270442 489580 270498
rect 489428 269850 489484 269906
rect 486740 268074 486796 268130
rect 480980 267926 481036 267982
rect 479348 266742 479404 266798
rect 479540 266742 479596 266798
rect 479444 266594 479500 266650
rect 479636 266594 479692 266650
rect 479540 266298 479596 266354
rect 479444 266150 479500 266206
rect 479348 266002 479404 266058
rect 479636 265854 479692 265910
rect 496148 277842 496204 277898
rect 498836 274142 498892 274198
rect 497684 265854 497740 265910
rect 439316 265410 439372 265466
rect 413204 265262 413260 265318
rect 455060 265262 455116 265318
rect 401588 264929 401644 264985
rect 412532 264966 412588 265022
rect 459572 265410 459628 265466
rect 503252 277694 503308 277750
rect 504404 274586 504460 274642
rect 504404 274142 504460 274198
rect 505940 274438 505996 274494
rect 502292 268814 502348 268870
rect 505268 266446 505324 266502
rect 501236 266150 501292 266206
rect 475124 265114 475180 265170
rect 483860 265114 483916 265170
rect 509780 276066 509836 276122
rect 509780 274438 509836 274494
rect 509780 270442 509836 270498
rect 509492 268962 509548 269018
rect 509780 268962 509836 269018
rect 513044 269110 513100 269166
rect 517748 277546 517804 277602
rect 518324 269741 518326 269758
rect 518326 269741 518378 269758
rect 518378 269741 518380 269758
rect 518324 269702 518380 269741
rect 511124 265114 511180 265170
rect 524948 277398 525004 277454
rect 524372 270442 524428 270498
rect 523796 270294 523852 270350
rect 524372 268962 524428 269018
rect 529844 276066 529900 276122
rect 529844 274438 529900 274494
rect 529940 269850 529996 269906
rect 529844 269702 529900 269758
rect 528500 267778 528556 267834
rect 532148 277250 532204 277306
rect 530900 267630 530956 267686
rect 535604 277102 535660 277158
rect 538004 267482 538060 267538
rect 534452 267334 534508 267390
rect 541556 267186 541612 267242
rect 546356 276954 546412 277010
rect 545684 276066 545740 276122
rect 545684 274438 545740 274494
rect 548756 271034 548812 271090
rect 545204 267038 545260 267094
rect 542804 266890 542860 266946
rect 521396 264966 521452 265022
rect 552980 274181 552982 274198
rect 552982 274181 553034 274198
rect 553034 274181 553036 274198
rect 552980 274142 553036 274181
rect 555860 271330 555916 271386
rect 552308 271182 552364 271238
rect 552980 270459 553036 270498
rect 552980 270442 552982 270459
rect 552982 270442 553034 270459
rect 553034 270442 553036 270459
rect 552980 269850 553036 269906
rect 553076 269702 553132 269758
rect 559412 271478 559468 271534
rect 563060 272662 563116 272718
rect 566516 272810 566572 272866
rect 570068 276066 570124 276122
rect 570068 274438 570124 274494
rect 570164 269554 570220 269610
rect 573044 274290 573100 274346
rect 573716 272218 573772 272274
rect 573044 270294 573100 270350
rect 573140 270146 573196 270202
rect 573140 269571 573196 269610
rect 573140 269554 573142 269571
rect 573142 269554 573194 269571
rect 573194 269554 573196 269571
rect 584756 274438 584812 274494
rect 584564 274290 584620 274346
rect 584372 273254 584428 273310
rect 582068 270590 582124 270646
rect 587924 276066 587980 276122
rect 591572 275918 591628 275974
rect 593300 274455 593356 274494
rect 593300 274438 593302 274455
rect 593302 274438 593354 274455
rect 593354 274438 593356 274455
rect 590420 270459 590476 270498
rect 590420 270442 590422 270459
rect 590422 270442 590474 270459
rect 590474 270442 590476 270459
rect 595124 275770 595180 275826
rect 598772 275622 598828 275678
rect 603380 276362 603436 276418
rect 602228 275474 602284 275530
rect 605780 273402 605836 273458
rect 600500 270459 600556 270498
rect 600500 270442 600502 270459
rect 600502 270442 600554 270459
rect 600554 270442 600556 270459
rect 596372 269998 596428 270054
rect 593204 269702 593260 269758
rect 580916 269258 580972 269314
rect 577268 268666 577324 268722
rect 610580 269702 610636 269758
rect 607028 265114 607084 265170
rect 612980 275326 613036 275382
rect 613364 274455 613420 274494
rect 613364 274438 613366 274455
rect 613366 274438 613418 274455
rect 613418 274438 613420 274455
rect 616532 275178 616588 275234
rect 619124 274290 619180 274346
rect 620564 275178 620620 275234
rect 620564 274734 620620 274790
rect 624884 276214 624940 276270
rect 623636 275030 623692 275086
rect 620084 268518 620140 268574
rect 632084 269406 632140 269462
rect 630836 268222 630892 268278
rect 637940 275178 637996 275234
rect 645140 274882 645196 274938
rect 642740 266742 642796 266798
rect 648692 273550 648748 273606
rect 647540 270738 647596 270794
rect 649556 941770 649612 941826
rect 646292 266594 646348 266650
rect 635540 265706 635596 265762
rect 216884 246762 216940 246818
rect 212084 244542 212140 244598
rect 211892 233738 211948 233794
rect 211028 233590 211084 233646
rect 211316 233590 211372 233646
rect 211700 233590 211756 233646
rect 211412 233442 211468 233498
rect 212180 233590 212236 233646
rect 212372 243654 212428 243710
rect 213236 235070 213292 235126
rect 214292 243506 214348 243562
rect 214868 237734 214924 237790
rect 214292 233442 214348 233498
rect 227924 246762 227980 246818
rect 215828 238030 215884 238086
rect 215252 237882 215308 237938
rect 214964 234922 215020 234978
rect 215924 237586 215980 237642
rect 218228 243802 218284 243858
rect 217172 235810 217228 235866
rect 219764 243950 219820 244006
rect 219188 235218 219244 235274
rect 221012 244394 221068 244450
rect 220820 235514 220876 235570
rect 223028 242914 223084 242970
rect 222164 235366 222220 235422
rect 224564 243062 224620 243118
rect 225812 244098 225868 244154
rect 226388 244690 226444 244746
rect 223988 235662 224044 235718
rect 227060 245025 227062 245042
rect 227062 245025 227114 245042
rect 227114 245025 227116 245042
rect 227060 244986 227116 245025
rect 227444 244690 227500 244746
rect 227636 244729 227638 244746
rect 227638 244729 227690 244746
rect 227690 244729 227692 244746
rect 227636 244690 227692 244729
rect 227540 244542 227596 244598
rect 246452 246762 246508 246818
rect 247796 246762 247852 246818
rect 248372 246762 248428 246818
rect 228116 244986 228172 245042
rect 228212 244690 228268 244746
rect 229556 244542 229612 244598
rect 228596 236106 228652 236162
rect 229748 235958 229804 236014
rect 232340 243210 232396 243266
rect 235700 242026 235756 242082
rect 240980 240546 241036 240602
rect 241364 238178 241420 238234
rect 241748 240694 241804 240750
rect 242324 238326 242380 238382
rect 243188 241138 243244 241194
rect 242708 240990 242764 241046
rect 242804 238622 242860 238678
rect 243572 238770 243628 238826
rect 243956 241286 244012 241342
rect 244340 238918 244396 238974
rect 245396 241730 245452 241786
rect 246164 241878 246220 241934
rect 247508 244986 247564 245042
rect 247700 244986 247756 245042
rect 247508 244690 247564 244746
rect 247700 244690 247756 244746
rect 259220 246762 259276 246818
rect 247124 240250 247180 240306
rect 247604 240102 247660 240158
rect 257684 244690 257740 244746
rect 257588 244246 257644 244302
rect 257684 244098 257740 244154
rect 257876 244098 257932 244154
rect 257588 243062 257644 243118
rect 257876 242914 257932 242970
rect 267956 246762 268012 246818
rect 258644 240842 258700 240898
rect 259988 241582 260044 241638
rect 259604 241434 259660 241490
rect 259028 238474 259084 238530
rect 262580 239954 262636 240010
rect 291956 246762 292012 246818
rect 292148 246762 292204 246818
rect 272948 234478 273004 234534
rect 282548 242174 282604 242230
rect 282260 240398 282316 240454
rect 283220 242322 283276 242378
rect 285140 242618 285196 242674
rect 286868 236846 286924 236902
rect 286772 234330 286828 234386
rect 287924 244986 287980 245042
rect 288116 244986 288172 245042
rect 290036 244986 290092 245042
rect 307988 246762 308044 246818
rect 289364 236271 289420 236310
rect 289364 236254 289366 236271
rect 289366 236254 289418 236271
rect 289418 236254 289420 236271
rect 290708 242470 290764 242526
rect 290804 242361 290806 242378
rect 290806 242361 290858 242378
rect 290858 242361 290860 242378
rect 290804 242322 290860 242361
rect 292340 244986 292396 245042
rect 292436 242213 292438 242230
rect 292438 242213 292490 242230
rect 292490 242213 292492 242230
rect 292436 242174 292492 242213
rect 293780 236254 293836 236310
rect 296660 243062 296716 243118
rect 297236 243062 297292 243118
rect 296756 242914 296812 242970
rect 295892 236846 295948 236902
rect 297524 242322 297580 242378
rect 297908 242618 297964 242674
rect 298196 242470 298252 242526
rect 298004 242322 298060 242378
rect 297428 234330 297484 234386
rect 311156 246779 311212 246818
rect 311156 246762 311158 246779
rect 311158 246762 311210 246779
rect 311210 246762 311212 246779
rect 327092 246762 327148 246818
rect 327956 246762 328012 246818
rect 328340 246762 328396 246818
rect 328532 246762 328588 246818
rect 305780 242914 305836 242970
rect 307796 244986 307852 245042
rect 307988 244986 308044 245042
rect 308180 244986 308236 245042
rect 308084 244394 308140 244450
rect 308276 244394 308332 244450
rect 308180 243062 308236 243118
rect 309428 244986 309484 245042
rect 321908 237438 321964 237494
rect 322292 237307 322348 237346
rect 322292 237290 322294 237307
rect 322294 237290 322346 237307
rect 322346 237290 322348 237307
rect 322772 237307 322828 237346
rect 322772 237290 322774 237307
rect 322774 237290 322826 237307
rect 322826 237290 322828 237307
rect 326804 244986 326860 245042
rect 328244 244986 328300 245042
rect 328436 244986 328492 245042
rect 328628 244986 328684 245042
rect 328724 244394 328780 244450
rect 328436 243506 328492 243562
rect 328436 242914 328492 242970
rect 335156 243654 335212 243710
rect 335348 237438 335404 237494
rect 348116 246779 348172 246818
rect 348116 246762 348118 246779
rect 348118 246762 348170 246779
rect 348170 246762 348172 246779
rect 348596 246779 348652 246818
rect 348596 246762 348598 246779
rect 348598 246762 348650 246779
rect 348650 246762 348652 246779
rect 367604 246762 367660 246818
rect 367988 246762 368044 246818
rect 369428 246762 369484 246818
rect 338996 235810 339052 235866
rect 341108 243802 341164 243858
rect 341588 243950 341644 244006
rect 341204 235218 341260 235274
rect 342548 243062 342604 243118
rect 342164 235514 342220 235570
rect 343316 244098 343372 244154
rect 342932 235366 342988 235422
rect 343796 244246 343852 244302
rect 343412 235662 343468 235718
rect 344468 244690 344524 244746
rect 344372 235070 344428 235126
rect 346004 243506 346060 243562
rect 345620 236106 345676 236162
rect 346580 235958 346636 236014
rect 347732 243210 347788 243266
rect 348212 244986 348268 245042
rect 348596 244690 348652 244746
rect 348404 244542 348460 244598
rect 348404 242914 348460 242970
rect 348884 244986 348940 245042
rect 348884 242026 348940 242082
rect 351380 239066 351436 239122
rect 352244 240102 352300 240158
rect 352244 234922 352300 234978
rect 353972 240250 354028 240306
rect 354452 234478 354508 234534
rect 355028 241878 355084 241934
rect 356756 241730 356812 241786
rect 360020 241286 360076 241342
rect 358964 238918 359020 238974
rect 359252 236550 359308 236606
rect 360692 238770 360748 238826
rect 361556 241138 361612 241194
rect 363092 240990 363148 241046
rect 362708 238622 362764 238678
rect 363860 238326 363916 238382
rect 364820 240694 364876 240750
rect 365780 238178 365836 238234
rect 366548 240546 366604 240602
rect 367604 240546 367660 240602
rect 368372 244986 368428 245042
rect 368468 244542 368524 244598
rect 368564 244394 368620 244450
rect 369908 246779 369964 246818
rect 369908 246762 369910 246779
rect 369910 246762 369962 246779
rect 369962 246762 369964 246779
rect 370196 246762 370252 246818
rect 370676 246762 370732 246818
rect 377204 246762 377260 246818
rect 369044 244986 369100 245042
rect 369140 244690 369196 244746
rect 368852 244542 368908 244598
rect 369140 244098 369196 244154
rect 388244 246762 388300 246818
rect 376148 241582 376204 241638
rect 370964 239954 371020 240010
rect 376820 241434 376876 241490
rect 392564 246762 392620 246818
rect 392948 246762 393004 246818
rect 378836 240842 378892 240898
rect 377684 238474 377740 238530
rect 379412 234774 379468 234830
rect 383060 241730 383116 241786
rect 383060 240119 383116 240158
rect 383060 240102 383062 240119
rect 383062 240102 383114 240119
rect 383114 240102 383116 240119
rect 383060 239971 383116 240010
rect 383060 239954 383062 239971
rect 383062 239954 383114 239971
rect 383114 239954 383116 239971
rect 383060 239066 383116 239122
rect 383060 238661 383062 238678
rect 383062 238661 383114 238678
rect 383114 238661 383116 238678
rect 383060 238622 383116 238661
rect 385268 243358 385324 243414
rect 388532 244986 388588 245042
rect 388724 244986 388780 245042
rect 388532 244690 388588 244746
rect 389012 244986 389068 245042
rect 389876 240102 389932 240158
rect 391412 238030 391468 238086
rect 393428 246762 393484 246818
rect 393140 237882 393196 237938
rect 395348 238622 395404 238678
rect 394676 237734 394732 237790
rect 400916 244690 400972 244746
rect 401492 244986 401548 245042
rect 403316 244986 403372 245042
rect 403892 244690 403948 244746
rect 403796 244542 403852 244598
rect 404372 244986 404428 245042
rect 404372 244707 404428 244746
rect 404372 244690 404374 244707
rect 404374 244690 404426 244707
rect 404426 244690 404428 244707
rect 405140 244986 405196 245042
rect 402356 239954 402412 240010
rect 407060 244986 407116 245042
rect 409172 244986 409228 245042
rect 409748 240546 409804 240602
rect 411476 240398 411532 240454
rect 411956 237586 412012 237642
rect 509780 242174 509836 242230
rect 504020 242026 504076 242082
rect 497492 236698 497548 236754
rect 420596 236402 420652 236458
rect 541460 234626 541516 234682
rect 637076 233590 637132 233646
rect 637556 233442 637612 233498
rect 638132 233738 638188 233794
rect 638708 233738 638764 233794
rect 637940 233442 637996 233498
rect 638516 233590 638572 233646
rect 638996 233442 639052 233498
rect 649652 801318 649708 801374
rect 212372 54214 212428 54270
rect 214388 54214 214444 54270
rect 214772 54066 214828 54122
rect 216596 53918 216652 53974
rect 209492 48886 209548 48942
rect 187604 41782 187660 41838
rect 194324 41782 194380 41838
rect 211892 51846 211948 51902
rect 212084 45038 212140 45094
rect 212660 51994 212716 52050
rect 213044 53474 213100 53530
rect 212852 44890 212908 44946
rect 215252 53326 215308 53382
rect 215924 53474 215980 53530
rect 216020 53069 216022 53086
rect 216022 53069 216074 53086
rect 216074 53069 216076 53086
rect 216020 53030 216076 53069
rect 216980 53770 217036 53826
rect 216788 53474 216844 53530
rect 220004 53474 220060 53530
rect 220340 53178 220396 53234
rect 220724 48886 220780 48942
rect 221876 51698 221932 51754
rect 222548 52142 222604 52198
rect 223316 51550 223372 51606
rect 229652 50366 229708 50422
rect 238196 51254 238252 51310
rect 242036 48590 242092 48646
rect 241940 48146 241996 48202
rect 243380 51402 243436 51458
rect 242996 48442 243052 48498
rect 243764 48294 243820 48350
rect 242612 47850 242668 47906
rect 302516 43262 302572 43318
rect 302324 42078 302380 42134
rect 306740 42078 306796 42134
rect 416564 43262 416620 43318
rect 466580 46074 466636 46130
rect 361460 41782 361516 41838
rect 364628 41782 364684 41838
rect 328052 40894 328108 40950
rect 210740 40746 210796 40802
rect 327284 40746 327340 40802
rect 461108 43114 461164 43170
rect 465620 43114 465676 43170
rect 471092 42078 471148 42134
rect 463700 41782 463756 41838
rect 645716 232406 645772 232462
rect 645140 232297 645142 232314
rect 645142 232297 645194 232314
rect 645194 232297 645196 232314
rect 645140 232258 645196 232297
rect 645140 231557 645142 231574
rect 645142 231557 645194 231574
rect 645194 231557 645196 231574
rect 645140 231518 645196 231557
rect 645140 231113 645142 231130
rect 645142 231113 645194 231130
rect 645194 231113 645196 231130
rect 645140 231074 645196 231113
rect 645140 230669 645142 230686
rect 645142 230669 645194 230686
rect 645194 230669 645196 230686
rect 645140 230630 645196 230669
rect 517844 43262 517900 43318
rect 520628 43262 520684 43318
rect 526964 42078 527020 42134
rect 528980 42078 529036 42134
rect 645428 78486 645484 78542
rect 645620 210354 645676 210410
rect 649748 707486 649804 707542
rect 650036 895150 650092 895206
rect 650132 848234 650188 848290
rect 649940 754550 649996 754606
rect 649844 660570 649900 660626
rect 655124 976698 655180 976754
rect 654452 953314 654508 953370
rect 655220 965006 655276 965062
rect 674324 967522 674380 967578
rect 674996 967522 675052 967578
rect 674516 967374 674572 967430
rect 675764 966338 675820 966394
rect 675668 965746 675724 965802
rect 675188 964858 675244 964914
rect 675764 963230 675820 963286
rect 675092 962490 675148 962546
rect 675092 962194 675148 962250
rect 675380 961454 675436 961510
rect 675380 961306 675436 961362
rect 675476 960122 675532 960178
rect 675764 959086 675820 959142
rect 654452 929782 654508 929838
rect 653972 918090 654028 918146
rect 654452 906398 654508 906454
rect 653972 882866 654028 882922
rect 654452 871174 654508 871230
rect 654164 859482 654220 859538
rect 653972 835950 654028 836006
rect 653972 824258 654028 824314
rect 654452 812566 654508 812622
rect 654068 789034 654124 789090
rect 654068 777342 654124 777398
rect 653972 765502 654028 765558
rect 653972 742118 654028 742174
rect 655220 730426 655276 730482
rect 654260 718586 654316 718642
rect 654452 695202 654508 695258
rect 654452 671670 654508 671726
rect 654260 648286 654316 648342
rect 654356 624754 654412 624810
rect 654356 613062 654412 613118
rect 654452 601370 654508 601426
rect 655124 589530 655180 589586
rect 654452 577838 654508 577894
rect 654356 566146 654412 566202
rect 654452 554454 654508 554510
rect 654164 542614 654220 542670
rect 654068 530922 654124 530978
rect 654068 519230 654124 519286
rect 654260 484006 654316 484062
rect 654452 472205 654454 472222
rect 654454 472205 654506 472222
rect 654506 472205 654508 472222
rect 654452 472166 654508 472205
rect 654452 460474 654508 460530
rect 654356 448782 654412 448838
rect 654452 436942 654508 436998
rect 654452 425398 654508 425454
rect 653876 413558 653932 413614
rect 655412 683510 655468 683566
rect 655316 636594 655372 636650
rect 655220 495698 655276 495754
rect 654452 401718 654508 401774
rect 654452 390026 654508 390082
rect 654452 378482 654508 378538
rect 654452 366494 654508 366550
rect 654452 343110 654508 343166
rect 654452 331566 654508 331622
rect 655124 319726 655180 319782
rect 656372 507390 656428 507446
rect 655316 354802 655372 354858
rect 654452 284650 654508 284706
rect 647924 210354 647980 210410
rect 646292 166546 646348 166602
rect 647924 166250 647980 166306
rect 647060 165954 647116 166010
rect 655220 307886 655276 307942
rect 655412 296194 655468 296250
rect 673844 942510 673900 942566
rect 672116 718438 672172 718494
rect 673172 755438 673228 755494
rect 673076 752330 673132 752386
rect 675380 957754 675436 957810
rect 675092 953462 675148 953518
rect 675476 955978 675532 956034
rect 675188 953314 675244 953370
rect 673940 939550 673996 939606
rect 674516 945322 674572 945378
rect 674516 944730 674572 944786
rect 674900 943990 674956 944046
rect 674516 942806 674572 942862
rect 674420 941957 674422 941974
rect 674422 941957 674474 941974
rect 674474 941957 674476 941974
rect 674420 941918 674476 941957
rect 674420 941143 674422 941160
rect 674422 941143 674474 941160
rect 674474 941143 674476 941160
rect 674420 941104 674476 941143
rect 676820 936590 676876 936646
rect 679796 928598 679852 928654
rect 679796 928006 679852 928062
rect 675764 876946 675820 877002
rect 675380 876502 675436 876558
rect 675380 875910 675436 875966
rect 675092 875762 675148 875818
rect 675188 875614 675244 875670
rect 675476 873986 675532 874042
rect 675380 873394 675436 873450
rect 675380 869842 675436 869898
rect 675764 864662 675820 864718
rect 675380 862886 675436 862942
rect 675668 787998 675724 788054
rect 675476 787110 675532 787166
rect 675764 786666 675820 786722
rect 675764 784742 675820 784798
rect 675476 780598 675532 780654
rect 674516 777490 674572 777546
rect 675764 779118 675820 779174
rect 675764 777342 675820 777398
rect 675764 775418 675820 775474
rect 675476 773642 675532 773698
rect 674132 773050 674188 773106
rect 674420 767465 674422 767482
rect 674422 767465 674474 767482
rect 674474 767465 674476 767482
rect 674420 767426 674476 767465
rect 674612 766873 674614 766890
rect 674614 766873 674666 766890
rect 674666 766873 674668 766890
rect 674612 766834 674668 766873
rect 674420 765837 674422 765854
rect 674422 765837 674474 765854
rect 674474 765837 674476 765854
rect 674420 765798 674476 765837
rect 673844 765058 673900 765114
rect 673844 764170 673900 764226
rect 674420 763521 674476 763560
rect 674420 763504 674422 763521
rect 674422 763504 674474 763521
rect 674474 763504 674476 763521
rect 673844 762690 673900 762746
rect 673364 753218 673420 753274
rect 673268 751590 673324 751646
rect 679796 750110 679852 750166
rect 679796 749518 679852 749574
rect 675380 743154 675436 743210
rect 673268 674038 673324 674094
rect 673172 661310 673228 661366
rect 673940 716997 673942 717014
rect 673942 716997 673994 717014
rect 673994 716997 673996 717014
rect 673940 716958 673996 716997
rect 673844 674778 673900 674834
rect 673748 673298 673804 673354
rect 673364 662198 673420 662254
rect 673268 629786 673324 629842
rect 673076 616318 673132 616374
rect 673076 530034 673132 530090
rect 673268 582278 673324 582334
rect 674420 722473 674422 722490
rect 674422 722473 674474 722490
rect 674474 722473 674476 722490
rect 674420 722434 674476 722473
rect 674420 720845 674422 720862
rect 674422 720845 674474 720862
rect 674474 720845 674476 720862
rect 674420 720806 674476 720845
rect 674420 710485 674422 710502
rect 674422 710485 674474 710502
rect 674474 710485 674476 710502
rect 674420 710446 674476 710485
rect 674420 707377 674422 707394
rect 674422 707377 674474 707394
rect 674474 707377 674476 707394
rect 674420 707338 674476 707377
rect 674324 668562 674380 668618
rect 674228 667748 674284 667804
rect 673844 664418 673900 664474
rect 673844 663826 673900 663882
rect 674132 630691 674188 630730
rect 674132 630674 674134 630691
rect 674134 630674 674186 630691
rect 674186 630674 674188 630691
rect 673844 629046 673900 629102
rect 673748 628306 673804 628362
rect 675764 742414 675820 742470
rect 675764 741674 675820 741730
rect 675476 740342 675532 740398
rect 675476 739306 675532 739362
rect 675380 738566 675436 738622
rect 674708 727910 674764 727966
rect 674708 721881 674710 721898
rect 674710 721881 674762 721898
rect 674762 721881 674764 721898
rect 674708 721842 674764 721881
rect 674708 720253 674710 720270
rect 674710 720253 674762 720270
rect 674762 720253 674764 720270
rect 674708 720214 674764 720253
rect 674708 719047 674764 719086
rect 674708 719030 674710 719047
rect 674710 719030 674762 719047
rect 674762 719030 674764 719047
rect 674708 711521 674710 711538
rect 674710 711521 674762 711538
rect 674762 711521 674764 711538
rect 674708 711482 674764 711521
rect 674708 708413 674710 708430
rect 674710 708413 674762 708430
rect 674762 708413 674764 708430
rect 674708 708374 674764 708413
rect 674708 706785 674710 706802
rect 674710 706785 674762 706802
rect 674762 706785 674764 706802
rect 674708 706746 674764 706785
rect 679796 705118 679852 705174
rect 679796 704526 679852 704582
rect 675476 697866 675532 697922
rect 675764 697274 675820 697330
rect 675764 697126 675820 697182
rect 675668 694758 675724 694814
rect 675476 694314 675532 694370
rect 675476 693426 675532 693482
rect 675764 691650 675820 691706
rect 674708 677481 674710 677498
rect 674710 677481 674762 677498
rect 674762 677481 674764 677498
rect 674708 677442 674764 677481
rect 674708 676719 674764 676758
rect 674708 676702 674710 676719
rect 674710 676702 674762 676719
rect 674762 676702 674764 676719
rect 675380 689134 675436 689190
rect 674900 687506 674956 687562
rect 674708 675853 674710 675870
rect 674710 675853 674762 675870
rect 674762 675853 674764 675870
rect 674708 675814 674764 675853
rect 674708 672262 674764 672318
rect 674516 671078 674572 671134
rect 674516 632489 674518 632506
rect 674518 632489 674570 632506
rect 674570 632489 674572 632506
rect 674516 632450 674572 632489
rect 674516 631749 674518 631766
rect 674518 631749 674570 631766
rect 674570 631749 674572 631766
rect 674516 631710 674572 631749
rect 674420 625864 674476 625920
rect 679700 659978 679756 660034
rect 679700 659238 679756 659294
rect 674804 653614 674860 653670
rect 675380 652578 675436 652634
rect 675476 652134 675532 652190
rect 675476 651394 675532 651450
rect 675764 649766 675820 649822
rect 675476 648878 675532 648934
rect 675764 645326 675820 645382
rect 675380 640294 675436 640350
rect 675476 638518 675532 638574
rect 675380 628010 675436 628066
rect 674612 623718 674668 623774
rect 674324 622682 674380 622738
rect 675380 620018 675436 620074
rect 674420 617985 674422 618002
rect 674422 617985 674474 618002
rect 674474 617985 674476 618002
rect 674420 617946 674476 617985
rect 675764 638074 675820 638130
rect 675764 630970 675820 631026
rect 675764 630822 675820 630878
rect 675764 630378 675820 630434
rect 679700 614986 679756 615042
rect 679700 614394 679756 614450
rect 673364 575174 673420 575230
rect 675380 607734 675436 607790
rect 675476 607142 675532 607198
rect 675668 606402 675724 606458
rect 675380 604774 675436 604830
rect 675476 600186 675532 600242
rect 674612 586718 674668 586774
rect 673844 586274 673900 586330
rect 674420 585425 674422 585442
rect 674422 585425 674474 585442
rect 674474 585425 674476 585442
rect 674420 585386 674476 585425
rect 673844 584646 673900 584702
rect 673844 583758 673900 583814
rect 674612 583353 674614 583370
rect 674614 583353 674666 583370
rect 674666 583353 674668 583370
rect 674612 583314 674668 583353
rect 674420 574325 674422 574342
rect 674422 574325 674474 574342
rect 674474 574325 674476 574342
rect 674420 574286 674476 574325
rect 673844 573546 673900 573602
rect 674420 572845 674422 572862
rect 674422 572845 674474 572862
rect 674474 572845 674476 572862
rect 674420 572806 674476 572845
rect 674420 571957 674422 571974
rect 674422 571957 674474 571974
rect 674474 571957 674476 571974
rect 674420 571918 674476 571957
rect 673844 571178 673900 571234
rect 675764 593378 675820 593434
rect 679796 570142 679852 570198
rect 679796 569254 679852 569310
rect 674900 568662 674956 568718
rect 673556 526926 673612 526982
rect 673172 526186 673228 526242
rect 673940 541430 673996 541486
rect 674324 542022 674380 542078
rect 674420 541430 674476 541486
rect 674612 541447 674668 541486
rect 674612 541430 674614 541447
rect 674614 541430 674666 541447
rect 674666 541430 674668 541447
rect 674612 540729 674614 540746
rect 674614 540729 674666 540746
rect 674666 540729 674668 540746
rect 674612 540690 674668 540729
rect 674612 539841 674614 539858
rect 674614 539841 674666 539858
rect 674666 539841 674668 539858
rect 674612 539802 674668 539841
rect 674420 497291 674422 497308
rect 674422 497291 674474 497308
rect 674474 497291 674476 497308
rect 674420 497252 674476 497291
rect 674420 496477 674422 496494
rect 674422 496477 674474 496494
rect 674474 496477 674476 496494
rect 674420 496438 674476 496477
rect 674516 491850 674572 491906
rect 674324 489334 674380 489390
rect 675476 562446 675532 562502
rect 675476 562002 675532 562058
rect 675476 561706 675532 561762
rect 675476 558746 675532 558802
rect 675380 558154 675436 558210
rect 675764 557562 675820 557618
rect 675380 554454 675436 554510
rect 676724 538618 676780 538674
rect 676532 537582 676588 537638
rect 676628 536990 676684 537046
rect 674804 531109 674806 531126
rect 674806 531109 674858 531126
rect 674858 531109 674860 531126
rect 674804 531070 674860 531109
rect 674804 529481 674806 529498
rect 674806 529481 674858 529498
rect 674858 529481 674860 529498
rect 674804 529442 674860 529481
rect 674804 528889 674806 528906
rect 674806 528889 674858 528906
rect 674858 528889 674860 528906
rect 674804 528850 674860 528889
rect 674804 528001 674806 528018
rect 674806 528001 674858 528018
rect 674858 528001 674860 528018
rect 674804 527962 674860 528001
rect 674708 497770 674764 497826
rect 674612 488742 674668 488798
rect 676532 493922 676588 493978
rect 674996 490222 675052 490278
rect 674900 485486 674956 485542
rect 674228 484598 674284 484654
rect 673748 482230 673804 482286
rect 679796 524706 679852 524762
rect 679796 524114 679852 524170
rect 676724 495846 676780 495902
rect 676724 494514 676780 494570
rect 676628 493034 676684 493090
rect 676532 412078 676588 412134
rect 676628 411930 676684 411986
rect 674708 409266 674764 409322
rect 674420 409044 674476 409100
rect 674708 408395 674764 408434
rect 674708 408378 674710 408395
rect 674710 408378 674762 408395
rect 674762 408378 674764 408395
rect 679796 480750 679852 480806
rect 679796 480010 679852 480066
rect 676724 407638 676780 407694
rect 673844 406602 673900 406658
rect 674036 404234 674092 404290
rect 673940 401866 673996 401922
rect 675380 402014 675436 402070
rect 675188 399350 675244 399406
rect 674612 398462 674668 398518
rect 674324 397870 674380 397926
rect 674132 397130 674188 397186
rect 674900 396094 674956 396150
rect 674708 393726 674764 393782
rect 675092 395354 675148 395410
rect 674996 394466 675052 394522
rect 679700 392542 679756 392598
rect 679700 392098 679756 392154
rect 675476 378778 675532 378834
rect 675188 374486 675244 374542
rect 675092 374042 675148 374098
rect 675476 373894 675532 373950
rect 675380 371970 675436 372026
rect 674708 364905 674710 364922
rect 674710 364905 674762 364922
rect 674762 364905 674764 364922
rect 674708 364866 674764 364905
rect 674420 363869 674422 363886
rect 674422 363869 674474 363886
rect 674474 363869 674476 363886
rect 674420 363830 674476 363869
rect 674708 363277 674710 363294
rect 674710 363277 674762 363294
rect 674762 363277 674764 363294
rect 674708 363238 674764 363277
rect 673844 362202 673900 362258
rect 673940 359094 673996 359150
rect 677108 358058 677164 358114
rect 674612 357170 674668 357226
rect 674324 352730 674380 352786
rect 674228 351250 674284 351306
rect 674036 349474 674092 349530
rect 674132 348734 674188 348790
rect 675188 356430 675244 356486
rect 675092 353322 675148 353378
rect 674804 350214 674860 350270
rect 676916 355690 676972 355746
rect 675284 354062 675340 354118
rect 676820 351694 676876 351750
rect 677012 354950 677068 355006
rect 676916 345330 676972 345386
rect 679796 347402 679852 347458
rect 679796 346662 679852 346718
rect 677108 345478 677164 345534
rect 677012 345182 677068 345238
rect 675476 335118 675532 335174
rect 675476 333786 675532 333842
rect 675764 333490 675820 333546
rect 675188 329494 675244 329550
rect 675764 328014 675820 328070
rect 675764 326830 675820 326886
rect 674420 319691 674422 319708
rect 674422 319691 674474 319708
rect 674474 319691 674476 319708
rect 674420 319652 674476 319691
rect 674420 318877 674422 318894
rect 674422 318877 674474 318894
rect 674474 318877 674476 318894
rect 674420 318838 674476 318877
rect 674708 318285 674710 318302
rect 674710 318285 674762 318302
rect 674762 318285 674764 318302
rect 674708 318246 674764 318285
rect 674036 314102 674092 314158
rect 673940 311586 673996 311642
rect 675092 312178 675148 312234
rect 674900 309070 674956 309126
rect 674228 308478 674284 308534
rect 674132 303742 674188 303798
rect 674612 307442 674668 307498
rect 674324 305370 674380 305426
rect 674420 304556 674476 304612
rect 676916 310698 676972 310754
rect 676820 305962 676876 306018
rect 677108 309958 677164 310014
rect 677012 306702 677068 306758
rect 677012 299450 677068 299506
rect 679796 302410 679852 302466
rect 679796 301670 679852 301726
rect 677108 299302 677164 299358
rect 675476 289682 675532 289738
rect 675380 289534 675436 289590
rect 675188 284946 675244 285002
rect 675764 284798 675820 284854
rect 675380 283614 675436 283670
rect 675764 281838 675820 281894
rect 674708 274921 674710 274938
rect 674710 274921 674762 274938
rect 674762 274921 674764 274938
rect 674708 274882 674764 274921
rect 674708 274033 674710 274050
rect 674710 274033 674762 274050
rect 674762 274033 674764 274050
rect 674708 273994 674764 274033
rect 674708 273293 674710 273310
rect 674710 273293 674762 273310
rect 674762 273293 674764 273310
rect 674708 273254 674764 273293
rect 674132 269110 674188 269166
rect 673940 266594 673996 266650
rect 674036 263486 674092 263542
rect 674516 267186 674572 267242
rect 674324 262746 674380 262802
rect 674228 258750 674284 258806
rect 673364 244690 673420 244746
rect 673844 244542 673900 244598
rect 673844 242174 673900 242230
rect 673364 242026 673420 242082
rect 678164 264966 678220 265022
rect 674612 264078 674668 264134
rect 676916 261710 676972 261766
rect 676820 260970 676876 261026
rect 675284 260082 675340 260138
rect 675188 259342 675244 259398
rect 674804 245874 674860 245930
rect 674900 245134 674956 245190
rect 674900 244838 674956 244894
rect 674900 241878 674956 241934
rect 679796 257418 679852 257474
rect 679796 256826 679852 256882
rect 678164 253422 678220 253478
rect 675476 245134 675532 245190
rect 675476 243506 675532 243562
rect 674804 238918 674860 238974
rect 675476 238622 675532 238678
rect 675764 236846 675820 236902
rect 674420 229485 674422 229502
rect 674422 229485 674474 229502
rect 674474 229485 674476 229502
rect 674420 229446 674476 229485
rect 674708 228893 674710 228910
rect 674710 228893 674762 228910
rect 674762 228893 674764 228910
rect 674708 228854 674764 228893
rect 674420 227857 674422 227874
rect 674422 227857 674474 227874
rect 674474 227857 674476 227874
rect 674420 227818 674476 227857
rect 674708 225785 674710 225802
rect 674710 225785 674762 225802
rect 674762 225785 674764 225802
rect 674708 225746 674764 225785
rect 673844 224727 673900 224766
rect 673844 224710 673846 224727
rect 673846 224710 673898 224727
rect 673898 224710 673900 224727
rect 673940 223822 673996 223878
rect 674420 222194 674476 222250
rect 674036 217458 674092 217514
rect 674996 221158 675052 221214
rect 674900 214646 674956 214702
rect 674804 214202 674860 214258
rect 674708 213314 674764 213370
rect 677012 220566 677068 220622
rect 675188 218938 675244 218994
rect 675092 217754 675148 217810
rect 676916 216422 676972 216478
rect 676820 215830 676876 215886
rect 677108 219678 677164 219734
rect 677012 207690 677068 207746
rect 679796 212130 679852 212186
rect 679796 211390 679852 211446
rect 680084 210206 680140 210262
rect 679988 210058 680044 210114
rect 677108 207542 677164 207598
rect 676916 207394 676972 207450
rect 675380 199254 675436 199310
rect 675476 198662 675532 198718
rect 675764 198366 675820 198422
rect 675764 195258 675820 195314
rect 675380 193482 675436 193538
rect 675764 191558 675820 191614
rect 674420 184454 674476 184510
rect 674708 183901 674710 183918
rect 674710 183901 674762 183918
rect 674762 183901 674764 183918
rect 674708 183862 674764 183901
rect 674420 182865 674422 182882
rect 674422 182865 674474 182882
rect 674474 182865 674476 182882
rect 674420 182826 674476 182865
rect 679700 179866 679756 179922
rect 674900 177054 674956 177110
rect 674804 173058 674860 173114
rect 674516 172318 674572 172374
rect 674228 169358 674284 169414
rect 674132 168470 674188 168526
rect 674708 167286 674764 167342
rect 674612 166546 674668 166602
rect 674708 165658 674764 165714
rect 677012 176166 677068 176222
rect 676916 175574 676972 175630
rect 674996 173946 675052 174002
rect 676820 170838 676876 170894
rect 675092 169950 675148 170006
rect 675764 166398 675820 166454
rect 675764 165510 675820 165566
rect 676916 162846 676972 162902
rect 677204 174686 677260 174742
rect 677108 171430 677164 171486
rect 679796 179422 679852 179478
rect 679700 166546 679756 166602
rect 679796 166398 679852 166454
rect 677204 164030 677260 164086
rect 677012 161366 677068 161422
rect 675380 159294 675436 159350
rect 675764 157666 675820 157722
rect 675380 154558 675436 154614
rect 675380 154262 675436 154318
rect 675764 153374 675820 153430
rect 675476 148490 675532 148546
rect 675188 148342 675244 148398
rect 675764 146566 675820 146622
rect 674708 139018 674764 139074
rect 674420 138443 674476 138482
rect 674420 138426 674422 138443
rect 674422 138426 674474 138443
rect 674474 138426 674476 138443
rect 674612 137242 674668 137298
rect 674708 135614 674764 135670
rect 673556 134874 673612 134930
rect 675476 131766 675532 131822
rect 675188 131026 675244 131082
rect 674804 128658 674860 128714
rect 674516 124810 674572 124866
rect 674324 124218 674380 124274
rect 674132 123330 674188 123386
rect 647732 121406 647788 121462
rect 647828 121110 647884 121166
rect 647924 120814 647980 120870
rect 646484 120370 646540 120426
rect 674420 121036 674476 121092
rect 674708 122294 674764 122350
rect 674612 121258 674668 121314
rect 675092 127918 675148 127974
rect 674900 127030 674956 127086
rect 677012 130286 677068 130342
rect 676916 126290 676972 126346
rect 676820 125550 676876 125606
rect 677108 129546 677164 129602
rect 677012 120370 677068 120426
rect 677108 118002 677164 118058
rect 675380 114154 675436 114210
rect 675380 110010 675436 110066
rect 675092 109270 675148 109326
rect 675764 108086 675820 108142
rect 675092 106458 675148 106514
rect 668180 105126 668236 105182
rect 665204 104551 665260 104590
rect 665204 104534 665206 104551
rect 665206 104534 665258 104551
rect 665258 104534 665260 104551
rect 647924 104238 647980 104294
rect 675380 103202 675436 103258
rect 675764 101426 675820 101482
rect 646196 85738 646252 85794
rect 645908 84110 645964 84166
rect 646484 76897 646486 76914
rect 646486 76897 646538 76914
rect 646538 76897 646540 76914
rect 646484 76858 646540 76897
rect 646484 75970 646540 76026
rect 646484 75417 646486 75434
rect 646486 75417 646538 75434
rect 646538 75417 646540 75434
rect 646484 75378 646540 75417
rect 646100 75230 646156 75286
rect 646100 72862 646156 72918
rect 646868 88106 646924 88162
rect 646868 84998 646924 85054
rect 647252 83814 647308 83870
rect 647444 87366 647500 87422
rect 647348 80854 647404 80910
rect 647636 88994 647692 89050
rect 647540 82186 647596 82242
rect 647924 87662 647980 87718
rect 647924 86495 647980 86534
rect 647924 86478 647926 86495
rect 647926 86478 647978 86495
rect 647978 86478 647980 86495
rect 647828 86182 647884 86238
rect 647732 85442 647788 85498
rect 650996 86922 651052 86978
rect 650900 85294 650956 85350
rect 650996 84258 651052 84314
rect 647924 83409 647926 83426
rect 647926 83409 647978 83426
rect 647978 83409 647980 83426
rect 647924 83370 647980 83409
rect 650900 82630 650956 82686
rect 647924 82482 647980 82538
rect 647924 81315 647980 81354
rect 647924 81298 647926 81315
rect 647926 81298 647978 81315
rect 647978 81298 647980 81315
rect 647828 80410 647884 80466
rect 647732 78930 647788 78986
rect 647924 80153 647926 80170
rect 647926 80153 647978 80170
rect 647978 80153 647980 80170
rect 647924 80114 647980 80153
rect 647924 79226 647980 79282
rect 647924 77637 647926 77654
rect 647926 77637 647978 77654
rect 647978 77637 647980 77654
rect 647924 77598 647980 77637
rect 647924 77006 647980 77062
rect 651188 86182 651244 86238
rect 651092 83370 651148 83426
rect 663380 85590 663436 85646
rect 663284 85146 663340 85202
rect 663476 84702 663532 84758
rect 662900 81150 662956 81206
rect 647252 74342 647308 74398
rect 646868 73750 646924 73806
rect 646676 72566 646732 72622
rect 663380 82778 663436 82834
rect 663284 82038 663340 82094
rect 646484 72122 646540 72178
rect 640724 40598 640780 40654
rect 454964 40302 455020 40358
rect 136532 40154 136588 40210
<< metal3 >>
rect 497826 1019912 499518 1019972
rect 115695 1005616 115761 1005619
rect 115488 1005614 115761 1005616
rect 115488 1005558 115700 1005614
rect 115756 1005558 115761 1005614
rect 115488 1005556 115761 1005558
rect 115695 1005553 115761 1005556
rect 102159 1005468 102225 1005471
rect 312783 1005468 312849 1005471
rect 313839 1005468 313905 1005471
rect 321039 1005468 321105 1005471
rect 102159 1005466 102720 1005468
rect 102159 1005410 102164 1005466
rect 102220 1005410 102720 1005466
rect 102159 1005408 102720 1005410
rect 312783 1005466 313248 1005468
rect 312783 1005410 312788 1005466
rect 312844 1005410 313248 1005466
rect 312783 1005408 313248 1005410
rect 313839 1005466 314016 1005468
rect 313839 1005410 313844 1005466
rect 313900 1005410 314016 1005466
rect 313839 1005408 314016 1005410
rect 320448 1005466 321105 1005468
rect 320448 1005410 321044 1005466
rect 321100 1005410 321105 1005466
rect 320448 1005408 321105 1005410
rect 102159 1005405 102225 1005408
rect 312783 1005405 312849 1005408
rect 313839 1005405 313905 1005408
rect 321039 1005405 321105 1005408
rect 321423 1005468 321489 1005471
rect 325455 1005468 325521 1005471
rect 365103 1005468 365169 1005471
rect 430863 1005468 430929 1005471
rect 433167 1005468 433233 1005471
rect 321423 1005466 325521 1005468
rect 321423 1005410 321428 1005466
rect 321484 1005410 325460 1005466
rect 325516 1005410 325521 1005466
rect 321423 1005408 325521 1005410
rect 364512 1005466 365169 1005468
rect 364512 1005410 365108 1005466
rect 365164 1005410 365169 1005466
rect 364512 1005408 365169 1005410
rect 430368 1005466 430929 1005468
rect 430368 1005410 430868 1005466
rect 430924 1005410 430929 1005466
rect 430368 1005408 430929 1005410
rect 432672 1005466 433233 1005468
rect 432672 1005410 433172 1005466
rect 433228 1005410 433233 1005466
rect 432672 1005408 433233 1005410
rect 321423 1005405 321489 1005408
rect 325455 1005405 325521 1005408
rect 365103 1005405 365169 1005408
rect 430863 1005405 430929 1005408
rect 433167 1005405 433233 1005408
rect 101487 1005320 101553 1005323
rect 114159 1005320 114225 1005323
rect 308751 1005320 308817 1005323
rect 309615 1005320 309681 1005323
rect 318639 1005320 318705 1005323
rect 358671 1005320 358737 1005323
rect 359919 1005320 359985 1005323
rect 425295 1005320 425361 1005323
rect 431535 1005320 431601 1005323
rect 101487 1005318 102048 1005320
rect 101487 1005262 101492 1005318
rect 101548 1005262 102048 1005318
rect 101487 1005260 102048 1005262
rect 114159 1005318 114720 1005320
rect 114159 1005262 114164 1005318
rect 114220 1005262 114720 1005318
rect 114159 1005260 114720 1005262
rect 308751 1005318 309312 1005320
rect 308751 1005262 308756 1005318
rect 308812 1005262 309312 1005318
rect 308751 1005260 309312 1005262
rect 309615 1005318 310176 1005320
rect 309615 1005262 309620 1005318
rect 309676 1005262 310176 1005318
rect 309615 1005260 310176 1005262
rect 318048 1005318 318705 1005320
rect 318048 1005262 318644 1005318
rect 318700 1005262 318705 1005318
rect 318048 1005260 318705 1005262
rect 358176 1005318 358737 1005320
rect 358176 1005262 358676 1005318
rect 358732 1005262 358737 1005318
rect 358176 1005260 358737 1005262
rect 359712 1005318 359985 1005320
rect 359712 1005262 359924 1005318
rect 359980 1005262 359985 1005318
rect 359712 1005260 359985 1005262
rect 424800 1005318 425361 1005320
rect 424800 1005262 425300 1005318
rect 425356 1005262 425361 1005318
rect 424800 1005260 425361 1005262
rect 431040 1005318 431601 1005320
rect 431040 1005262 431540 1005318
rect 431596 1005262 431601 1005318
rect 431040 1005260 431601 1005262
rect 101487 1005257 101553 1005260
rect 114159 1005257 114225 1005260
rect 308751 1005257 308817 1005260
rect 309615 1005257 309681 1005260
rect 318639 1005257 318705 1005260
rect 358671 1005257 358737 1005260
rect 359919 1005257 359985 1005260
rect 425295 1005257 425361 1005260
rect 431535 1005257 431601 1005260
rect 105423 1005172 105489 1005175
rect 209007 1005172 209073 1005175
rect 310287 1005172 310353 1005175
rect 357039 1005172 357105 1005175
rect 364239 1005172 364305 1005175
rect 427599 1005172 427665 1005175
rect 435567 1005172 435633 1005175
rect 105423 1005170 105984 1005172
rect 105423 1005114 105428 1005170
rect 105484 1005114 105984 1005170
rect 105423 1005112 105984 1005114
rect 209007 1005170 209568 1005172
rect 209007 1005114 209012 1005170
rect 209068 1005114 209568 1005170
rect 209007 1005112 209568 1005114
rect 310287 1005170 310944 1005172
rect 310287 1005114 310292 1005170
rect 310348 1005114 310944 1005170
rect 310287 1005112 310944 1005114
rect 356640 1005170 357105 1005172
rect 356640 1005114 357044 1005170
rect 357100 1005114 357105 1005170
rect 356640 1005112 357105 1005114
rect 363648 1005170 364305 1005172
rect 363648 1005114 364244 1005170
rect 364300 1005114 364305 1005170
rect 363648 1005112 364305 1005114
rect 427104 1005170 427665 1005172
rect 427104 1005114 427604 1005170
rect 427660 1005114 427665 1005170
rect 427104 1005112 427665 1005114
rect 435168 1005170 435633 1005172
rect 435168 1005114 435572 1005170
rect 435628 1005114 435633 1005170
rect 497826 1005172 497886 1019912
rect 499458 1019824 499518 1019912
rect 499296 1019764 499518 1019824
rect 554511 1005468 554577 1005471
rect 554016 1005466 554577 1005468
rect 554016 1005410 554516 1005466
rect 554572 1005410 554577 1005466
rect 554016 1005408 554577 1005410
rect 554511 1005405 554577 1005408
rect 500655 1005320 500721 1005323
rect 556911 1005320 556977 1005323
rect 500160 1005318 500721 1005320
rect 500160 1005262 500660 1005318
rect 500716 1005262 500721 1005318
rect 500160 1005260 500721 1005262
rect 556320 1005318 556977 1005320
rect 556320 1005262 556916 1005318
rect 556972 1005262 556977 1005318
rect 556320 1005260 556977 1005262
rect 500655 1005257 500721 1005260
rect 556911 1005257 556977 1005260
rect 498159 1005172 498225 1005175
rect 501135 1005172 501201 1005175
rect 553743 1005172 553809 1005175
rect 562479 1005172 562545 1005175
rect 497826 1005170 498225 1005172
rect 497826 1005142 498164 1005170
rect 435168 1005112 435633 1005114
rect 497856 1005114 498164 1005142
rect 498220 1005114 498225 1005170
rect 497856 1005112 498225 1005114
rect 501024 1005170 501201 1005172
rect 501024 1005114 501140 1005170
rect 501196 1005114 501201 1005170
rect 501024 1005112 501201 1005114
rect 553248 1005170 553809 1005172
rect 553248 1005114 553748 1005170
rect 553804 1005114 553809 1005170
rect 553248 1005112 553809 1005114
rect 561888 1005170 562545 1005172
rect 561888 1005114 562484 1005170
rect 562540 1005114 562545 1005170
rect 561888 1005112 562545 1005114
rect 105423 1005109 105489 1005112
rect 209007 1005109 209073 1005112
rect 310287 1005109 310353 1005112
rect 357039 1005109 357105 1005112
rect 364239 1005109 364305 1005112
rect 427599 1005109 427665 1005112
rect 435567 1005109 435633 1005112
rect 498159 1005109 498225 1005112
rect 501135 1005109 501201 1005112
rect 553743 1005109 553809 1005112
rect 562479 1005109 562545 1005112
rect 428079 1003988 428145 1003991
rect 427872 1003986 428145 1003988
rect 427872 1003930 428084 1003986
rect 428140 1003930 428145 1003986
rect 427872 1003928 428145 1003930
rect 428079 1003925 428145 1003928
rect 357615 1003840 357681 1003843
rect 359055 1003840 359121 1003843
rect 423375 1003840 423441 1003843
rect 426447 1003840 426513 1003843
rect 554895 1003840 554961 1003843
rect 357408 1003838 357681 1003840
rect 357408 1003782 357620 1003838
rect 357676 1003782 357681 1003838
rect 357408 1003780 357681 1003782
rect 358944 1003838 359121 1003840
rect 358944 1003782 359060 1003838
rect 359116 1003782 359121 1003838
rect 358944 1003780 359121 1003782
rect 423168 1003838 423441 1003840
rect 423168 1003782 423380 1003838
rect 423436 1003782 423441 1003838
rect 423168 1003780 423441 1003782
rect 426336 1003838 426513 1003840
rect 426336 1003782 426452 1003838
rect 426508 1003782 426513 1003838
rect 426336 1003780 426513 1003782
rect 554688 1003838 554961 1003840
rect 554688 1003782 554900 1003838
rect 554956 1003782 554961 1003838
rect 554688 1003780 554961 1003782
rect 357615 1003777 357681 1003780
rect 359055 1003777 359121 1003780
rect 423375 1003777 423441 1003780
rect 426447 1003777 426513 1003780
rect 554895 1003777 554961 1003780
rect 108879 1003692 108945 1003695
rect 355983 1003692 356049 1003695
rect 425775 1003692 425841 1003695
rect 555663 1003692 555729 1003695
rect 108879 1003690 109152 1003692
rect 108879 1003634 108884 1003690
rect 108940 1003634 109152 1003690
rect 108879 1003632 109152 1003634
rect 355776 1003690 356049 1003692
rect 355776 1003634 355988 1003690
rect 356044 1003634 356049 1003690
rect 355776 1003632 356049 1003634
rect 425568 1003690 425841 1003692
rect 425568 1003634 425780 1003690
rect 425836 1003634 425841 1003690
rect 425568 1003632 425841 1003634
rect 555552 1003690 555729 1003692
rect 555552 1003634 555668 1003690
rect 555724 1003634 555729 1003690
rect 555552 1003632 555729 1003634
rect 108879 1003629 108945 1003632
rect 355983 1003629 356049 1003632
rect 425775 1003629 425841 1003632
rect 555663 1003629 555729 1003632
rect 308079 1002656 308145 1002659
rect 308079 1002654 308448 1002656
rect 308079 1002598 308084 1002654
rect 308140 1002598 308448 1002654
rect 308079 1002596 308448 1002598
rect 308079 1002593 308145 1002596
rect 102831 1002508 102897 1002511
rect 151215 1002508 151281 1002511
rect 157935 1002508 158001 1002511
rect 503439 1002508 503505 1002511
rect 559119 1002508 559185 1002511
rect 560559 1002508 560625 1002511
rect 102831 1002506 103488 1002508
rect 102831 1002450 102836 1002506
rect 102892 1002450 103488 1002506
rect 102831 1002448 103488 1002450
rect 151215 1002506 151776 1002508
rect 151215 1002450 151220 1002506
rect 151276 1002450 151776 1002506
rect 151215 1002448 151776 1002450
rect 157935 1002506 158208 1002508
rect 157935 1002450 157940 1002506
rect 157996 1002450 158208 1002506
rect 157935 1002448 158208 1002450
rect 503328 1002506 503505 1002508
rect 503328 1002450 503444 1002506
rect 503500 1002450 503505 1002506
rect 503328 1002448 503505 1002450
rect 558816 1002506 559185 1002508
rect 558816 1002450 559124 1002506
rect 559180 1002450 559185 1002506
rect 558816 1002448 559185 1002450
rect 560256 1002506 560625 1002508
rect 560256 1002450 560564 1002506
rect 560620 1002450 560625 1002506
rect 560256 1002448 560625 1002450
rect 102831 1002445 102897 1002448
rect 151215 1002445 151281 1002448
rect 157935 1002445 158001 1002448
rect 503439 1002445 503505 1002448
rect 559119 1002445 559185 1002448
rect 560559 1002445 560625 1002448
rect 100527 1002360 100593 1002363
rect 103791 1002360 103857 1002363
rect 104463 1002360 104529 1002363
rect 150351 1002360 150417 1002363
rect 505071 1002360 505137 1002363
rect 560079 1002360 560145 1002363
rect 561519 1002360 561585 1002363
rect 564783 1002360 564849 1002363
rect 100527 1002358 101184 1002360
rect 100527 1002302 100532 1002358
rect 100588 1002302 101184 1002358
rect 100527 1002300 101184 1002302
rect 103791 1002358 104352 1002360
rect 103791 1002302 103796 1002358
rect 103852 1002302 104352 1002358
rect 103791 1002300 104352 1002302
rect 104463 1002358 105120 1002360
rect 104463 1002302 104468 1002358
rect 104524 1002302 105120 1002358
rect 104463 1002300 105120 1002302
rect 150351 1002358 151008 1002360
rect 150351 1002302 150356 1002358
rect 150412 1002302 151008 1002358
rect 150351 1002300 151008 1002302
rect 504960 1002358 505137 1002360
rect 504960 1002302 505076 1002358
rect 505132 1002302 505137 1002358
rect 504960 1002300 505137 1002302
rect 559488 1002358 560145 1002360
rect 559488 1002302 560084 1002358
rect 560140 1002302 560145 1002358
rect 559488 1002300 560145 1002302
rect 561120 1002358 561585 1002360
rect 561120 1002302 561524 1002358
rect 561580 1002302 561585 1002358
rect 561120 1002300 561585 1002302
rect 564192 1002358 564849 1002360
rect 564192 1002302 564788 1002358
rect 564844 1002302 564849 1002358
rect 564192 1002300 564849 1002302
rect 100527 1002297 100593 1002300
rect 103791 1002297 103857 1002300
rect 104463 1002297 104529 1002300
rect 150351 1002297 150417 1002300
rect 505071 1002297 505137 1002300
rect 560079 1002297 560145 1002300
rect 561519 1002297 561585 1002300
rect 564783 1002297 564849 1002300
rect 434031 1001176 434097 1001179
rect 433536 1001174 434097 1001176
rect 433536 1001118 434036 1001174
rect 434092 1001118 434097 1001174
rect 433536 1001116 434097 1001118
rect 434031 1001113 434097 1001116
rect 208335 1001028 208401 1001031
rect 432495 1001028 432561 1001031
rect 208335 1001026 208800 1001028
rect 208335 1000970 208340 1001026
rect 208396 1000970 208800 1001026
rect 208335 1000968 208800 1000970
rect 431904 1001026 432561 1001028
rect 431904 1000970 432500 1001026
rect 432556 1000970 432561 1001026
rect 431904 1000968 432561 1000970
rect 208335 1000965 208401 1000968
rect 432495 1000965 432561 1000968
rect 160239 1000880 160305 1000883
rect 211695 1000880 211761 1000883
rect 360687 1000880 360753 1000883
rect 361551 1000880 361617 1000883
rect 424143 1000880 424209 1000883
rect 428943 1000880 429009 1000883
rect 160239 1000878 160512 1000880
rect 160239 1000822 160244 1000878
rect 160300 1000822 160512 1000878
rect 160239 1000820 160512 1000822
rect 211695 1000878 211872 1000880
rect 211695 1000822 211700 1000878
rect 211756 1000822 211872 1000878
rect 211695 1000820 211872 1000822
rect 360480 1000878 360753 1000880
rect 360480 1000822 360692 1000878
rect 360748 1000822 360753 1000878
rect 360480 1000820 360753 1000822
rect 361344 1000878 361617 1000880
rect 361344 1000822 361556 1000878
rect 361612 1000822 361617 1000878
rect 361344 1000820 361617 1000822
rect 424032 1000878 424209 1000880
rect 424032 1000822 424148 1000878
rect 424204 1000822 424209 1000878
rect 424032 1000820 424209 1000822
rect 428736 1000878 429009 1000880
rect 428736 1000822 428948 1000878
rect 429004 1000822 429009 1000878
rect 428736 1000820 429009 1000822
rect 160239 1000817 160305 1000820
rect 211695 1000817 211761 1000820
rect 360687 1000817 360753 1000820
rect 361551 1000817 361617 1000820
rect 424143 1000817 424209 1000820
rect 428943 1000817 429009 1000820
rect 509391 1000732 509457 1000735
rect 508896 1000730 509457 1000732
rect 508896 1000674 509396 1000730
rect 509452 1000674 509457 1000730
rect 508896 1000672 509457 1000674
rect 509391 1000669 509457 1000672
rect 516687 1000288 516753 1000291
rect 523791 1000288 523857 1000291
rect 516687 1000286 523857 1000288
rect 516687 1000230 516692 1000286
rect 516748 1000230 523796 1000286
rect 523852 1000230 523857 1000286
rect 516687 1000228 523857 1000230
rect 516687 1000225 516753 1000228
rect 523791 1000225 523857 1000228
rect 503055 999992 503121 999995
rect 502560 999990 503121 999992
rect 502560 999934 503060 999990
rect 503116 999934 503121 999990
rect 502560 999932 503121 999934
rect 503055 999929 503121 999932
rect 509871 999844 509937 999847
rect 509664 999842 509937 999844
rect 509664 999786 509876 999842
rect 509932 999786 509937 999842
rect 509664 999784 509937 999786
rect 509871 999781 509937 999784
rect 516879 999844 516945 999847
rect 523503 999844 523569 999847
rect 516879 999842 523569 999844
rect 516879 999786 516884 999842
rect 516940 999786 523508 999842
rect 523564 999786 523569 999842
rect 516879 999784 523569 999786
rect 516879 999781 516945 999784
rect 523503 999781 523569 999784
rect 506223 999696 506289 999699
rect 507759 999696 507825 999699
rect 505728 999694 506289 999696
rect 505728 999638 506228 999694
rect 506284 999638 506289 999694
rect 505728 999636 506289 999638
rect 507360 999694 507825 999696
rect 507360 999638 507764 999694
rect 507820 999638 507825 999694
rect 507360 999636 507825 999638
rect 506223 999633 506289 999636
rect 507759 999633 507825 999636
rect 516783 999696 516849 999699
rect 523887 999696 523953 999699
rect 516783 999694 523953 999696
rect 516783 999638 516788 999694
rect 516844 999638 523892 999694
rect 523948 999638 523953 999694
rect 516783 999636 523953 999638
rect 516783 999633 516849 999636
rect 523887 999633 523953 999636
rect 256431 999548 256497 999551
rect 314703 999548 314769 999551
rect 315471 999548 315537 999551
rect 502383 999548 502449 999551
rect 508623 999548 508689 999551
rect 256431 999546 256896 999548
rect 256431 999490 256436 999546
rect 256492 999490 256896 999546
rect 256431 999488 256896 999490
rect 314703 999546 314880 999548
rect 314703 999490 314708 999546
rect 314764 999490 314880 999546
rect 314703 999488 314880 999490
rect 315471 999546 315744 999548
rect 315471 999490 315476 999546
rect 315532 999490 315744 999546
rect 315471 999488 315744 999490
rect 501792 999546 502449 999548
rect 501792 999490 502388 999546
rect 502444 999490 502449 999546
rect 501792 999488 502449 999490
rect 508032 999546 508689 999548
rect 508032 999490 508628 999546
rect 508684 999490 508689 999546
rect 508032 999488 508689 999490
rect 256431 999485 256497 999488
rect 314703 999485 314769 999488
rect 315471 999485 315537 999488
rect 502383 999485 502449 999488
rect 508623 999485 508689 999488
rect 516783 999548 516849 999551
rect 523695 999548 523761 999551
rect 516783 999546 523761 999548
rect 516783 999490 516788 999546
rect 516844 999490 523700 999546
rect 523756 999490 523761 999546
rect 516783 999488 523761 999490
rect 516783 999485 516849 999488
rect 523695 999485 523761 999488
rect 156879 999400 156945 999403
rect 259503 999400 259569 999403
rect 311439 999400 311505 999403
rect 488847 999400 488913 999403
rect 497583 999400 497649 999403
rect 156879 999398 157344 999400
rect 156879 999342 156884 999398
rect 156940 999342 157344 999398
rect 156879 999340 157344 999342
rect 259503 999398 260160 999400
rect 259503 999342 259508 999398
rect 259564 999342 260160 999398
rect 259503 999340 260160 999342
rect 311439 999398 311712 999400
rect 311439 999342 311444 999398
rect 311500 999342 311712 999398
rect 311439 999340 311712 999342
rect 488847 999398 497649 999400
rect 488847 999342 488852 999398
rect 488908 999342 497588 999398
rect 497644 999342 497649 999398
rect 488847 999340 497649 999342
rect 156879 999337 156945 999340
rect 259503 999337 259569 999340
rect 311439 999337 311505 999340
rect 488847 999337 488913 999340
rect 497583 999337 497649 999340
rect 516687 999400 516753 999403
rect 524079 999400 524145 999403
rect 552975 999400 553041 999403
rect 516687 999398 524145 999400
rect 516687 999342 516692 999398
rect 516748 999342 524084 999398
rect 524140 999342 524145 999398
rect 516687 999340 524145 999342
rect 552384 999398 553041 999400
rect 552384 999342 552980 999398
rect 553036 999342 553041 999398
rect 552384 999340 553041 999342
rect 516687 999337 516753 999340
rect 524079 999337 524145 999340
rect 552975 999337 553041 999340
rect 367887 997920 367953 997923
rect 557295 997920 557361 997923
rect 367776 997918 367953 997920
rect 367776 997862 367892 997918
rect 367948 997862 367953 997918
rect 367776 997860 367953 997862
rect 557088 997918 557361 997920
rect 557088 997862 557300 997918
rect 557356 997862 557361 997918
rect 557088 997860 557361 997862
rect 367887 997857 367953 997860
rect 557295 997857 557361 997860
rect 369039 997772 369105 997775
rect 369039 997770 369216 997772
rect 369039 997714 369044 997770
rect 369100 997714 369216 997770
rect 369039 997712 369216 997714
rect 369039 997709 369105 997712
rect 204207 996588 204273 996591
rect 263055 996588 263121 996591
rect 204207 996586 204768 996588
rect 204207 996530 204212 996586
rect 204268 996530 204768 996586
rect 204207 996528 204768 996530
rect 263055 996586 263328 996588
rect 263055 996530 263060 996586
rect 263116 996530 263328 996586
rect 263055 996528 263328 996530
rect 204207 996525 204273 996528
rect 263055 996525 263121 996528
rect 573039 996440 573105 996443
rect 604815 996440 604881 996443
rect 573039 996438 604881 996440
rect 573039 996382 573044 996438
rect 573100 996382 604820 996438
rect 604876 996382 604881 996438
rect 573039 996380 604881 996382
rect 573039 996377 573105 996380
rect 604815 996377 604881 996380
rect 436335 996292 436401 996295
rect 436335 996290 436608 996292
rect 436335 996234 436340 996290
rect 436396 996234 436608 996290
rect 436335 996232 436608 996234
rect 436335 996229 436401 996232
rect 162255 996144 162321 996147
rect 163119 996144 163185 996147
rect 162144 996142 162321 996144
rect 162144 996086 162260 996142
rect 162316 996086 162321 996142
rect 162144 996084 162321 996086
rect 162912 996142 163185 996144
rect 162912 996086 163124 996142
rect 163180 996086 163185 996142
rect 162912 996084 163185 996086
rect 162255 996081 162321 996084
rect 163119 996081 163185 996084
rect 164079 996144 164145 996147
rect 213327 996144 213393 996147
rect 214095 996144 214161 996147
rect 215631 996144 215697 996147
rect 265935 996144 266001 996147
rect 164079 996142 164448 996144
rect 164079 996086 164084 996142
rect 164140 996086 164448 996142
rect 164079 996084 164448 996086
rect 213327 996142 213504 996144
rect 213327 996086 213332 996142
rect 213388 996086 213504 996142
rect 213327 996084 213504 996086
rect 214095 996142 214368 996144
rect 214095 996086 214100 996142
rect 214156 996086 214368 996142
rect 214095 996084 214368 996086
rect 215040 996142 215697 996144
rect 215040 996086 215636 996142
rect 215692 996086 215697 996142
rect 215040 996084 215697 996086
rect 265728 996142 266001 996144
rect 265728 996086 265940 996142
rect 265996 996086 266001 996142
rect 265728 996084 266001 996086
rect 164079 996081 164145 996084
rect 213327 996081 213393 996084
rect 214095 996081 214161 996084
rect 215631 996081 215697 996084
rect 265935 996081 266001 996084
rect 266991 996144 267057 996147
rect 317103 996144 317169 996147
rect 318639 996144 318705 996147
rect 399855 996144 399921 996147
rect 436431 996144 436497 996147
rect 266991 996142 267264 996144
rect 266991 996086 266996 996142
rect 267052 996086 267264 996142
rect 266991 996084 267264 996086
rect 317103 996142 317280 996144
rect 317103 996086 317108 996142
rect 317164 996086 317280 996142
rect 317103 996084 317280 996086
rect 318639 996142 318816 996144
rect 318639 996086 318644 996142
rect 318700 996086 318816 996142
rect 318639 996084 318816 996086
rect 399855 996142 418878 996144
rect 399855 996086 399860 996142
rect 399916 996086 418878 996142
rect 399855 996084 418878 996086
rect 435840 996142 436497 996144
rect 435840 996086 436436 996142
rect 436492 996086 436497 996142
rect 435840 996084 436497 996086
rect 266991 996081 267057 996084
rect 317103 996081 317169 996084
rect 318639 996081 318705 996084
rect 399855 996081 399921 996084
rect 106959 995996 107025 995999
rect 113295 995996 113361 995999
rect 144015 995996 144081 995999
rect 106959 995994 107424 995996
rect 106959 995938 106964 995994
rect 107020 995938 107424 995994
rect 106959 995936 107424 995938
rect 113295 995994 113856 995996
rect 113295 995938 113300 995994
rect 113356 995938 113856 995994
rect 113295 995936 113856 995938
rect 136770 995994 144081 995996
rect 136770 995938 144020 995994
rect 144076 995938 144081 995994
rect 136770 995936 144081 995938
rect 106959 995933 107025 995936
rect 113295 995933 113361 995936
rect 136770 995851 136830 995936
rect 144015 995933 144081 995936
rect 145263 995996 145329 995999
rect 149103 995996 149169 995999
rect 145263 995994 149169 995996
rect 145263 995938 145268 995994
rect 145324 995938 149108 995994
rect 149164 995938 149169 995994
rect 145263 995936 149169 995938
rect 145263 995933 145329 995936
rect 149103 995933 149169 995936
rect 149487 995996 149553 995999
rect 151983 995996 152049 995999
rect 152847 995996 152913 995999
rect 155343 995996 155409 995999
rect 164175 995996 164241 995999
rect 198639 995996 198705 995999
rect 203439 995996 203505 995999
rect 205647 995996 205713 995999
rect 206511 995996 206577 995999
rect 215439 995996 215505 995999
rect 217071 995996 217137 995999
rect 221775 995996 221841 995999
rect 246927 995996 246993 995999
rect 149487 995994 150144 995996
rect 149487 995938 149492 995994
rect 149548 995938 150144 995994
rect 149487 995936 150144 995938
rect 151983 995994 152544 995996
rect 151983 995938 151988 995994
rect 152044 995938 152544 995994
rect 151983 995936 152544 995938
rect 152847 995994 153408 995996
rect 152847 995938 152852 995994
rect 152908 995938 153408 995994
rect 152847 995936 153408 995938
rect 155343 995994 155712 995996
rect 155343 995938 155348 995994
rect 155404 995938 155712 995994
rect 155343 995936 155712 995938
rect 163680 995994 164241 995996
rect 163680 995938 164180 995994
rect 164236 995938 164241 995994
rect 163680 995936 164241 995938
rect 149487 995933 149553 995936
rect 151983 995933 152049 995936
rect 152847 995933 152913 995936
rect 155343 995933 155409 995936
rect 164175 995933 164241 995936
rect 185922 995994 198705 995996
rect 185922 995938 198644 995994
rect 198700 995938 198705 995994
rect 185922 995936 198705 995938
rect 87855 995848 87921 995851
rect 92559 995848 92625 995851
rect 113391 995848 113457 995851
rect 87855 995846 92625 995848
rect 87855 995790 87860 995846
rect 87916 995790 92564 995846
rect 92620 995790 92625 995846
rect 87855 995788 92625 995790
rect 87855 995785 87921 995788
rect 92559 995785 92625 995788
rect 85935 995700 86001 995703
rect 92655 995700 92721 995703
rect 85935 995698 92721 995700
rect 85935 995642 85940 995698
rect 85996 995642 92660 995698
rect 92716 995642 92721 995698
rect 85935 995640 92721 995642
rect 85935 995637 86001 995640
rect 92655 995637 92721 995640
rect 94959 995700 95025 995703
rect 97218 995700 97278 995818
rect 98754 995700 98814 995818
rect 94959 995698 98814 995700
rect 94959 995642 94964 995698
rect 95020 995642 98814 995698
rect 94959 995640 98814 995642
rect 94959 995637 95025 995640
rect 86511 995552 86577 995555
rect 99522 995552 99582 995818
rect 86511 995550 99582 995552
rect 86511 995494 86516 995550
rect 86572 995494 99582 995550
rect 86511 995492 99582 995494
rect 86511 995489 86577 995492
rect 85359 995404 85425 995407
rect 100386 995404 100446 995818
rect 85359 995402 100446 995404
rect 85359 995346 85364 995402
rect 85420 995346 100446 995402
rect 85359 995344 100446 995346
rect 85359 995341 85425 995344
rect 80751 995256 80817 995259
rect 99759 995256 99825 995259
rect 80751 995254 99825 995256
rect 80751 995198 80756 995254
rect 80812 995198 99764 995254
rect 99820 995198 99825 995254
rect 80751 995196 99825 995198
rect 80751 995193 80817 995196
rect 99759 995193 99825 995196
rect 84495 993924 84561 993927
rect 106722 993924 106782 995818
rect 108258 995407 108318 995818
rect 108207 995402 108318 995407
rect 108207 995346 108212 995402
rect 108268 995346 108318 995402
rect 108207 995344 108318 995346
rect 108207 995341 108273 995344
rect 109890 995259 109950 995818
rect 110688 995788 111294 995848
rect 112992 995846 113457 995848
rect 111234 995404 111294 995788
rect 111522 995552 111582 995818
rect 112194 995700 112254 995818
rect 112992 995790 113396 995846
rect 113452 995790 113457 995846
rect 112992 995788 113457 995790
rect 113391 995785 113457 995788
rect 136719 995846 136830 995851
rect 136719 995790 136724 995846
rect 136780 995790 136830 995846
rect 136719 995788 136830 995790
rect 137967 995848 138033 995851
rect 143919 995848 143985 995851
rect 137967 995846 143985 995848
rect 137967 995790 137972 995846
rect 138028 995790 143924 995846
rect 143980 995790 143985 995846
rect 154287 995848 154353 995851
rect 156303 995848 156369 995851
rect 165615 995848 165681 995851
rect 166191 995848 166257 995851
rect 185103 995848 185169 995851
rect 185922 995848 185982 995936
rect 198639 995933 198705 995936
rect 200898 995936 201504 995996
rect 203439 995994 204000 995996
rect 203439 995938 203444 995994
rect 203500 995938 204000 995994
rect 203439 995936 204000 995938
rect 205647 995994 206304 995996
rect 205647 995938 205652 995994
rect 205708 995938 206304 995994
rect 205647 995936 206304 995938
rect 206511 995994 207072 995996
rect 206511 995938 206516 995994
rect 206572 995938 207072 995994
rect 206511 995936 207072 995938
rect 215439 995994 215808 995996
rect 215439 995938 215444 995994
rect 215500 995938 215808 995994
rect 215439 995936 215808 995938
rect 217071 995994 217440 995996
rect 217071 995938 217076 995994
rect 217132 995938 217440 995994
rect 217071 995936 217440 995938
rect 218304 995994 221841 995996
rect 218304 995938 221780 995994
rect 221836 995938 221841 995994
rect 218304 995936 221841 995938
rect 154287 995846 154944 995848
rect 137967 995788 143985 995790
rect 136719 995785 136785 995788
rect 137967 995785 138033 995788
rect 143919 995785 143985 995788
rect 137583 995700 137649 995703
rect 112194 995698 137649 995700
rect 112194 995642 137588 995698
rect 137644 995642 137649 995698
rect 112194 995640 137649 995642
rect 137583 995637 137649 995640
rect 139215 995700 139281 995703
rect 139215 995698 153342 995700
rect 139215 995642 139220 995698
rect 139276 995642 153342 995698
rect 139215 995640 153342 995642
rect 139215 995637 139281 995640
rect 115215 995552 115281 995555
rect 111522 995550 115281 995552
rect 111522 995494 115220 995550
rect 115276 995494 115281 995550
rect 111522 995492 115281 995494
rect 115215 995489 115281 995492
rect 137391 995552 137457 995555
rect 152847 995552 152913 995555
rect 137391 995550 152913 995552
rect 137391 995494 137396 995550
rect 137452 995494 152852 995550
rect 152908 995494 152913 995550
rect 137391 995492 152913 995494
rect 153282 995552 153342 995640
rect 154050 995552 154110 995818
rect 154287 995790 154292 995846
rect 154348 995790 154944 995846
rect 154287 995788 154944 995790
rect 156303 995846 156576 995848
rect 156303 995790 156308 995846
rect 156364 995790 156576 995846
rect 156303 995788 156576 995790
rect 154287 995785 154353 995788
rect 156303 995785 156369 995788
rect 158850 995555 158910 995818
rect 159618 995703 159678 995818
rect 159567 995698 159678 995703
rect 159567 995642 159572 995698
rect 159628 995642 159678 995698
rect 159567 995640 159678 995642
rect 159567 995637 159633 995640
rect 153282 995492 154110 995552
rect 158799 995550 158910 995555
rect 158799 995494 158804 995550
rect 158860 995494 158910 995550
rect 158799 995492 158910 995494
rect 158991 995552 159057 995555
rect 161250 995552 161310 995818
rect 165216 995788 165438 995848
rect 165378 995700 165438 995788
rect 165615 995846 166080 995848
rect 165615 995790 165620 995846
rect 165676 995790 166080 995846
rect 165615 995788 166080 995790
rect 166191 995846 166944 995848
rect 166191 995790 166196 995846
rect 166252 995790 166944 995846
rect 166191 995788 166944 995790
rect 185103 995846 185982 995848
rect 185103 995790 185108 995846
rect 185164 995790 185982 995846
rect 185103 995788 185982 995790
rect 188751 995848 188817 995851
rect 195183 995848 195249 995851
rect 188751 995846 195249 995848
rect 188751 995790 188756 995846
rect 188812 995790 195188 995846
rect 195244 995790 195249 995846
rect 188751 995788 195249 995790
rect 165615 995785 165681 995788
rect 166191 995785 166257 995788
rect 185103 995785 185169 995788
rect 188751 995785 188817 995788
rect 195183 995785 195249 995788
rect 170319 995700 170385 995703
rect 165378 995698 170385 995700
rect 165378 995642 170324 995698
rect 170380 995642 170385 995698
rect 165378 995640 170385 995642
rect 170319 995637 170385 995640
rect 178479 995700 178545 995703
rect 185199 995700 185265 995703
rect 178479 995698 185265 995700
rect 178479 995642 178484 995698
rect 178540 995642 185204 995698
rect 185260 995642 185265 995698
rect 178479 995640 185265 995642
rect 178479 995637 178545 995640
rect 185199 995637 185265 995640
rect 195087 995700 195153 995703
rect 200034 995700 200094 995818
rect 200898 995700 200958 995936
rect 203439 995933 203505 995936
rect 205647 995933 205713 995936
rect 206511 995933 206577 995936
rect 215439 995933 215505 995936
rect 217071 995933 217137 995936
rect 221775 995933 221841 995936
rect 243714 995994 246993 995996
rect 243714 995938 246932 995994
rect 246988 995938 246993 995994
rect 243714 995936 246993 995938
rect 201711 995848 201777 995851
rect 202863 995848 202929 995851
rect 204975 995848 205041 995851
rect 241839 995848 241905 995851
rect 243714 995848 243774 995936
rect 246927 995933 246993 995936
rect 247503 995996 247569 995999
rect 258831 995996 258897 995999
rect 264687 995996 264753 995999
rect 298383 995996 298449 995999
rect 247503 995994 251424 995996
rect 247503 995938 247508 995994
rect 247564 995966 251424 995994
rect 258831 995994 259296 995996
rect 247564 995938 251454 995966
rect 247503 995936 251454 995938
rect 247503 995933 247569 995936
rect 201711 995846 202368 995848
rect 201711 995790 201716 995846
rect 201772 995790 202368 995846
rect 201711 995788 202368 995790
rect 202863 995846 203232 995848
rect 202863 995790 202868 995846
rect 202924 995790 203232 995846
rect 202863 995788 203232 995790
rect 204975 995846 205536 995848
rect 204975 995790 204980 995846
rect 205036 995790 205536 995846
rect 241839 995846 243774 995848
rect 204975 995788 205536 995790
rect 201711 995785 201777 995788
rect 202863 995785 202929 995788
rect 204975 995785 205041 995788
rect 195087 995698 200958 995700
rect 195087 995642 195092 995698
rect 195148 995642 200958 995698
rect 195087 995640 200958 995642
rect 206991 995700 207057 995703
rect 207906 995700 207966 995818
rect 206991 995698 207966 995700
rect 206991 995642 206996 995698
rect 207052 995642 207966 995698
rect 206991 995640 207966 995642
rect 195087 995637 195153 995640
rect 206991 995637 207057 995640
rect 158991 995550 161310 995552
rect 158991 995494 158996 995550
rect 159052 995494 161310 995550
rect 158991 995492 161310 995494
rect 184335 995552 184401 995555
rect 189423 995552 189489 995555
rect 201711 995552 201777 995555
rect 184335 995550 189246 995552
rect 184335 995494 184340 995550
rect 184396 995494 189246 995550
rect 184335 995492 189246 995494
rect 137391 995489 137457 995492
rect 152847 995489 152913 995492
rect 158799 995489 158865 995492
rect 158991 995489 159057 995492
rect 184335 995489 184401 995492
rect 115311 995404 115377 995407
rect 111234 995402 115377 995404
rect 111234 995346 115316 995402
rect 115372 995346 115377 995402
rect 111234 995344 115377 995346
rect 115311 995341 115377 995344
rect 140367 995404 140433 995407
rect 141135 995404 141201 995407
rect 140367 995402 141201 995404
rect 140367 995346 140372 995402
rect 140428 995346 141140 995402
rect 141196 995346 141201 995402
rect 140367 995344 141201 995346
rect 189186 995404 189246 995492
rect 189423 995550 201777 995552
rect 189423 995494 189428 995550
rect 189484 995494 201716 995550
rect 201772 995494 201777 995550
rect 189423 995492 201777 995494
rect 189423 995489 189489 995492
rect 201711 995489 201777 995492
rect 210210 995407 210270 995818
rect 211074 995407 211134 995818
rect 212706 995407 212766 995818
rect 216642 995700 216702 995818
rect 241839 995790 241844 995846
rect 241900 995790 243774 995846
rect 241839 995788 243774 995790
rect 243855 995848 243921 995851
rect 251247 995848 251313 995851
rect 243855 995846 251313 995848
rect 243855 995790 243860 995846
rect 243916 995790 251252 995846
rect 251308 995790 251313 995846
rect 251394 995848 251454 995936
rect 258831 995938 258836 995994
rect 258892 995938 259296 995994
rect 258831 995936 259296 995938
rect 264687 995994 264864 995996
rect 264687 995938 264692 995994
rect 264748 995938 264864 995994
rect 264687 995936 264864 995938
rect 294594 995994 298449 995996
rect 294594 995938 298388 995994
rect 298444 995938 298449 995994
rect 294594 995936 298449 995938
rect 258831 995933 258897 995936
rect 264687 995933 264753 995936
rect 254799 995848 254865 995851
rect 255567 995848 255633 995851
rect 257487 995848 257553 995851
rect 258255 995848 258321 995851
rect 260751 995848 260817 995851
rect 268239 995848 268305 995851
rect 251394 995818 251838 995848
rect 243855 995788 251313 995790
rect 251424 995788 251838 995818
rect 241839 995785 241905 995788
rect 243855 995785 243921 995788
rect 251247 995785 251313 995788
rect 222927 995700 222993 995703
rect 216642 995698 222993 995700
rect 216642 995642 222932 995698
rect 222988 995642 222993 995698
rect 216642 995640 222993 995642
rect 222927 995637 222993 995640
rect 240783 995700 240849 995703
rect 251778 995700 251838 995788
rect 252930 995700 252990 995818
rect 253728 995788 253950 995848
rect 254799 995846 255456 995848
rect 253890 995700 253950 995788
rect 240783 995698 250494 995700
rect 240783 995642 240788 995698
rect 240844 995642 250494 995698
rect 240783 995640 250494 995642
rect 251778 995640 252990 995700
rect 253698 995640 253950 995700
rect 240783 995637 240849 995640
rect 239535 995552 239601 995555
rect 250434 995552 250494 995640
rect 253698 995552 253758 995640
rect 239535 995550 250302 995552
rect 239535 995494 239540 995550
rect 239596 995494 250302 995550
rect 239535 995492 250302 995494
rect 250434 995492 253758 995552
rect 239535 995489 239601 995492
rect 205647 995404 205713 995407
rect 189186 995402 205713 995404
rect 189186 995346 205652 995402
rect 205708 995346 205713 995402
rect 189186 995344 205713 995346
rect 210210 995402 210321 995407
rect 210210 995346 210260 995402
rect 210316 995346 210321 995402
rect 210210 995344 210321 995346
rect 140367 995341 140433 995344
rect 141135 995341 141201 995344
rect 205647 995341 205713 995344
rect 210255 995341 210321 995344
rect 211023 995402 211134 995407
rect 211023 995346 211028 995402
rect 211084 995346 211134 995402
rect 211023 995344 211134 995346
rect 212655 995402 212766 995407
rect 212655 995346 212660 995402
rect 212716 995346 212766 995402
rect 212655 995344 212766 995346
rect 240207 995404 240273 995407
rect 250095 995404 250161 995407
rect 240207 995402 250161 995404
rect 240207 995346 240212 995402
rect 240268 995346 250100 995402
rect 250156 995346 250161 995402
rect 240207 995344 250161 995346
rect 250242 995404 250302 995492
rect 254562 995404 254622 995818
rect 254799 995790 254804 995846
rect 254860 995790 255456 995846
rect 254799 995788 255456 995790
rect 255567 995846 256224 995848
rect 255567 995790 255572 995846
rect 255628 995790 256224 995846
rect 255567 995788 256224 995790
rect 257487 995846 257760 995848
rect 257487 995790 257492 995846
rect 257548 995790 257760 995846
rect 257487 995788 257760 995790
rect 258255 995846 258528 995848
rect 258255 995790 258260 995846
rect 258316 995790 258528 995846
rect 258255 995788 258528 995790
rect 260751 995846 261024 995848
rect 260751 995790 260756 995846
rect 260812 995790 261024 995846
rect 260751 995788 261024 995790
rect 261600 995788 261822 995848
rect 268032 995846 268305 995848
rect 254799 995785 254865 995788
rect 255567 995785 255633 995788
rect 257487 995785 257553 995788
rect 258255 995785 258321 995788
rect 260751 995785 260817 995788
rect 261762 995700 261822 995788
rect 262434 995703 262494 995818
rect 261570 995640 261822 995700
rect 262383 995698 262494 995703
rect 262383 995642 262388 995698
rect 262444 995642 262494 995698
rect 262383 995640 262494 995642
rect 250242 995344 254622 995404
rect 254703 995404 254769 995407
rect 261570 995404 261630 995640
rect 262383 995637 262449 995640
rect 264066 995407 264126 995818
rect 266370 995700 266430 995818
rect 268032 995790 268244 995846
rect 268300 995790 268305 995846
rect 268032 995788 268305 995790
rect 268239 995785 268305 995788
rect 268431 995848 268497 995851
rect 273615 995848 273681 995851
rect 268431 995846 268896 995848
rect 268431 995790 268436 995846
rect 268492 995790 268896 995846
rect 268431 995788 268896 995790
rect 269664 995846 273681 995848
rect 269664 995790 273620 995846
rect 273676 995790 273681 995846
rect 269664 995788 273681 995790
rect 268431 995785 268497 995788
rect 273615 995785 273681 995788
rect 283119 995848 283185 995851
rect 294594 995848 294654 995936
rect 298383 995933 298449 995936
rect 305583 995996 305649 995999
rect 316335 995996 316401 995999
rect 328239 995996 328305 995999
rect 362319 995996 362385 995999
rect 367119 995996 367185 995999
rect 377295 995996 377361 995999
rect 305583 995994 306144 995996
rect 305583 995938 305588 995994
rect 305644 995938 306144 995994
rect 305583 995936 306144 995938
rect 316335 995994 316512 995996
rect 316335 995938 316340 995994
rect 316396 995938 316512 995994
rect 316335 995936 316512 995938
rect 321312 995994 328305 995996
rect 321312 995938 328244 995994
rect 328300 995938 328305 995994
rect 321312 995936 328305 995938
rect 362208 995994 362385 995996
rect 362208 995938 362324 995994
rect 362380 995938 362385 995994
rect 362208 995936 362385 995938
rect 366912 995994 367185 995996
rect 366912 995938 367124 995994
rect 367180 995938 367185 995994
rect 366912 995936 367185 995938
rect 371712 995994 377361 995996
rect 371712 995938 377300 995994
rect 377356 995938 377361 995994
rect 371712 995936 377361 995938
rect 305583 995933 305649 995936
rect 316335 995933 316401 995936
rect 328239 995933 328305 995936
rect 362319 995933 362385 995936
rect 367119 995933 367185 995936
rect 377295 995933 377361 995936
rect 379311 995996 379377 995999
rect 379311 995994 391422 995996
rect 379311 995938 379316 995994
rect 379372 995938 391422 995994
rect 379311 995936 391422 995938
rect 379311 995933 379377 995936
rect 283119 995846 294654 995848
rect 283119 995790 283124 995846
rect 283180 995790 294654 995846
rect 283119 995788 294654 995790
rect 294831 995848 294897 995851
rect 298287 995848 298353 995851
rect 306447 995848 306513 995851
rect 307407 995848 307473 995851
rect 311919 995848 311985 995851
rect 348687 995848 348753 995851
rect 365871 995848 365937 995851
rect 366639 995848 366705 995851
rect 294831 995846 298353 995848
rect 294831 995790 294836 995846
rect 294892 995790 298292 995846
rect 298348 995790 298353 995846
rect 294831 995788 298353 995790
rect 283119 995785 283185 995788
rect 294831 995785 294897 995788
rect 298287 995785 298353 995788
rect 270735 995700 270801 995703
rect 266370 995698 270801 995700
rect 266370 995642 270740 995698
rect 270796 995642 270801 995698
rect 266370 995640 270801 995642
rect 270735 995637 270801 995640
rect 286287 995700 286353 995703
rect 298479 995700 298545 995703
rect 286287 995698 298545 995700
rect 286287 995642 286292 995698
rect 286348 995642 298484 995698
rect 298540 995642 298545 995698
rect 286287 995640 298545 995642
rect 286287 995637 286353 995640
rect 298479 995637 298545 995640
rect 299151 995700 299217 995703
rect 303042 995700 303102 995818
rect 304002 995788 304608 995848
rect 306447 995846 307008 995848
rect 304002 995700 304062 995788
rect 299151 995698 304062 995700
rect 299151 995642 299156 995698
rect 299212 995642 304062 995698
rect 299151 995640 304062 995642
rect 299151 995637 299217 995640
rect 292527 995552 292593 995555
rect 305346 995552 305406 995818
rect 306447 995790 306452 995846
rect 306508 995790 307008 995846
rect 306447 995788 307008 995790
rect 307407 995846 307872 995848
rect 307407 995790 307412 995846
rect 307468 995790 307872 995846
rect 307407 995788 307872 995790
rect 311919 995846 312576 995848
rect 311919 995790 311924 995846
rect 311980 995790 312576 995846
rect 348687 995846 353472 995848
rect 311919 995788 312576 995790
rect 306447 995785 306513 995788
rect 307407 995785 307473 995788
rect 311919 995785 311985 995788
rect 319650 995700 319710 995818
rect 348687 995790 348692 995846
rect 348748 995818 353472 995846
rect 348748 995790 353502 995818
rect 348687 995788 353502 995790
rect 354912 995788 355134 995848
rect 365280 995846 365937 995848
rect 348687 995785 348753 995788
rect 325263 995700 325329 995703
rect 319650 995698 325329 995700
rect 319650 995642 325268 995698
rect 325324 995642 325329 995698
rect 319650 995640 325329 995642
rect 353442 995700 353502 995788
rect 355074 995700 355134 995788
rect 353442 995640 355134 995700
rect 325263 995637 325329 995640
rect 292527 995550 305406 995552
rect 292527 995494 292532 995550
rect 292588 995494 305406 995550
rect 292527 995492 305406 995494
rect 292527 995489 292593 995492
rect 254703 995402 261630 995404
rect 254703 995346 254708 995402
rect 254764 995346 261630 995402
rect 254703 995344 261630 995346
rect 264015 995402 264126 995407
rect 264015 995346 264020 995402
rect 264076 995346 264126 995402
rect 264015 995344 264126 995346
rect 362946 995404 363006 995818
rect 365280 995790 365876 995846
rect 365932 995790 365937 995846
rect 365280 995788 365937 995790
rect 366048 995846 366705 995848
rect 366048 995790 366644 995846
rect 366700 995790 366705 995846
rect 371823 995848 371889 995851
rect 385839 995848 385905 995851
rect 389103 995848 389169 995851
rect 371823 995846 385905 995848
rect 366048 995788 366705 995790
rect 365871 995785 365937 995788
rect 366639 995785 366705 995788
rect 368418 995700 368478 995818
rect 368655 995700 368721 995703
rect 368418 995698 368721 995700
rect 368418 995642 368660 995698
rect 368716 995642 368721 995698
rect 368418 995640 368721 995642
rect 368655 995637 368721 995640
rect 370050 995552 370110 995818
rect 370818 995700 370878 995818
rect 371823 995790 371828 995846
rect 371884 995790 385844 995846
rect 385900 995790 385905 995846
rect 371823 995788 385905 995790
rect 371823 995785 371889 995788
rect 385839 995785 385905 995788
rect 385986 995846 389169 995848
rect 385986 995790 389108 995846
rect 389164 995790 389169 995846
rect 385986 995788 389169 995790
rect 391362 995848 391422 995936
rect 393711 995848 393777 995851
rect 391362 995846 393777 995848
rect 391362 995790 393716 995846
rect 393772 995790 393777 995846
rect 391362 995788 393777 995790
rect 374415 995700 374481 995703
rect 370818 995698 374481 995700
rect 370818 995642 374420 995698
rect 374476 995642 374481 995698
rect 370818 995640 374481 995642
rect 374415 995637 374481 995640
rect 381711 995700 381777 995703
rect 385986 995700 386046 995788
rect 389103 995785 389169 995788
rect 393711 995785 393777 995788
rect 389391 995700 389457 995703
rect 381711 995698 386046 995700
rect 381711 995642 381716 995698
rect 381772 995642 386046 995698
rect 381711 995640 386046 995642
rect 386178 995698 389457 995700
rect 386178 995642 389396 995698
rect 389452 995642 389457 995698
rect 386178 995640 389457 995642
rect 381711 995637 381777 995640
rect 374511 995552 374577 995555
rect 370050 995550 374577 995552
rect 370050 995494 374516 995550
rect 374572 995494 374577 995550
rect 370050 995492 374577 995494
rect 374511 995489 374577 995492
rect 380271 995552 380337 995555
rect 386178 995552 386238 995640
rect 389391 995637 389457 995640
rect 380271 995550 386238 995552
rect 380271 995494 380276 995550
rect 380332 995494 386238 995550
rect 380271 995492 386238 995494
rect 386319 995552 386385 995555
rect 391791 995552 391857 995555
rect 386319 995550 391857 995552
rect 386319 995494 386324 995550
rect 386380 995494 391796 995550
rect 391852 995494 391857 995550
rect 386319 995492 391857 995494
rect 418818 995552 418878 996084
rect 436431 996081 436497 996084
rect 511119 996144 511185 996147
rect 513423 996144 513489 996147
rect 517167 996144 517233 996147
rect 511119 996142 511296 996144
rect 511119 996086 511124 996142
rect 511180 996086 511296 996142
rect 511119 996084 511296 996086
rect 513423 996142 513696 996144
rect 513423 996086 513428 996142
rect 513484 996086 513696 996142
rect 513423 996084 513696 996086
rect 517167 996142 532734 996144
rect 517167 996086 517172 996142
rect 517228 996086 532734 996142
rect 517167 996084 532734 996086
rect 511119 996081 511185 996084
rect 513423 996081 513489 996084
rect 517167 996081 517233 996084
rect 429711 995996 429777 995999
rect 429600 995994 429777 995996
rect 429600 995938 429716 995994
rect 429772 995938 429777 995994
rect 429600 995936 429777 995938
rect 429711 995933 429777 995936
rect 434127 995996 434193 995999
rect 446223 995996 446289 995999
rect 434127 995994 434304 995996
rect 434127 995938 434132 995994
rect 434188 995938 434304 995994
rect 434127 995936 434304 995938
rect 439104 995994 446289 995996
rect 439104 995938 446228 995994
rect 446284 995938 446289 995994
rect 439104 995936 446289 995938
rect 434127 995933 434193 995936
rect 446223 995933 446289 995936
rect 471855 995996 471921 995999
rect 511887 995996 511953 995999
rect 513327 995996 513393 995999
rect 521391 995996 521457 995999
rect 471855 995994 477822 995996
rect 471855 995938 471860 995994
rect 471916 995938 477822 995994
rect 471855 995936 477822 995938
rect 471855 995933 471921 995936
rect 422511 995848 422577 995851
rect 438735 995848 438801 995851
rect 422304 995846 422656 995848
rect 420834 995700 420894 995818
rect 422304 995790 422516 995846
rect 422572 995790 422656 995846
rect 438240 995846 438801 995848
rect 422304 995788 422656 995790
rect 422466 995785 422577 995788
rect 422466 995700 422526 995785
rect 420834 995640 422526 995700
rect 437442 995700 437502 995818
rect 438240 995790 438740 995846
rect 438796 995790 438801 995846
rect 438240 995788 438801 995790
rect 438735 995785 438801 995788
rect 472239 995848 472305 995851
rect 477039 995848 477105 995851
rect 472239 995846 477105 995848
rect 472239 995790 472244 995846
rect 472300 995790 477044 995846
rect 477100 995790 477105 995846
rect 472239 995788 477105 995790
rect 477762 995848 477822 995936
rect 511887 995994 512160 995996
rect 511887 995938 511892 995994
rect 511948 995938 512160 995994
rect 511887 995936 512160 995938
rect 512832 995994 513393 995996
rect 512832 995938 513332 995994
rect 513388 995938 513393 995994
rect 512832 995936 513393 995938
rect 516096 995994 521457 995996
rect 516096 995938 521396 995994
rect 521452 995938 521457 995994
rect 516096 995936 521457 995938
rect 511887 995933 511953 995936
rect 513327 995933 513393 995936
rect 521391 995933 521457 995936
rect 521583 995996 521649 995999
rect 521583 995994 528126 995996
rect 521583 995938 521588 995994
rect 521644 995938 528126 995994
rect 521583 995936 528126 995938
rect 521583 995933 521649 995936
rect 485775 995848 485841 995851
rect 504687 995848 504753 995851
rect 523983 995848 524049 995851
rect 527919 995848 527985 995851
rect 477762 995846 485841 995848
rect 477762 995790 485780 995846
rect 485836 995790 485841 995846
rect 477762 995788 485841 995790
rect 504096 995846 504753 995848
rect 504096 995790 504692 995846
rect 504748 995790 504753 995846
rect 504096 995788 504753 995790
rect 472239 995785 472305 995788
rect 477039 995785 477105 995788
rect 485775 995785 485841 995788
rect 504687 995785 504753 995788
rect 440751 995700 440817 995703
rect 437442 995698 440817 995700
rect 437442 995642 440756 995698
rect 440812 995642 440817 995698
rect 437442 995640 440817 995642
rect 440751 995637 440817 995640
rect 467055 995700 467121 995703
rect 480975 995700 481041 995703
rect 467055 995698 481041 995700
rect 467055 995642 467060 995698
rect 467116 995642 480980 995698
rect 481036 995642 481041 995698
rect 467055 995640 481041 995642
rect 467055 995637 467121 995640
rect 480975 995637 481041 995640
rect 472143 995552 472209 995555
rect 478383 995552 478449 995555
rect 418818 995492 429054 995552
rect 380271 995489 380337 995492
rect 386319 995489 386385 995492
rect 391791 995489 391857 995492
rect 377391 995404 377457 995407
rect 396687 995404 396753 995407
rect 362946 995344 372990 995404
rect 211023 995341 211089 995344
rect 212655 995341 212721 995344
rect 240207 995341 240273 995344
rect 250095 995341 250161 995344
rect 254703 995341 254769 995344
rect 264015 995341 264081 995344
rect 109839 995254 109950 995259
rect 109839 995198 109844 995254
rect 109900 995198 109950 995254
rect 109839 995196 109950 995198
rect 161199 995256 161265 995259
rect 166959 995256 167025 995259
rect 161199 995254 167025 995256
rect 161199 995198 161204 995254
rect 161260 995198 166964 995254
rect 167020 995198 167025 995254
rect 161199 995196 167025 995198
rect 109839 995193 109905 995196
rect 161199 995193 161265 995196
rect 166959 995193 167025 995196
rect 183759 995256 183825 995259
rect 201711 995256 201777 995259
rect 183759 995254 201777 995256
rect 183759 995198 183764 995254
rect 183820 995198 201716 995254
rect 201772 995198 201777 995254
rect 183759 995196 201777 995198
rect 183759 995193 183825 995196
rect 201711 995193 201777 995196
rect 316719 995256 316785 995259
rect 339759 995256 339825 995259
rect 362799 995256 362865 995259
rect 368463 995256 368529 995259
rect 316719 995254 319710 995256
rect 316719 995198 316724 995254
rect 316780 995198 319710 995254
rect 316719 995196 319710 995198
rect 316719 995193 316785 995196
rect 167151 995108 167217 995111
rect 181455 995108 181521 995111
rect 167151 995106 181521 995108
rect 167151 995050 167156 995106
rect 167212 995050 181460 995106
rect 181516 995050 181521 995106
rect 167151 995048 181521 995050
rect 167151 995045 167217 995048
rect 181455 995045 181521 995048
rect 201519 995108 201585 995111
rect 227343 995108 227409 995111
rect 201519 995106 201726 995108
rect 201519 995050 201524 995106
rect 201580 995050 201726 995106
rect 201519 995048 201726 995050
rect 201519 995045 201585 995048
rect 201666 994960 201726 995048
rect 221634 995106 227409 995108
rect 221634 995050 227348 995106
rect 227404 995050 227409 995106
rect 221634 995048 227409 995050
rect 221634 994960 221694 995048
rect 227343 995045 227409 995048
rect 227535 995108 227601 995111
rect 247407 995108 247473 995111
rect 227535 995106 247473 995108
rect 227535 995050 227540 995106
rect 227596 995050 247412 995106
rect 247468 995050 247473 995106
rect 227535 995048 247473 995050
rect 227535 995045 227601 995048
rect 247407 995045 247473 995048
rect 259119 995108 259185 995111
rect 262191 995108 262257 995111
rect 316719 995108 316785 995111
rect 259119 995106 262257 995108
rect 259119 995050 259124 995106
rect 259180 995050 262196 995106
rect 262252 995050 262257 995106
rect 259119 995048 262257 995050
rect 259119 995045 259185 995048
rect 262191 995045 262257 995048
rect 296658 995106 316785 995108
rect 296658 995050 316724 995106
rect 316780 995050 316785 995106
rect 296658 995048 316785 995050
rect 201666 994900 221694 994960
rect 262191 994812 262257 994815
rect 296658 994812 296718 995048
rect 316719 995045 316785 995048
rect 319650 994960 319710 995196
rect 339759 995254 342846 995256
rect 339759 995198 339764 995254
rect 339820 995198 342846 995254
rect 339759 995196 342846 995198
rect 339759 995193 339825 995196
rect 342786 995108 342846 995196
rect 362799 995254 368529 995256
rect 362799 995198 362804 995254
rect 362860 995198 368468 995254
rect 368524 995198 368529 995254
rect 362799 995196 368529 995198
rect 372930 995256 372990 995344
rect 377391 995402 396753 995404
rect 377391 995346 377396 995402
rect 377452 995346 396692 995402
rect 396748 995346 396753 995402
rect 377391 995344 396753 995346
rect 377391 995341 377457 995344
rect 396687 995341 396753 995344
rect 386319 995256 386385 995259
rect 372930 995254 386385 995256
rect 372930 995198 386324 995254
rect 386380 995198 386385 995254
rect 372930 995196 386385 995198
rect 428994 995256 429054 995492
rect 472143 995550 478449 995552
rect 472143 995494 472148 995550
rect 472204 995494 478388 995550
rect 478444 995494 478449 995550
rect 472143 995492 478449 995494
rect 472143 995489 472209 995492
rect 478383 995489 478449 995492
rect 479919 995552 479985 995555
rect 488847 995552 488913 995555
rect 479919 995550 488913 995552
rect 479919 995494 479924 995550
rect 479980 995494 488852 995550
rect 488908 995494 488913 995550
rect 479919 995492 488913 995494
rect 479919 995489 479985 995492
rect 488847 995489 488913 995492
rect 463599 995404 463665 995407
rect 471759 995404 471825 995407
rect 482031 995404 482097 995407
rect 463599 995402 469566 995404
rect 463599 995346 463604 995402
rect 463660 995346 469566 995402
rect 463599 995344 469566 995346
rect 463599 995341 463665 995344
rect 443535 995256 443601 995259
rect 428994 995254 443601 995256
rect 428994 995198 443540 995254
rect 443596 995198 443601 995254
rect 428994 995196 443601 995198
rect 469506 995256 469566 995344
rect 471759 995402 482097 995404
rect 471759 995346 471764 995402
rect 471820 995346 482036 995402
rect 482092 995346 482097 995402
rect 471759 995344 482097 995346
rect 471759 995341 471825 995344
rect 482031 995341 482097 995344
rect 506562 995259 506622 995818
rect 510498 995404 510558 995818
rect 514434 995552 514494 995818
rect 515232 995788 515838 995848
rect 515778 995700 515838 995788
rect 523983 995846 527985 995848
rect 523983 995790 523988 995846
rect 524044 995790 527924 995846
rect 527980 995790 527985 995846
rect 523983 995788 527985 995790
rect 528066 995848 528126 995936
rect 532239 995848 532305 995851
rect 528066 995846 532305 995848
rect 528066 995790 532244 995846
rect 532300 995790 532305 995846
rect 528066 995788 532305 995790
rect 532674 995848 532734 996084
rect 562863 995996 562929 995999
rect 562752 995994 562929 995996
rect 562752 995938 562868 995994
rect 562924 995938 562929 995994
rect 562752 995936 562929 995938
rect 562863 995933 562929 995936
rect 564783 995996 564849 995999
rect 567087 995996 567153 995999
rect 564783 995994 565056 995996
rect 564783 995938 564788 995994
rect 564844 995938 565056 995994
rect 564783 995936 565056 995938
rect 566688 995994 567153 995996
rect 566688 995938 567092 995994
rect 567148 995938 567153 995994
rect 566688 995936 567153 995938
rect 564783 995933 564849 995936
rect 567087 995933 567153 995936
rect 624879 995996 624945 995999
rect 624879 995994 634110 995996
rect 624879 995938 624884 995994
rect 624940 995938 634110 995994
rect 624879 995936 634110 995938
rect 624879 995933 624945 995936
rect 634050 995851 634110 995936
rect 535311 995848 535377 995851
rect 558159 995848 558225 995851
rect 563727 995848 563793 995851
rect 566319 995848 566385 995851
rect 573135 995848 573201 995851
rect 532674 995846 535377 995848
rect 532674 995790 535316 995846
rect 535372 995790 535377 995846
rect 532674 995788 535377 995790
rect 549216 995788 549438 995848
rect 523983 995785 524049 995788
rect 527919 995785 527985 995788
rect 532239 995785 532305 995788
rect 535311 995785 535377 995788
rect 518511 995700 518577 995703
rect 515778 995698 518577 995700
rect 515778 995642 518516 995698
rect 518572 995642 518577 995698
rect 515778 995640 518577 995642
rect 518511 995637 518577 995640
rect 518703 995700 518769 995703
rect 529071 995700 529137 995703
rect 534063 995700 534129 995703
rect 518703 995698 529137 995700
rect 518703 995642 518708 995698
rect 518764 995642 529076 995698
rect 529132 995642 529137 995698
rect 518703 995640 529137 995642
rect 518703 995637 518769 995640
rect 529071 995637 529137 995640
rect 529218 995698 534129 995700
rect 529218 995642 534068 995698
rect 534124 995642 534129 995698
rect 529218 995640 534129 995642
rect 518703 995552 518769 995555
rect 514434 995550 518769 995552
rect 514434 995494 518708 995550
rect 518764 995494 518769 995550
rect 514434 995492 518769 995494
rect 518703 995489 518769 995492
rect 521487 995552 521553 995555
rect 529218 995552 529278 995640
rect 534063 995637 534129 995640
rect 544239 995700 544305 995703
rect 549378 995700 549438 995788
rect 550722 995700 550782 995818
rect 551520 995788 551742 995848
rect 557952 995846 558225 995848
rect 557952 995790 558164 995846
rect 558220 995790 558225 995846
rect 557952 995788 558225 995790
rect 563520 995846 563793 995848
rect 563520 995790 563732 995846
rect 563788 995790 563793 995846
rect 563520 995788 563793 995790
rect 565824 995846 566385 995848
rect 565824 995790 566324 995846
rect 566380 995790 566385 995846
rect 565824 995788 566385 995790
rect 567456 995846 573201 995848
rect 567456 995790 573140 995846
rect 573196 995790 573201 995846
rect 567456 995788 573201 995790
rect 634050 995846 634161 995851
rect 634050 995790 634100 995846
rect 634156 995790 634161 995846
rect 634050 995788 634161 995790
rect 544239 995698 550782 995700
rect 544239 995642 544244 995698
rect 544300 995642 550782 995698
rect 544239 995640 550782 995642
rect 551682 995700 551742 995788
rect 558159 995785 558225 995788
rect 563727 995785 563793 995788
rect 566319 995785 566385 995788
rect 573135 995785 573201 995788
rect 634095 995785 634161 995788
rect 635823 995700 635889 995703
rect 551682 995698 635889 995700
rect 551682 995642 635828 995698
rect 635884 995642 635889 995698
rect 551682 995640 635889 995642
rect 544239 995637 544305 995640
rect 635823 995637 635889 995640
rect 521487 995550 529278 995552
rect 521487 995494 521492 995550
rect 521548 995494 529278 995550
rect 521487 995492 529278 995494
rect 521487 995489 521553 995492
rect 526095 995404 526161 995407
rect 510498 995402 526161 995404
rect 510498 995346 526100 995402
rect 526156 995346 526161 995402
rect 510498 995344 526161 995346
rect 526095 995341 526161 995344
rect 526479 995404 526545 995407
rect 530703 995404 530769 995407
rect 536847 995404 536913 995407
rect 561615 995404 561681 995407
rect 526479 995402 536913 995404
rect 526479 995346 526484 995402
rect 526540 995346 530708 995402
rect 530764 995346 536852 995402
rect 536908 995346 536913 995402
rect 526479 995344 536913 995346
rect 526479 995341 526545 995344
rect 530703 995341 530769 995344
rect 536847 995341 536913 995344
rect 550146 995402 561681 995404
rect 550146 995346 561620 995402
rect 561676 995346 561681 995402
rect 550146 995344 561681 995346
rect 469506 995196 499710 995256
rect 506562 995254 506673 995259
rect 506562 995198 506612 995254
rect 506668 995198 506673 995254
rect 506562 995196 506673 995198
rect 362799 995193 362865 995196
rect 368463 995193 368529 995196
rect 386319 995193 386385 995196
rect 443535 995193 443601 995196
rect 362799 995108 362865 995111
rect 342786 995106 362865 995108
rect 342786 995050 362804 995106
rect 362860 995050 362865 995106
rect 342786 995048 362865 995050
rect 362799 995045 362865 995048
rect 383247 995108 383313 995111
rect 393039 995108 393105 995111
rect 383247 995106 393105 995108
rect 383247 995050 383252 995106
rect 383308 995050 393044 995106
rect 393100 995050 393105 995106
rect 383247 995048 393105 995050
rect 499650 995108 499710 995196
rect 506607 995193 506673 995196
rect 521679 995256 521745 995259
rect 537135 995256 537201 995259
rect 521679 995254 537201 995256
rect 521679 995198 521684 995254
rect 521740 995198 537140 995254
rect 537196 995198 537201 995254
rect 521679 995196 537201 995198
rect 521679 995193 521745 995196
rect 537135 995193 537201 995196
rect 509679 995108 509745 995111
rect 550146 995108 550206 995344
rect 561615 995341 561681 995344
rect 581679 995404 581745 995407
rect 581679 995402 584766 995404
rect 581679 995346 581684 995402
rect 581740 995346 584766 995402
rect 581679 995344 584766 995346
rect 581679 995341 581745 995344
rect 584706 995259 584766 995344
rect 584706 995254 584817 995259
rect 584706 995198 584756 995254
rect 584812 995198 584817 995254
rect 584706 995196 584817 995198
rect 584751 995193 584817 995196
rect 604719 995256 604785 995259
rect 604719 995254 630270 995256
rect 604719 995198 604724 995254
rect 604780 995198 630270 995254
rect 604719 995196 630270 995198
rect 604719 995193 604785 995196
rect 499650 995106 509745 995108
rect 499650 995050 509684 995106
rect 509740 995050 509745 995106
rect 499650 995048 509745 995050
rect 383247 995045 383313 995048
rect 393039 995045 393105 995048
rect 509679 995045 509745 995048
rect 549954 995048 550206 995108
rect 570447 995108 570513 995111
rect 629967 995108 630033 995111
rect 570447 995106 630033 995108
rect 570447 995050 570452 995106
rect 570508 995050 629972 995106
rect 630028 995050 630033 995106
rect 570447 995048 630033 995050
rect 630210 995108 630270 995196
rect 641103 995108 641169 995111
rect 630210 995106 641169 995108
rect 630210 995050 641108 995106
rect 641164 995050 641169 995106
rect 630210 995048 641169 995050
rect 339759 994960 339825 994963
rect 319650 994958 339825 994960
rect 319650 994902 339764 994958
rect 339820 994902 339825 994958
rect 319650 994900 339825 994902
rect 339759 994897 339825 994900
rect 519279 994960 519345 994963
rect 526479 994960 526545 994963
rect 549954 994960 550014 995048
rect 570447 995045 570513 995048
rect 629967 995045 630033 995048
rect 641103 995045 641169 995048
rect 519279 994958 526545 994960
rect 519279 994902 519284 994958
rect 519340 994902 526484 994958
rect 526540 994902 526545 994958
rect 519279 994900 526545 994902
rect 519279 994897 519345 994900
rect 526479 994897 526545 994900
rect 539970 994900 550014 994960
rect 575439 994960 575505 994963
rect 630927 994960 630993 994963
rect 575439 994958 630993 994960
rect 575439 994902 575444 994958
rect 575500 994902 630932 994958
rect 630988 994902 630993 994958
rect 575439 994900 630993 994902
rect 262191 994810 296718 994812
rect 262191 994754 262196 994810
rect 262252 994754 296718 994810
rect 262191 994752 296718 994754
rect 368463 994812 368529 994815
rect 399855 994812 399921 994815
rect 368463 994810 399921 994812
rect 368463 994754 368468 994810
rect 368524 994754 399860 994810
rect 399916 994754 399921 994810
rect 368463 994752 399921 994754
rect 262191 994749 262257 994752
rect 368463 994749 368529 994752
rect 399855 994749 399921 994752
rect 509871 994812 509937 994815
rect 539970 994812 540030 994900
rect 575439 994897 575505 994900
rect 630927 994897 630993 994900
rect 509871 994810 540030 994812
rect 509871 994754 509876 994810
rect 509932 994754 540030 994810
rect 509871 994752 540030 994754
rect 572847 994812 572913 994815
rect 631791 994812 631857 994815
rect 572847 994810 631857 994812
rect 572847 994754 572852 994810
rect 572908 994754 631796 994810
rect 631852 994754 631857 994810
rect 572847 994752 631857 994754
rect 509871 994749 509937 994752
rect 572847 994749 572913 994752
rect 631791 994749 631857 994752
rect 242319 994664 242385 994667
rect 250479 994664 250545 994667
rect 242319 994662 250545 994664
rect 242319 994606 242324 994662
rect 242380 994606 250484 994662
rect 250540 994606 250545 994662
rect 242319 994604 250545 994606
rect 242319 994601 242385 994604
rect 250479 994601 250545 994604
rect 575343 994664 575409 994667
rect 637359 994664 637425 994667
rect 575343 994662 637425 994664
rect 575343 994606 575348 994662
rect 575404 994606 637364 994662
rect 637420 994606 637425 994662
rect 575343 994604 637425 994606
rect 575343 994601 575409 994604
rect 637359 994601 637425 994604
rect 638511 994664 638577 994667
rect 649839 994664 649905 994667
rect 638511 994662 649905 994664
rect 638511 994606 638516 994662
rect 638572 994606 649844 994662
rect 649900 994606 649905 994662
rect 638511 994604 649905 994606
rect 638511 994601 638577 994604
rect 649839 994601 649905 994604
rect 235791 994516 235857 994519
rect 247599 994516 247665 994519
rect 235791 994514 247665 994516
rect 235791 994458 235796 994514
rect 235852 994458 247604 994514
rect 247660 994458 247665 994514
rect 235791 994456 247665 994458
rect 235791 994453 235857 994456
rect 247599 994453 247665 994456
rect 572943 994516 573009 994519
rect 639183 994516 639249 994519
rect 572943 994514 639249 994516
rect 572943 994458 572948 994514
rect 573004 994458 639188 994514
rect 639244 994458 639249 994514
rect 572943 994456 639249 994458
rect 572943 994453 573009 994456
rect 639183 994453 639249 994456
rect 232143 994368 232209 994371
rect 242319 994368 242385 994371
rect 232143 994366 242385 994368
rect 232143 994310 232148 994366
rect 232204 994310 242324 994366
rect 242380 994310 242385 994366
rect 232143 994308 242385 994310
rect 232143 994305 232209 994308
rect 242319 994305 242385 994308
rect 242511 994368 242577 994371
rect 244815 994368 244881 994371
rect 242511 994366 244881 994368
rect 242511 994310 242516 994366
rect 242572 994310 244820 994366
rect 244876 994310 244881 994366
rect 242511 994308 244881 994310
rect 242511 994305 242577 994308
rect 244815 994305 244881 994308
rect 561423 994368 561489 994371
rect 634863 994368 634929 994371
rect 561423 994366 634929 994368
rect 561423 994310 561428 994366
rect 561484 994310 634868 994366
rect 634924 994310 634929 994366
rect 561423 994308 634929 994310
rect 561423 994305 561489 994308
rect 634863 994305 634929 994308
rect 182991 994220 183057 994223
rect 210255 994220 210321 994223
rect 182991 994218 210321 994220
rect 182991 994162 182996 994218
rect 183052 994162 210260 994218
rect 210316 994162 210321 994218
rect 182991 994160 210321 994162
rect 182991 994157 183057 994160
rect 210255 994157 210321 994160
rect 234351 994220 234417 994223
rect 254703 994220 254769 994223
rect 234351 994218 254769 994220
rect 234351 994162 234356 994218
rect 234412 994162 254708 994218
rect 254764 994162 254769 994218
rect 234351 994160 254769 994162
rect 234351 994157 234417 994160
rect 254703 994157 254769 994160
rect 296655 994220 296721 994223
rect 390831 994220 390897 994223
rect 479823 994220 479889 994223
rect 296655 994218 479889 994220
rect 296655 994162 296660 994218
rect 296716 994162 390836 994218
rect 390892 994162 479828 994218
rect 479884 994162 479889 994218
rect 296655 994160 479889 994162
rect 296655 994157 296721 994160
rect 390831 994157 390897 994160
rect 479823 994157 479889 994160
rect 536847 994220 536913 994223
rect 632367 994220 632433 994223
rect 536847 994218 632433 994220
rect 536847 994162 536852 994218
rect 536908 994162 632372 994218
rect 632428 994162 632433 994218
rect 536847 994160 632433 994162
rect 536847 994157 536913 994160
rect 632367 994157 632433 994160
rect 185391 994072 185457 994075
rect 236751 994072 236817 994075
rect 242511 994072 242577 994075
rect 185391 994070 242577 994072
rect 185391 994014 185396 994070
rect 185452 994014 236756 994070
rect 236812 994014 242516 994070
rect 242572 994014 242577 994070
rect 185391 994012 242577 994014
rect 185391 994009 185457 994012
rect 236751 994009 236817 994012
rect 242511 994009 242577 994012
rect 243183 994072 243249 994075
rect 640911 994072 640977 994075
rect 243183 994070 640977 994072
rect 243183 994014 243188 994070
rect 243244 994014 640916 994070
rect 640972 994014 640977 994070
rect 243183 994012 640977 994014
rect 243183 994009 243249 994012
rect 640911 994009 640977 994012
rect 84495 993922 106782 993924
rect 84495 993866 84500 993922
rect 84556 993866 106782 993922
rect 84495 993864 106782 993866
rect 129711 993924 129777 993927
rect 158991 993924 159057 993927
rect 129711 993922 159057 993924
rect 129711 993866 129716 993922
rect 129772 993866 158996 993922
rect 159052 993866 159057 993922
rect 129711 993864 159057 993866
rect 84495 993861 84561 993864
rect 129711 993861 129777 993864
rect 158991 993861 159057 993864
rect 191535 993924 191601 993927
rect 640527 993924 640593 993927
rect 191535 993922 640593 993924
rect 191535 993866 191540 993922
rect 191596 993866 640532 993922
rect 640588 993866 640593 993922
rect 191535 993864 640593 993866
rect 191535 993861 191601 993864
rect 640527 993861 640593 993864
rect 80175 993776 80241 993779
rect 106479 993776 106545 993779
rect 80175 993774 106545 993776
rect 80175 993718 80180 993774
rect 80236 993718 106484 993774
rect 106540 993718 106545 993774
rect 80175 993716 106545 993718
rect 80175 993713 80241 993716
rect 106479 993713 106545 993716
rect 83439 993630 83505 993631
rect 83386 993628 83392 993630
rect 83312 993568 83392 993628
rect 83456 993628 83505 993630
rect 92847 993628 92913 993631
rect 83456 993626 92913 993628
rect 83500 993570 92852 993626
rect 92908 993570 92913 993626
rect 83386 993566 83392 993568
rect 83456 993568 92913 993570
rect 83456 993566 83505 993568
rect 83439 993565 83505 993566
rect 92847 993565 92913 993568
rect 62031 992148 62097 992151
rect 83386 992148 83392 992150
rect 62031 992146 83392 992148
rect 62031 992090 62036 992146
rect 62092 992090 83392 992146
rect 62031 992088 83392 992090
rect 62031 992085 62097 992088
rect 83386 992086 83392 992088
rect 83456 992086 83462 992150
rect 655119 976756 655185 976759
rect 650208 976754 655185 976756
rect 650208 976698 655124 976754
rect 655180 976698 655185 976754
rect 650208 976696 655185 976698
rect 655119 976693 655185 976696
rect 59439 975424 59505 975427
rect 59439 975422 64416 975424
rect 59439 975366 59444 975422
rect 59500 975366 64416 975422
rect 59439 975364 64416 975366
rect 59439 975361 59505 975364
rect 40954 968702 40960 968766
rect 41024 968764 41030 968766
rect 41775 968764 41841 968767
rect 41024 968762 41841 968764
rect 41024 968706 41780 968762
rect 41836 968706 41841 968762
rect 41024 968704 41841 968706
rect 41024 968702 41030 968704
rect 41775 968701 41841 968704
rect 674319 967580 674385 967583
rect 674991 967580 675057 967583
rect 674319 967578 675057 967580
rect 674319 967522 674324 967578
rect 674380 967522 674996 967578
rect 675052 967522 675057 967578
rect 674319 967520 675057 967522
rect 674319 967517 674385 967520
rect 674991 967517 675057 967520
rect 674511 967432 674577 967435
rect 675322 967432 675328 967434
rect 674511 967430 675328 967432
rect 674511 967374 674516 967430
rect 674572 967374 675328 967430
rect 674511 967372 675328 967374
rect 674511 967369 674577 967372
rect 675322 967370 675328 967372
rect 675392 967370 675398 967434
rect 40570 967074 40576 967138
rect 40640 967136 40646 967138
rect 41775 967136 41841 967139
rect 40640 967134 41841 967136
rect 40640 967078 41780 967134
rect 41836 967078 41841 967134
rect 40640 967076 41841 967078
rect 40640 967074 40646 967076
rect 41775 967073 41841 967076
rect 675759 966396 675825 966399
rect 676666 966396 676672 966398
rect 675759 966394 676672 966396
rect 675759 966338 675764 966394
rect 675820 966338 676672 966394
rect 675759 966336 676672 966338
rect 675759 966333 675825 966336
rect 676666 966334 676672 966336
rect 676736 966334 676742 966398
rect 675663 965806 675729 965807
rect 675663 965802 675712 965806
rect 675776 965804 675782 965806
rect 675663 965746 675668 965802
rect 675663 965742 675712 965746
rect 675776 965744 675820 965804
rect 675776 965742 675782 965744
rect 675663 965741 675729 965742
rect 40762 965002 40768 965066
rect 40832 965064 40838 965066
rect 41775 965064 41841 965067
rect 655215 965064 655281 965067
rect 40832 965062 41841 965064
rect 40832 965006 41780 965062
rect 41836 965006 41841 965062
rect 40832 965004 41841 965006
rect 650208 965062 655281 965064
rect 650208 965006 655220 965062
rect 655276 965006 655281 965062
rect 650208 965004 655281 965006
rect 40832 965002 40838 965004
rect 41775 965001 41841 965004
rect 655215 965001 655281 965004
rect 675183 964918 675249 964919
rect 675130 964916 675136 964918
rect 675092 964856 675136 964916
rect 675200 964914 675249 964918
rect 675244 964858 675249 964914
rect 675130 964854 675136 964856
rect 675200 964854 675249 964858
rect 675183 964853 675249 964854
rect 40378 963966 40384 964030
rect 40448 964028 40454 964030
rect 41775 964028 41841 964031
rect 40448 964026 41841 964028
rect 40448 963970 41780 964026
rect 41836 963970 41841 964026
rect 40448 963968 41841 963970
rect 40448 963966 40454 963968
rect 41775 963965 41841 963968
rect 41530 963226 41536 963290
rect 41600 963288 41606 963290
rect 41775 963288 41841 963291
rect 41600 963286 41841 963288
rect 41600 963230 41780 963286
rect 41836 963230 41841 963286
rect 41600 963228 41841 963230
rect 41600 963226 41606 963228
rect 41775 963225 41841 963228
rect 675759 963288 675825 963291
rect 676474 963288 676480 963290
rect 675759 963286 676480 963288
rect 675759 963230 675764 963286
rect 675820 963230 676480 963286
rect 675759 963228 676480 963230
rect 675759 963225 675825 963228
rect 676474 963226 676480 963228
rect 676544 963226 676550 963290
rect 42159 962844 42225 962847
rect 42298 962844 42304 962846
rect 42159 962842 42304 962844
rect 42159 962786 42164 962842
rect 42220 962786 42304 962842
rect 42159 962784 42304 962786
rect 42159 962781 42225 962784
rect 42298 962782 42304 962784
rect 42368 962782 42374 962846
rect 674362 962486 674368 962550
rect 674432 962548 674438 962550
rect 675087 962548 675153 962551
rect 674432 962546 675153 962548
rect 674432 962490 675092 962546
rect 675148 962490 675153 962546
rect 674432 962488 675153 962490
rect 674432 962486 674438 962488
rect 675087 962485 675153 962488
rect 42063 962254 42129 962255
rect 42063 962250 42112 962254
rect 42176 962252 42182 962254
rect 43066 962252 43072 962254
rect 42063 962194 42068 962250
rect 42063 962190 42112 962194
rect 42176 962192 42220 962252
rect 42306 962192 43072 962252
rect 42176 962190 42182 962192
rect 42063 962189 42129 962190
rect 42159 962104 42225 962107
rect 42306 962104 42366 962192
rect 43066 962190 43072 962192
rect 43136 962252 43142 962254
rect 62031 962252 62097 962255
rect 43136 962250 62097 962252
rect 43136 962194 62036 962250
rect 62092 962194 62097 962250
rect 43136 962192 62097 962194
rect 43136 962190 43142 962192
rect 62031 962189 62097 962192
rect 674554 962190 674560 962254
rect 674624 962252 674630 962254
rect 675087 962252 675153 962255
rect 674624 962250 675153 962252
rect 674624 962194 675092 962250
rect 675148 962194 675153 962250
rect 674624 962192 675153 962194
rect 674624 962190 674630 962192
rect 675087 962189 675153 962192
rect 42159 962102 42366 962104
rect 42159 962046 42164 962102
rect 42220 962046 42366 962102
rect 42159 962044 42366 962046
rect 42447 962104 42513 962107
rect 42874 962104 42880 962106
rect 42447 962102 42880 962104
rect 42447 962046 42452 962102
rect 42508 962046 42880 962102
rect 42447 962044 42880 962046
rect 42159 962041 42225 962044
rect 42447 962041 42513 962044
rect 42874 962042 42880 962044
rect 42944 962104 42950 962106
rect 61839 962104 61905 962107
rect 42944 962102 61905 962104
rect 42944 962046 61844 962102
rect 61900 962046 61905 962102
rect 42944 962044 61905 962046
rect 42944 962042 42950 962044
rect 61839 962041 61905 962044
rect 674170 961450 674176 961514
rect 674240 961512 674246 961514
rect 675375 961512 675441 961515
rect 674240 961510 675441 961512
rect 674240 961454 675380 961510
rect 675436 961454 675441 961510
rect 674240 961452 675441 961454
rect 674240 961450 674246 961452
rect 675375 961449 675441 961452
rect 675375 961366 675441 961367
rect 675322 961302 675328 961366
rect 675392 961364 675441 961366
rect 675392 961362 675484 961364
rect 675436 961306 675484 961362
rect 675392 961304 675484 961306
rect 675392 961302 675441 961304
rect 675375 961301 675441 961302
rect 59535 960920 59601 960923
rect 59535 960918 64416 960920
rect 59535 960862 59540 960918
rect 59596 960862 64416 960918
rect 59535 960860 64416 960862
rect 59535 960857 59601 960860
rect 675471 960182 675537 960183
rect 675471 960180 675520 960182
rect 675428 960178 675520 960180
rect 675428 960122 675476 960178
rect 675428 960120 675520 960122
rect 675471 960118 675520 960120
rect 675584 960118 675590 960182
rect 675471 960117 675537 960118
rect 42159 959588 42225 959591
rect 42682 959588 42688 959590
rect 42159 959586 42688 959588
rect 42159 959530 42164 959586
rect 42220 959530 42688 959586
rect 42159 959528 42688 959530
rect 42159 959525 42225 959528
rect 42682 959526 42688 959528
rect 42752 959526 42758 959590
rect 41775 959146 41841 959147
rect 41722 959144 41728 959146
rect 41684 959084 41728 959144
rect 41792 959142 41841 959146
rect 41836 959086 41841 959142
rect 41722 959082 41728 959084
rect 41792 959082 41841 959086
rect 41775 959081 41841 959082
rect 675759 959144 675825 959147
rect 676090 959144 676096 959146
rect 675759 959142 676096 959144
rect 675759 959086 675764 959142
rect 675820 959086 676096 959142
rect 675759 959084 676096 959086
rect 675759 959081 675825 959084
rect 676090 959082 676096 959084
rect 676160 959082 676166 959146
rect 41967 958406 42033 958407
rect 41914 958404 41920 958406
rect 41876 958344 41920 958404
rect 41984 958402 42033 958406
rect 42028 958346 42033 958402
rect 41914 958342 41920 958344
rect 41984 958342 42033 958346
rect 41967 958341 42033 958342
rect 42159 957812 42225 957815
rect 42490 957812 42496 957814
rect 42159 957810 42496 957812
rect 42159 957754 42164 957810
rect 42220 957754 42496 957810
rect 42159 957752 42496 957754
rect 42159 957749 42225 957752
rect 42490 957750 42496 957752
rect 42560 957750 42566 957814
rect 674746 957750 674752 957814
rect 674816 957812 674822 957814
rect 675375 957812 675441 957815
rect 674816 957810 675441 957812
rect 674816 957754 675380 957810
rect 675436 957754 675441 957810
rect 674816 957752 675441 957754
rect 674816 957750 674822 957752
rect 675375 957749 675441 957752
rect 41146 956566 41152 956630
rect 41216 956628 41222 956630
rect 41775 956628 41841 956631
rect 41216 956626 41841 956628
rect 41216 956570 41780 956626
rect 41836 956570 41841 956626
rect 41216 956568 41841 956570
rect 41216 956566 41222 956568
rect 41775 956565 41841 956568
rect 674938 955974 674944 956038
rect 675008 956036 675014 956038
rect 675471 956036 675537 956039
rect 675008 956034 675537 956036
rect 675008 955978 675476 956034
rect 675532 955978 675537 956034
rect 675008 955976 675537 955978
rect 675008 955974 675014 955976
rect 675471 955973 675537 955976
rect 675087 953520 675153 953523
rect 677050 953520 677056 953522
rect 675087 953518 677056 953520
rect 675087 953462 675092 953518
rect 675148 953462 677056 953518
rect 675087 953460 677056 953462
rect 675087 953457 675153 953460
rect 677050 953458 677056 953460
rect 677120 953458 677126 953522
rect 654447 953372 654513 953375
rect 650208 953370 654513 953372
rect 650208 953314 654452 953370
rect 654508 953314 654513 953370
rect 650208 953312 654513 953314
rect 654447 953309 654513 953312
rect 675183 953372 675249 953375
rect 676858 953372 676864 953374
rect 675183 953370 676864 953372
rect 675183 953314 675188 953370
rect 675244 953314 676864 953370
rect 675183 953312 676864 953314
rect 675183 953309 675249 953312
rect 676858 953310 676864 953312
rect 676928 953310 676934 953374
rect 42306 949376 42366 949494
rect 42447 949376 42513 949379
rect 42306 949374 42513 949376
rect 42306 949318 42452 949374
rect 42508 949318 42513 949374
rect 42306 949316 42513 949318
rect 42447 949313 42513 949316
rect 42306 948491 42366 948680
rect 42306 948486 42417 948491
rect 42306 948430 42356 948486
rect 42412 948430 42417 948486
rect 42306 948428 42417 948430
rect 42351 948425 42417 948428
rect 42639 947896 42705 947899
rect 42336 947894 42705 947896
rect 42336 947838 42644 947894
rect 42700 947838 42705 947894
rect 42336 947836 42705 947838
rect 42639 947833 42705 947836
rect 40578 946567 40638 947052
rect 57807 946712 57873 946715
rect 57807 946710 64416 946712
rect 57807 946654 57812 946710
rect 57868 946654 64416 946710
rect 57807 946652 64416 946654
rect 57807 946649 57873 946652
rect 40578 946562 40689 946567
rect 40578 946506 40628 946562
rect 40684 946506 40689 946562
rect 40578 946504 40689 946506
rect 40623 946501 40689 946504
rect 47439 946268 47505 946271
rect 42336 946266 47505 946268
rect 42336 946210 47444 946266
rect 47500 946210 47505 946266
rect 42336 946208 47505 946210
rect 47439 946205 47505 946208
rect 47727 946120 47793 946123
rect 42306 946118 47793 946120
rect 42306 946062 47732 946118
rect 47788 946062 47793 946118
rect 42306 946060 47793 946062
rect 40239 945084 40305 945087
rect 42306 945084 42366 946060
rect 47727 946057 47793 946060
rect 674511 945380 674577 945383
rect 674754 945380 674814 945942
rect 674511 945378 674814 945380
rect 674511 945322 674516 945378
rect 674572 945322 674814 945378
rect 674511 945320 674814 945322
rect 674511 945317 674577 945320
rect 40239 945082 42366 945084
rect 40239 945026 40244 945082
rect 40300 945026 42366 945082
rect 40239 945024 42366 945026
rect 40239 945021 40305 945024
rect 40431 944936 40497 944939
rect 40431 944934 42366 944936
rect 40431 944878 40436 944934
rect 40492 944878 42366 944934
rect 40431 944876 42366 944878
rect 40431 944873 40497 944876
rect 42306 944788 42366 944876
rect 47919 944788 47985 944791
rect 42306 944786 47985 944788
rect 42306 944758 47924 944786
rect 42336 944730 47924 944758
rect 47980 944730 47985 944786
rect 42336 944728 47985 944730
rect 47919 944725 47985 944728
rect 674511 944788 674577 944791
rect 674754 944788 674814 945054
rect 674511 944786 674814 944788
rect 674511 944730 674516 944786
rect 674572 944730 674814 944786
rect 674511 944728 674814 944730
rect 674511 944725 674577 944728
rect 41146 944430 41152 944494
rect 41216 944430 41222 944494
rect 41154 943944 41214 944430
rect 674946 944051 675006 944240
rect 674895 944046 675006 944051
rect 674895 943990 674900 944046
rect 674956 943990 675006 944046
rect 674895 943988 675006 943990
rect 674895 943985 674961 943988
rect 40570 943690 40576 943754
rect 40640 943690 40646 943754
rect 40578 943130 40638 943690
rect 37359 942864 37425 942867
rect 37314 942862 37425 942864
rect 37314 942806 37364 942862
rect 37420 942806 37425 942862
rect 37314 942801 37425 942806
rect 674511 942864 674577 942867
rect 674754 942864 674814 943426
rect 674511 942862 674814 942864
rect 674511 942806 674516 942862
rect 674572 942806 674814 942862
rect 674511 942804 674814 942806
rect 674511 942801 674577 942804
rect 37314 942242 37374 942801
rect 673839 942568 673905 942571
rect 674754 942568 674814 942612
rect 673839 942566 674814 942568
rect 673839 942510 673844 942566
rect 673900 942510 674814 942566
rect 673839 942508 674814 942510
rect 673839 942505 673905 942508
rect 674415 941976 674481 941979
rect 674415 941974 674784 941976
rect 674415 941918 674420 941974
rect 674476 941918 674784 941974
rect 674415 941916 674784 941918
rect 674415 941913 674481 941916
rect 649551 941828 649617 941831
rect 649551 941826 649662 941828
rect 649551 941770 649556 941826
rect 649612 941770 649662 941826
rect 649551 941765 649662 941770
rect 42490 941680 42496 941682
rect 42306 941620 42496 941680
rect 42306 941502 42366 941620
rect 42490 941618 42496 941620
rect 42560 941618 42566 941682
rect 649602 941502 649662 941765
rect 42106 941174 42112 941238
rect 42176 941174 42182 941238
rect 42114 940762 42174 941174
rect 674415 941162 674481 941165
rect 674415 941160 674784 941162
rect 674415 941104 674420 941160
rect 674476 941104 674784 941160
rect 674415 941102 674784 941104
rect 674415 941099 674481 941102
rect 675130 940878 675136 940942
rect 675200 940878 675206 940942
rect 40954 940582 40960 940646
rect 41024 940582 41030 940646
rect 40962 940022 41022 940582
rect 675138 940318 675198 940878
rect 673935 939608 674001 939611
rect 673935 939606 674814 939608
rect 673935 939550 673940 939606
rect 673996 939550 674814 939606
rect 673935 939548 674814 939550
rect 673935 939545 674001 939548
rect 674754 939504 674814 939548
rect 676666 939250 676672 939314
rect 676736 939250 676742 939314
rect 42831 939164 42897 939167
rect 42336 939162 42897 939164
rect 42336 939106 42836 939162
rect 42892 939106 42897 939162
rect 42336 939104 42897 939106
rect 42831 939101 42897 939104
rect 41914 938806 41920 938870
rect 41984 938806 41990 938870
rect 41922 938394 41982 938806
rect 676674 938690 676734 939250
rect 41722 938066 41728 938130
rect 41792 938066 41798 938130
rect 676474 938066 676480 938130
rect 676544 938066 676550 938130
rect 41730 937506 41790 938066
rect 676482 937802 676542 938066
rect 40762 937326 40768 937390
rect 40832 937326 40838 937390
rect 676090 937326 676096 937390
rect 676160 937326 676166 937390
rect 40770 936766 40830 937326
rect 676098 937210 676158 937326
rect 676815 936648 676881 936651
rect 676815 936646 676926 936648
rect 676815 936590 676820 936646
rect 676876 936590 676926 936646
rect 676815 936585 676926 936590
rect 41530 936438 41536 936502
rect 41600 936438 41606 936502
rect 41538 936026 41598 936438
rect 676866 936322 676926 936585
rect 675706 935846 675712 935910
rect 675776 935846 675782 935910
rect 675714 935582 675774 935846
rect 42682 935316 42688 935318
rect 42336 935256 42688 935316
rect 42682 935254 42688 935256
rect 42752 935254 42758 935318
rect 42298 934958 42304 935022
rect 42368 934958 42374 935022
rect 42306 934398 42366 934958
rect 674362 934662 674368 934726
rect 674432 934724 674438 934726
rect 674432 934664 674784 934724
rect 674432 934662 674438 934664
rect 674554 934514 674560 934578
rect 674624 934576 674630 934578
rect 674624 934516 674814 934576
rect 674624 934514 674630 934516
rect 40378 934070 40384 934134
rect 40448 934070 40454 934134
rect 40386 933584 40446 934070
rect 674754 933954 674814 934516
rect 674938 933330 674944 933394
rect 675008 933330 675014 933394
rect 674946 933066 675006 933330
rect 674746 932886 674752 932950
rect 674816 932886 674822 932950
rect 42306 932507 42366 932770
rect 42306 932502 42417 932507
rect 42306 932446 42356 932502
rect 42412 932446 42417 932502
rect 674754 932474 674814 932886
rect 42306 932444 42417 932446
rect 42351 932441 42417 932444
rect 59535 932356 59601 932359
rect 59535 932354 64416 932356
rect 59535 932298 59540 932354
rect 59596 932298 64416 932354
rect 59535 932296 64416 932298
rect 59535 932293 59601 932296
rect 674170 931554 674176 931618
rect 674240 931616 674246 931618
rect 674240 931556 674784 931616
rect 674240 931554 674246 931556
rect 677050 931406 677056 931470
rect 677120 931406 677126 931470
rect 42306 931027 42366 931290
rect 42306 931022 42417 931027
rect 42306 930966 42356 931022
rect 42412 930966 42417 931022
rect 42306 930964 42417 930966
rect 42351 930961 42417 930964
rect 677058 930846 677118 931406
rect 676858 930222 676864 930286
rect 676928 930222 676934 930286
rect 676866 929958 676926 930222
rect 654447 929840 654513 929843
rect 650208 929838 654513 929840
rect 650208 929782 654452 929838
rect 654508 929782 654513 929838
rect 650208 929780 654513 929782
rect 654447 929777 654513 929780
rect 679746 928659 679806 929144
rect 679746 928654 679857 928659
rect 679746 928598 679796 928654
rect 679852 928598 679857 928654
rect 679746 928596 679857 928598
rect 679791 928593 679857 928596
rect 679791 928064 679857 928067
rect 679746 928062 679857 928064
rect 679746 928006 679796 928062
rect 679852 928006 679857 928062
rect 679746 928001 679857 928006
rect 679746 927664 679806 928001
rect 653967 918148 654033 918151
rect 650208 918146 654033 918148
rect 650208 918090 653972 918146
rect 654028 918090 654033 918146
rect 650208 918088 654033 918090
rect 653967 918085 654033 918088
rect 59535 917852 59601 917855
rect 59535 917850 64416 917852
rect 59535 917794 59540 917850
rect 59596 917794 64416 917850
rect 59535 917792 64416 917794
rect 59535 917789 59601 917792
rect 654447 906456 654513 906459
rect 650208 906454 654513 906456
rect 650208 906398 654452 906454
rect 654508 906398 654513 906454
rect 650208 906396 654513 906398
rect 654447 906393 654513 906396
rect 59535 903496 59601 903499
rect 59535 903494 64416 903496
rect 59535 903438 59540 903494
rect 59596 903438 64416 903494
rect 59535 903436 64416 903438
rect 59535 903433 59601 903436
rect 650031 895208 650097 895211
rect 649986 895206 650097 895208
rect 649986 895150 650036 895206
rect 650092 895150 650097 895206
rect 649986 895145 650097 895150
rect 649986 894586 650046 895145
rect 59535 889140 59601 889143
rect 59535 889138 64416 889140
rect 59535 889082 59540 889138
rect 59596 889082 64416 889138
rect 59535 889080 64416 889082
rect 59535 889077 59601 889080
rect 653967 882924 654033 882927
rect 650208 882922 654033 882924
rect 650208 882866 653972 882922
rect 654028 882866 654033 882922
rect 650208 882864 654033 882866
rect 653967 882861 654033 882864
rect 675759 877004 675825 877007
rect 676090 877004 676096 877006
rect 675759 877002 676096 877004
rect 675759 876946 675764 877002
rect 675820 876946 676096 877002
rect 675759 876944 676096 876946
rect 675759 876941 675825 876944
rect 676090 876942 676096 876944
rect 676160 876942 676166 877006
rect 673978 876498 673984 876562
rect 674048 876560 674054 876562
rect 675375 876560 675441 876563
rect 674048 876558 675441 876560
rect 674048 876502 675380 876558
rect 675436 876502 675441 876558
rect 674048 876500 675441 876502
rect 674048 876498 674054 876500
rect 675375 876497 675441 876500
rect 674746 875906 674752 875970
rect 674816 875968 674822 875970
rect 675375 875968 675441 875971
rect 674816 875966 675441 875968
rect 674816 875910 675380 875966
rect 675436 875910 675441 875966
rect 674816 875908 675441 875910
rect 674816 875906 674822 875908
rect 675375 875905 675441 875908
rect 675087 875820 675153 875823
rect 675322 875820 675328 875822
rect 675087 875818 675328 875820
rect 675087 875762 675092 875818
rect 675148 875762 675328 875818
rect 675087 875760 675328 875762
rect 675087 875757 675153 875760
rect 675322 875758 675328 875760
rect 675392 875758 675398 875822
rect 675183 875672 675249 875675
rect 675514 875672 675520 875674
rect 675183 875670 675520 875672
rect 675183 875614 675188 875670
rect 675244 875614 675520 875670
rect 675183 875612 675520 875614
rect 675183 875609 675249 875612
rect 675514 875610 675520 875612
rect 675584 875610 675590 875674
rect 59535 874784 59601 874787
rect 59535 874782 64416 874784
rect 59535 874726 59540 874782
rect 59596 874726 64416 874782
rect 59535 874724 64416 874726
rect 59535 874721 59601 874724
rect 674554 873982 674560 874046
rect 674624 874044 674630 874046
rect 675471 874044 675537 874047
rect 674624 874042 675537 874044
rect 674624 873986 675476 874042
rect 675532 873986 675537 874042
rect 674624 873984 675537 873986
rect 674624 873982 674630 873984
rect 675471 873981 675537 873984
rect 674170 873390 674176 873454
rect 674240 873452 674246 873454
rect 675375 873452 675441 873455
rect 674240 873450 675441 873452
rect 674240 873394 675380 873450
rect 675436 873394 675441 873450
rect 674240 873392 675441 873394
rect 674240 873390 674246 873392
rect 675375 873389 675441 873392
rect 654447 871232 654513 871235
rect 650208 871230 654513 871232
rect 650208 871174 654452 871230
rect 654508 871174 654513 871230
rect 650208 871172 654513 871174
rect 654447 871169 654513 871172
rect 674938 869838 674944 869902
rect 675008 869900 675014 869902
rect 675375 869900 675441 869903
rect 675008 869898 675441 869900
rect 675008 869842 675380 869898
rect 675436 869842 675441 869898
rect 675008 869840 675441 869842
rect 675008 869838 675014 869840
rect 675375 869837 675441 869840
rect 675759 864720 675825 864723
rect 676666 864720 676672 864722
rect 675759 864718 676672 864720
rect 675759 864662 675764 864718
rect 675820 864662 676672 864718
rect 675759 864660 676672 864662
rect 675759 864657 675825 864660
rect 676666 864658 676672 864660
rect 676736 864658 676742 864722
rect 675375 862946 675441 862947
rect 675322 862944 675328 862946
rect 675284 862884 675328 862944
rect 675392 862942 675441 862946
rect 675436 862886 675441 862942
rect 675322 862882 675328 862884
rect 675392 862882 675441 862886
rect 675375 862881 675441 862882
rect 58575 860428 58641 860431
rect 58575 860426 64416 860428
rect 58575 860370 58580 860426
rect 58636 860370 64416 860426
rect 58575 860368 64416 860370
rect 58575 860365 58641 860368
rect 654159 859540 654225 859543
rect 650208 859538 654225 859540
rect 650208 859482 654164 859538
rect 654220 859482 654225 859538
rect 650208 859480 654225 859482
rect 654159 859477 654225 859480
rect 650127 848292 650193 848295
rect 650127 848290 650238 848292
rect 650127 848234 650132 848290
rect 650188 848234 650238 848290
rect 650127 848229 650238 848234
rect 650178 847670 650238 848229
rect 59535 846072 59601 846075
rect 59535 846070 64416 846072
rect 59535 846014 59540 846070
rect 59596 846014 64416 846070
rect 59535 846012 64416 846014
rect 59535 846009 59601 846012
rect 653967 836008 654033 836011
rect 650208 836006 654033 836008
rect 650208 835950 653972 836006
rect 654028 835950 654033 836006
rect 650208 835948 654033 835950
rect 653967 835945 654033 835948
rect 59535 831716 59601 831719
rect 59535 831714 64416 831716
rect 59535 831658 59540 831714
rect 59596 831658 64416 831714
rect 59535 831656 64416 831658
rect 59535 831653 59601 831656
rect 653967 824316 654033 824319
rect 650208 824314 654033 824316
rect 650208 824258 653972 824314
rect 654028 824258 654033 824314
rect 650208 824256 654033 824258
rect 653967 824253 654033 824256
rect 42159 823872 42225 823875
rect 42114 823870 42225 823872
rect 42114 823814 42164 823870
rect 42220 823814 42225 823870
rect 42114 823809 42225 823814
rect 42114 823694 42174 823809
rect 42159 823132 42225 823135
rect 42114 823130 42225 823132
rect 42114 823074 42164 823130
rect 42220 823074 42225 823130
rect 42114 823069 42225 823074
rect 42114 822880 42174 823069
rect 42159 822244 42225 822247
rect 42114 822242 42225 822244
rect 42114 822186 42164 822242
rect 42220 822186 42225 822242
rect 42114 822181 42225 822186
rect 42114 822066 42174 822181
rect 43215 821208 43281 821211
rect 42336 821206 43281 821208
rect 42336 821150 43220 821206
rect 43276 821150 43281 821206
rect 42336 821148 43281 821150
rect 43215 821145 43281 821148
rect 40623 820764 40689 820767
rect 40578 820762 40689 820764
rect 40578 820706 40628 820762
rect 40684 820706 40689 820762
rect 40578 820701 40689 820706
rect 40578 820438 40638 820701
rect 40239 820024 40305 820027
rect 40194 820022 40305 820024
rect 40194 819966 40244 820022
rect 40300 819966 40305 820022
rect 40194 819961 40305 819966
rect 37263 819136 37329 819139
rect 40194 819136 40254 819961
rect 40431 819580 40497 819583
rect 37263 819134 40254 819136
rect 37263 819078 37268 819134
rect 37324 819078 40254 819134
rect 37263 819076 40254 819078
rect 40386 819578 40497 819580
rect 40386 819522 40436 819578
rect 40492 819522 40497 819578
rect 40386 819517 40497 819522
rect 37263 819073 37329 819076
rect 40386 818988 40446 819517
rect 40386 818958 41376 818988
rect 40416 818928 41406 818958
rect 41346 818694 41406 818928
rect 41338 818630 41344 818694
rect 41408 818630 41414 818694
rect 41730 817955 41790 818070
rect 41679 817950 41790 817955
rect 41679 817894 41684 817950
rect 41740 817894 41790 817950
rect 41679 817892 41790 817894
rect 41679 817889 41745 817892
rect 59535 817360 59601 817363
rect 59535 817358 64416 817360
rect 40194 816771 40254 817330
rect 59535 817302 59540 817358
rect 59596 817302 64416 817358
rect 59535 817300 64416 817302
rect 59535 817297 59601 817300
rect 40143 816766 40254 816771
rect 40143 816710 40148 816766
rect 40204 816710 40254 816766
rect 40143 816708 40254 816710
rect 40143 816705 40209 816708
rect 40194 815883 40254 816442
rect 40194 815878 40305 815883
rect 40194 815822 40244 815878
rect 40300 815822 40305 815878
rect 40194 815820 40305 815822
rect 40239 815817 40305 815820
rect 42831 815732 42897 815735
rect 42336 815730 42897 815732
rect 42336 815674 42836 815730
rect 42892 815674 42897 815730
rect 42336 815672 42897 815674
rect 42831 815669 42897 815672
rect 43023 814992 43089 814995
rect 42336 814990 43089 814992
rect 42336 814934 43028 814990
rect 43084 814934 43089 814990
rect 42336 814932 43089 814934
rect 43023 814929 43089 814932
rect 41922 813663 41982 814222
rect 41871 813658 41982 813663
rect 41871 813602 41876 813658
rect 41932 813602 41982 813658
rect 41871 813600 41982 813602
rect 41871 813597 41937 813600
rect 37314 812775 37374 813334
rect 37314 812770 37425 812775
rect 37314 812714 37364 812770
rect 37420 812714 37425 812770
rect 37314 812712 37425 812714
rect 37359 812709 37425 812712
rect 654447 812624 654513 812627
rect 650208 812622 654513 812624
rect 650208 812566 654452 812622
rect 654508 812566 654513 812622
rect 650208 812564 654513 812566
rect 654447 812561 654513 812564
rect 41922 812331 41982 812520
rect 41922 812326 42033 812331
rect 41922 812270 41972 812326
rect 42028 812270 42033 812326
rect 41922 812268 42033 812270
rect 41967 812265 42033 812268
rect 41538 811147 41598 811706
rect 41487 811142 41598 811147
rect 41487 811086 41492 811142
rect 41548 811086 41598 811142
rect 41487 811084 41598 811086
rect 41487 811081 41553 811084
rect 42306 810404 42366 810892
rect 43023 810404 43089 810407
rect 42306 810402 43089 810404
rect 42306 810346 43028 810402
rect 43084 810346 43089 810402
rect 42306 810344 43089 810346
rect 43023 810341 43089 810344
rect 41730 809667 41790 810226
rect 41730 809662 41841 809667
rect 41730 809606 41780 809662
rect 41836 809606 41841 809662
rect 41730 809604 41841 809606
rect 41775 809601 41841 809604
rect 41538 809223 41598 809412
rect 41538 809218 41649 809223
rect 41538 809162 41588 809218
rect 41644 809162 41649 809218
rect 41538 809160 41649 809162
rect 41583 809157 41649 809160
rect 42114 808335 42174 808598
rect 42063 808330 42174 808335
rect 42063 808274 42068 808330
rect 42124 808274 42174 808330
rect 42063 808272 42174 808274
rect 42063 808269 42129 808272
rect 42306 807740 42366 807784
rect 43119 807740 43185 807743
rect 42306 807738 43185 807740
rect 42306 807682 43124 807738
rect 43180 807682 43185 807738
rect 42306 807680 43185 807682
rect 43119 807677 43185 807680
rect 42831 807000 42897 807003
rect 42336 806998 42897 807000
rect 42336 806942 42836 806998
rect 42892 806942 42897 806998
rect 42336 806940 42897 806942
rect 42831 806937 42897 806940
rect 42831 805520 42897 805523
rect 42336 805518 42897 805520
rect 42336 805462 42836 805518
rect 42892 805462 42897 805518
rect 42336 805460 42897 805462
rect 42831 805457 42897 805460
rect 59535 802856 59601 802859
rect 59535 802854 64416 802856
rect 59535 802798 59540 802854
rect 59596 802798 64416 802854
rect 59535 802796 64416 802798
rect 59535 802793 59601 802796
rect 37359 802264 37425 802267
rect 41530 802264 41536 802266
rect 37359 802262 41536 802264
rect 37359 802206 37364 802262
rect 37420 802206 41536 802262
rect 37359 802204 41536 802206
rect 37359 802201 37425 802204
rect 41530 802202 41536 802204
rect 41600 802202 41606 802266
rect 42447 802264 42513 802267
rect 42682 802264 42688 802266
rect 42447 802262 42688 802264
rect 42447 802206 42452 802262
rect 42508 802206 42688 802262
rect 42447 802204 42688 802206
rect 42447 802201 42513 802204
rect 42682 802202 42688 802204
rect 42752 802202 42758 802266
rect 37263 802116 37329 802119
rect 41146 802116 41152 802118
rect 37263 802114 41152 802116
rect 37263 802058 37268 802114
rect 37324 802058 41152 802114
rect 37263 802056 41152 802058
rect 37263 802053 37329 802056
rect 41146 802054 41152 802056
rect 41216 802054 41222 802118
rect 40239 801968 40305 801971
rect 41722 801968 41728 801970
rect 40239 801966 41728 801968
rect 40239 801910 40244 801966
rect 40300 801910 41728 801966
rect 40239 801908 41728 801910
rect 40239 801905 40305 801908
rect 41722 801906 41728 801908
rect 41792 801906 41798 801970
rect 649647 801376 649713 801379
rect 649602 801374 649713 801376
rect 649602 801318 649652 801374
rect 649708 801318 649713 801374
rect 649602 801313 649713 801318
rect 649602 800754 649662 801313
rect 41679 800488 41745 800491
rect 42298 800488 42304 800490
rect 41679 800486 42304 800488
rect 41679 800430 41684 800486
rect 41740 800430 42304 800486
rect 41679 800428 42304 800430
rect 41679 800425 41745 800428
rect 42298 800426 42304 800428
rect 42368 800426 42374 800490
rect 41775 800340 41841 800343
rect 42063 800342 42129 800343
rect 41914 800340 41920 800342
rect 41775 800338 41920 800340
rect 41775 800282 41780 800338
rect 41836 800282 41920 800338
rect 41775 800280 41920 800282
rect 41775 800277 41841 800280
rect 41914 800278 41920 800280
rect 41984 800278 41990 800342
rect 42063 800338 42112 800342
rect 42176 800340 42182 800342
rect 42063 800282 42068 800338
rect 42063 800278 42112 800282
rect 42176 800280 42220 800340
rect 42176 800278 42182 800280
rect 42063 800277 42129 800278
rect 42447 799750 42513 799751
rect 42447 799748 42496 799750
rect 42404 799746 42496 799748
rect 42404 799690 42452 799746
rect 42404 799688 42496 799690
rect 42447 799686 42496 799688
rect 42560 799686 42566 799750
rect 42447 799685 42513 799686
rect 42682 798354 42688 798418
rect 42752 798416 42758 798418
rect 43023 798416 43089 798419
rect 42752 798414 43089 798416
rect 42752 798358 43028 798414
rect 43084 798358 43089 798414
rect 42752 798356 43089 798358
rect 42752 798354 42758 798356
rect 43023 798353 43089 798356
rect 41871 794274 41937 794275
rect 41871 794272 41920 794274
rect 41828 794270 41920 794272
rect 41828 794214 41876 794270
rect 41828 794212 41920 794214
rect 41871 794210 41920 794212
rect 41984 794210 41990 794274
rect 41871 794209 41937 794210
rect 42063 793830 42129 793831
rect 42063 793828 42112 793830
rect 42020 793826 42112 793828
rect 42020 793770 42068 793826
rect 42020 793768 42112 793770
rect 42063 793766 42112 793768
rect 42176 793766 42182 793830
rect 42063 793765 42129 793766
rect 42447 792498 42513 792499
rect 42447 792494 42496 792498
rect 42560 792496 42566 792498
rect 42447 792438 42452 792494
rect 42447 792434 42496 792438
rect 42560 792436 42604 792496
rect 42560 792434 42566 792436
rect 42447 792433 42513 792434
rect 42298 792286 42304 792350
rect 42368 792348 42374 792350
rect 43023 792348 43089 792351
rect 42368 792346 43089 792348
rect 42368 792290 43028 792346
rect 43084 792290 43089 792346
rect 42368 792288 43089 792290
rect 42368 792286 42374 792288
rect 43023 792285 43089 792288
rect 41530 791842 41536 791906
rect 41600 791904 41606 791906
rect 42831 791904 42897 791907
rect 41600 791902 42897 791904
rect 41600 791846 42836 791902
rect 42892 791846 42897 791902
rect 41600 791844 42897 791846
rect 41600 791842 41606 791844
rect 42831 791841 42897 791844
rect 42106 791694 42112 791758
rect 42176 791756 42182 791758
rect 42927 791756 42993 791759
rect 42176 791754 42993 791756
rect 42176 791698 42932 791754
rect 42988 791698 42993 791754
rect 42176 791696 42993 791698
rect 42176 791694 42182 791696
rect 42927 791693 42993 791696
rect 42063 791166 42129 791167
rect 42063 791164 42112 791166
rect 42020 791162 42112 791164
rect 42176 791164 42182 791166
rect 43066 791164 43072 791166
rect 42020 791106 42068 791162
rect 42020 791104 42112 791106
rect 42063 791102 42112 791104
rect 42176 791104 43072 791164
rect 42176 791102 42182 791104
rect 43066 791102 43072 791104
rect 43136 791102 43142 791166
rect 42063 791101 42129 791102
rect 41530 790954 41536 791018
rect 41600 791016 41606 791018
rect 42159 791016 42225 791019
rect 42874 791016 42880 791018
rect 41600 791014 42880 791016
rect 41600 790958 42164 791014
rect 42220 790958 42880 791014
rect 41600 790956 42880 790958
rect 41600 790954 41606 790956
rect 42159 790953 42225 790956
rect 42874 790954 42880 790956
rect 42944 790954 42950 791018
rect 41722 790510 41728 790574
rect 41792 790572 41798 790574
rect 42735 790572 42801 790575
rect 41792 790570 42801 790572
rect 41792 790514 42740 790570
rect 42796 790514 42801 790570
rect 41792 790512 42801 790514
rect 41792 790510 41798 790512
rect 42735 790509 42801 790512
rect 654063 789092 654129 789095
rect 650208 789090 654129 789092
rect 650208 789034 654068 789090
rect 654124 789034 654129 789090
rect 650208 789032 654129 789034
rect 654063 789029 654129 789032
rect 42159 788648 42225 788651
rect 42298 788648 42304 788650
rect 42159 788646 42304 788648
rect 42159 788590 42164 788646
rect 42220 788590 42304 788646
rect 42159 788588 42304 788590
rect 42159 788585 42225 788588
rect 42298 788586 42304 788588
rect 42368 788586 42374 788650
rect 59535 788648 59601 788651
rect 59535 788646 64416 788648
rect 59535 788590 59540 788646
rect 59596 788590 64416 788646
rect 59535 788588 64416 788590
rect 59535 788585 59601 788588
rect 675663 788058 675729 788059
rect 675663 788054 675712 788058
rect 675776 788056 675782 788058
rect 675663 787998 675668 788054
rect 675663 787994 675712 787998
rect 675776 787996 675820 788056
rect 675776 787994 675782 787996
rect 675663 787993 675729 787994
rect 675471 787170 675537 787171
rect 675471 787166 675520 787170
rect 675584 787168 675590 787170
rect 675471 787110 675476 787166
rect 675471 787106 675520 787110
rect 675584 787108 675628 787168
rect 675584 787106 675590 787108
rect 675471 787105 675537 787106
rect 675759 786724 675825 786727
rect 676474 786724 676480 786726
rect 675759 786722 676480 786724
rect 675759 786666 675764 786722
rect 675820 786666 676480 786722
rect 675759 786664 676480 786666
rect 675759 786661 675825 786664
rect 676474 786662 676480 786664
rect 676544 786662 676550 786726
rect 675759 784800 675825 784803
rect 675898 784800 675904 784802
rect 675759 784798 675904 784800
rect 675759 784742 675764 784798
rect 675820 784742 675904 784798
rect 675759 784740 675904 784742
rect 675759 784737 675825 784740
rect 675898 784738 675904 784740
rect 675968 784738 675974 784802
rect 674362 780594 674368 780658
rect 674432 780656 674438 780658
rect 675471 780656 675537 780659
rect 674432 780654 675537 780656
rect 674432 780598 675476 780654
rect 675532 780598 675537 780654
rect 674432 780596 675537 780598
rect 674432 780594 674438 780596
rect 675471 780593 675537 780596
rect 42735 780508 42801 780511
rect 42336 780506 42801 780508
rect 42336 780450 42740 780506
rect 42796 780450 42801 780506
rect 42336 780448 42801 780450
rect 42735 780445 42801 780448
rect 42735 779694 42801 779697
rect 42336 779692 42801 779694
rect 42336 779636 42740 779692
rect 42796 779636 42801 779692
rect 42336 779634 42801 779636
rect 42735 779631 42801 779634
rect 675759 779176 675825 779179
rect 676858 779176 676864 779178
rect 675759 779174 676864 779176
rect 675759 779118 675764 779174
rect 675820 779118 676864 779174
rect 675759 779116 676864 779118
rect 675759 779113 675825 779116
rect 676858 779114 676864 779116
rect 676928 779114 676934 779178
rect 42735 778880 42801 778883
rect 42336 778878 42801 778880
rect 42336 778822 42740 778878
rect 42796 778822 42801 778878
rect 42336 778820 42801 778822
rect 42735 778817 42801 778820
rect 42306 777992 42366 778036
rect 43311 777992 43377 777995
rect 42306 777990 43377 777992
rect 42306 777934 43316 777990
rect 43372 777934 43377 777990
rect 42306 777932 43377 777934
rect 43311 777929 43377 777932
rect 674511 777548 674577 777551
rect 677050 777548 677056 777550
rect 674511 777546 677056 777548
rect 674511 777490 674516 777546
rect 674572 777490 677056 777546
rect 674511 777488 677056 777490
rect 674511 777485 674577 777488
rect 677050 777486 677056 777488
rect 677120 777486 677126 777550
rect 654063 777400 654129 777403
rect 650208 777398 654129 777400
rect 650208 777342 654068 777398
rect 654124 777342 654129 777398
rect 650208 777340 654129 777342
rect 654063 777337 654129 777340
rect 675759 777400 675825 777403
rect 677050 777400 677056 777402
rect 675759 777398 677056 777400
rect 675759 777342 675764 777398
rect 675820 777342 677056 777398
rect 675759 777340 677056 777342
rect 675759 777337 675825 777340
rect 677050 777338 677056 777340
rect 677120 777338 677126 777402
rect 43215 777252 43281 777255
rect 42336 777250 43281 777252
rect 42336 777194 43220 777250
rect 43276 777194 43281 777250
rect 42336 777192 43281 777194
rect 43215 777189 43281 777192
rect 41146 776746 41152 776810
rect 41216 776746 41222 776810
rect 41154 776512 41214 776746
rect 41154 776482 41568 776512
rect 41184 776452 41598 776482
rect 41538 775922 41598 776452
rect 41530 775858 41536 775922
rect 41600 775858 41606 775922
rect 41346 775182 41406 775742
rect 675759 775476 675825 775479
rect 676282 775476 676288 775478
rect 675759 775474 676288 775476
rect 675759 775418 675764 775474
rect 675820 775418 676288 775474
rect 675759 775416 676288 775418
rect 675759 775413 675825 775416
rect 676282 775414 676288 775416
rect 676352 775414 676358 775478
rect 41338 775118 41344 775182
rect 41408 775118 41414 775182
rect 42927 774884 42993 774887
rect 42336 774882 42993 774884
rect 42336 774826 42932 774882
rect 42988 774826 42993 774882
rect 42336 774824 42993 774826
rect 42927 774821 42993 774824
rect 59535 774144 59601 774147
rect 59535 774142 64416 774144
rect 39042 773555 39102 774114
rect 59535 774086 59540 774142
rect 59596 774086 64416 774142
rect 59535 774084 64416 774086
rect 59535 774081 59601 774084
rect 675130 773638 675136 773702
rect 675200 773700 675206 773702
rect 675471 773700 675537 773703
rect 675200 773698 675537 773700
rect 675200 773642 675476 773698
rect 675532 773642 675537 773698
rect 675200 773640 675537 773642
rect 675200 773638 675206 773640
rect 675471 773637 675537 773640
rect 38991 773550 39102 773555
rect 38991 773494 38996 773550
rect 39052 773494 39102 773550
rect 38991 773492 39102 773494
rect 38991 773489 39057 773492
rect 38850 772667 38910 773226
rect 674127 773108 674193 773111
rect 677818 773108 677824 773110
rect 674127 773106 677824 773108
rect 674127 773050 674132 773106
rect 674188 773050 677824 773106
rect 674127 773048 677824 773050
rect 674127 773045 674193 773048
rect 677818 773046 677824 773048
rect 677888 773046 677894 773110
rect 38799 772662 38910 772667
rect 38799 772606 38804 772662
rect 38860 772606 38910 772662
rect 38799 772604 38910 772606
rect 38799 772601 38865 772604
rect 43023 772516 43089 772519
rect 42336 772514 43089 772516
rect 42336 772458 43028 772514
rect 43084 772458 43089 772514
rect 42336 772456 43089 772458
rect 43023 772453 43089 772456
rect 41538 771187 41598 771746
rect 41487 771182 41598 771187
rect 41487 771126 41492 771182
rect 41548 771126 41598 771182
rect 41487 771124 41598 771126
rect 41487 771121 41553 771124
rect 41922 770447 41982 771006
rect 41871 770442 41982 770447
rect 41871 770386 41876 770442
rect 41932 770386 41982 770442
rect 41871 770384 41982 770386
rect 41871 770381 41937 770384
rect 37314 769559 37374 770118
rect 37314 769554 37425 769559
rect 37314 769498 37364 769554
rect 37420 769498 37425 769554
rect 37314 769496 37425 769498
rect 37359 769493 37425 769496
rect 41346 769115 41406 769378
rect 41346 769110 41457 769115
rect 41346 769054 41396 769110
rect 41452 769054 41457 769110
rect 41346 769052 41457 769054
rect 41391 769049 41457 769052
rect 41538 767931 41598 768490
rect 41538 767926 41649 767931
rect 41538 767870 41588 767926
rect 41644 767870 41649 767926
rect 41538 767868 41649 767870
rect 41583 767865 41649 767868
rect 42114 767339 42174 767750
rect 674415 767484 674481 767487
rect 674415 767482 674784 767484
rect 674415 767426 674420 767482
rect 674476 767426 674784 767482
rect 674415 767424 674784 767426
rect 674415 767421 674481 767424
rect 42063 767334 42174 767339
rect 42063 767278 42068 767334
rect 42124 767278 42174 767334
rect 42063 767276 42174 767278
rect 42063 767273 42129 767276
rect 41922 766451 41982 767010
rect 674607 766892 674673 766895
rect 674607 766890 674814 766892
rect 674607 766834 674612 766890
rect 674668 766834 674814 766890
rect 674607 766832 674814 766834
rect 674607 766829 674673 766832
rect 674754 766714 674814 766832
rect 41922 766446 42033 766451
rect 41922 766390 41972 766446
rect 42028 766390 42033 766446
rect 41922 766388 42033 766390
rect 41967 766385 42033 766388
rect 41730 766007 41790 766196
rect 41730 766002 41841 766007
rect 41730 765946 41780 766002
rect 41836 765946 41841 766002
rect 41730 765944 41841 765946
rect 41775 765941 41841 765944
rect 674415 765856 674481 765859
rect 674415 765854 674784 765856
rect 674415 765798 674420 765854
rect 674476 765798 674784 765854
rect 674415 765796 674784 765798
rect 674415 765793 674481 765796
rect 653967 765560 654033 765563
rect 650208 765558 654033 765560
rect 650208 765502 653972 765558
rect 654028 765502 654033 765558
rect 650208 765500 654033 765502
rect 653967 765497 654033 765500
rect 41730 765267 41790 765382
rect 41679 765262 41790 765267
rect 41679 765206 41684 765262
rect 41740 765206 41790 765262
rect 41679 765204 41790 765206
rect 41679 765201 41745 765204
rect 673839 765116 673905 765119
rect 673839 765114 674784 765116
rect 673839 765058 673844 765114
rect 673900 765058 674784 765114
rect 673839 765056 674784 765058
rect 673839 765053 673905 765056
rect 42306 764080 42366 764568
rect 673839 764228 673905 764231
rect 673839 764226 674784 764228
rect 673839 764170 673844 764226
rect 673900 764170 674784 764226
rect 673839 764168 674784 764170
rect 673839 764165 673905 764168
rect 42490 764080 42496 764082
rect 42306 764020 42496 764080
rect 42490 764018 42496 764020
rect 42560 764018 42566 764082
rect 42114 763491 42174 763754
rect 674415 763562 674481 763565
rect 674415 763560 674784 763562
rect 674415 763504 674420 763560
rect 674476 763504 674784 763560
rect 674415 763502 674784 763504
rect 674415 763499 674481 763502
rect 42114 763486 42225 763491
rect 42114 763430 42164 763486
rect 42220 763430 42225 763486
rect 42114 763428 42225 763430
rect 42159 763425 42225 763428
rect 673839 762748 673905 762751
rect 673839 762746 674784 762748
rect 673839 762690 673844 762746
rect 673900 762690 674784 762746
rect 673839 762688 674784 762690
rect 673839 762685 673905 762688
rect 674746 762390 674752 762454
rect 674816 762390 674822 762454
rect 42114 762011 42174 762274
rect 42114 762006 42225 762011
rect 42114 761950 42164 762006
rect 42220 761950 42225 762006
rect 42114 761948 42225 761950
rect 42159 761945 42225 761948
rect 674754 761904 674814 762390
rect 676666 761650 676672 761714
rect 676736 761650 676742 761714
rect 676674 761090 676734 761650
rect 42874 760466 42880 760530
rect 42944 760528 42950 760530
rect 43023 760528 43089 760531
rect 42944 760526 43089 760528
rect 42944 760470 43028 760526
rect 43084 760470 43089 760526
rect 42944 760468 43089 760470
rect 42944 760466 42950 760468
rect 43023 760465 43089 760468
rect 676090 760466 676096 760530
rect 676160 760466 676166 760530
rect 676098 760276 676158 760466
rect 38799 760232 38865 760235
rect 41146 760232 41152 760234
rect 38799 760230 41152 760232
rect 38799 760174 38804 760230
rect 38860 760174 41152 760230
rect 38799 760172 41152 760174
rect 38799 760169 38865 760172
rect 41146 760170 41152 760172
rect 41216 760170 41222 760234
rect 674554 760022 674560 760086
rect 674624 760084 674630 760086
rect 674624 760024 674814 760084
rect 674624 760022 674630 760024
rect 59535 759788 59601 759791
rect 59535 759786 64416 759788
rect 59535 759730 59540 759786
rect 59596 759730 64416 759786
rect 59535 759728 64416 759730
rect 59535 759725 59601 759728
rect 674754 759462 674814 760024
rect 674938 759134 674944 759198
rect 675008 759134 675014 759198
rect 37359 758752 37425 758755
rect 40762 758752 40768 758754
rect 37359 758750 40768 758752
rect 37359 758694 37364 758750
rect 37420 758694 40768 758750
rect 37359 758692 40768 758694
rect 37359 758689 37425 758692
rect 40762 758690 40768 758692
rect 40832 758690 40838 758754
rect 674946 758722 675006 759134
rect 675322 758542 675328 758606
rect 675392 758542 675398 758606
rect 41967 758456 42033 758459
rect 42682 758456 42688 758458
rect 41967 758454 42688 758456
rect 41967 758398 41972 758454
rect 42028 758398 42688 758454
rect 41967 758396 42688 758398
rect 41967 758393 42033 758396
rect 42682 758394 42688 758396
rect 42752 758394 42758 758458
rect 675330 757982 675390 758542
rect 41583 757420 41649 757423
rect 43066 757420 43072 757422
rect 41583 757418 43072 757420
rect 41583 757362 41588 757418
rect 41644 757362 43072 757418
rect 41583 757360 43072 757362
rect 41583 757357 41649 757360
rect 43066 757358 43072 757360
rect 43136 757358 43142 757422
rect 40954 757210 40960 757274
rect 41024 757272 41030 757274
rect 42106 757272 42112 757274
rect 41024 757212 42112 757272
rect 41024 757210 41030 757212
rect 42106 757210 42112 757212
rect 42176 757210 42182 757274
rect 41775 757126 41841 757127
rect 41722 757124 41728 757126
rect 41684 757064 41728 757124
rect 41792 757122 41841 757126
rect 41836 757066 41841 757122
rect 41722 757062 41728 757064
rect 41792 757062 41841 757066
rect 41775 757061 41841 757062
rect 42063 757126 42129 757127
rect 42063 757122 42112 757126
rect 42176 757124 42182 757126
rect 42063 757066 42068 757122
rect 42063 757062 42112 757066
rect 42176 757064 42220 757124
rect 42176 757062 42182 757064
rect 673978 757062 673984 757126
rect 674048 757124 674054 757126
rect 674048 757064 674784 757124
rect 674048 757062 674054 757064
rect 42063 757061 42129 757062
rect 674170 756322 674176 756386
rect 674240 756384 674246 756386
rect 674240 756324 674784 756384
rect 674240 756322 674246 756324
rect 673167 755496 673233 755499
rect 673167 755494 674784 755496
rect 673167 755438 673172 755494
rect 673228 755438 674784 755494
rect 673167 755436 674784 755438
rect 673167 755433 673233 755436
rect 677818 755286 677824 755350
rect 677888 755286 677894 755350
rect 677826 754726 677886 755286
rect 649935 754608 650001 754611
rect 649935 754606 650046 754608
rect 649935 754550 649940 754606
rect 649996 754550 650046 754606
rect 649935 754545 650046 754550
rect 649986 753838 650046 754545
rect 677242 754398 677248 754462
rect 677312 754398 677318 754462
rect 677250 753986 677310 754398
rect 673359 753276 673425 753279
rect 673359 753274 674784 753276
rect 673359 753218 673364 753274
rect 673420 753218 674784 753274
rect 673359 753216 674784 753218
rect 673359 753213 673425 753216
rect 42063 753130 42129 753131
rect 42063 753128 42112 753130
rect 42020 753126 42112 753128
rect 42020 753070 42068 753126
rect 42020 753068 42112 753070
rect 42063 753066 42112 753068
rect 42176 753066 42182 753130
rect 42063 753065 42129 753066
rect 673071 752388 673137 752391
rect 673071 752386 674784 752388
rect 673071 752330 673076 752386
rect 673132 752330 674784 752386
rect 673071 752328 674784 752330
rect 673071 752325 673137 752328
rect 42063 751796 42129 751799
rect 42490 751796 42496 751798
rect 42063 751794 42496 751796
rect 42063 751738 42068 751794
rect 42124 751738 42496 751794
rect 42063 751736 42496 751738
rect 42063 751733 42129 751736
rect 42490 751734 42496 751736
rect 42560 751734 42566 751798
rect 43066 751734 43072 751798
rect 43136 751796 43142 751798
rect 43215 751796 43281 751799
rect 43136 751794 43281 751796
rect 43136 751738 43220 751794
rect 43276 751738 43281 751794
rect 43136 751736 43281 751738
rect 43136 751734 43142 751736
rect 43215 751733 43281 751736
rect 673263 751648 673329 751651
rect 673263 751646 674784 751648
rect 673263 751590 673268 751646
rect 673324 751590 674784 751646
rect 673263 751588 674784 751590
rect 673263 751585 673329 751588
rect 42063 751056 42129 751059
rect 42682 751056 42688 751058
rect 42063 751054 42688 751056
rect 42063 750998 42068 751054
rect 42124 750998 42688 751054
rect 42063 750996 42688 750998
rect 42063 750993 42129 750996
rect 42682 750994 42688 750996
rect 42752 750994 42758 751058
rect 679746 750171 679806 750730
rect 679746 750166 679857 750171
rect 679746 750110 679796 750166
rect 679852 750110 679857 750166
rect 679746 750108 679857 750110
rect 679791 750105 679857 750108
rect 679791 749576 679857 749579
rect 679746 749574 679857 749576
rect 679746 749518 679796 749574
rect 679852 749518 679857 749574
rect 679746 749513 679857 749518
rect 679746 749250 679806 749513
rect 40954 748626 40960 748690
rect 41024 748688 41030 748690
rect 41775 748688 41841 748691
rect 41914 748688 41920 748690
rect 41024 748686 41920 748688
rect 41024 748630 41780 748686
rect 41836 748630 41920 748686
rect 41024 748628 41920 748630
rect 41024 748626 41030 748628
rect 41775 748625 41841 748628
rect 41914 748626 41920 748628
rect 41984 748626 41990 748690
rect 41775 747506 41841 747507
rect 41722 747504 41728 747506
rect 41684 747444 41728 747504
rect 41792 747502 41841 747506
rect 41836 747446 41841 747502
rect 41722 747442 41728 747444
rect 41792 747442 41841 747446
rect 41775 747441 41841 747442
rect 41722 747294 41728 747358
rect 41792 747356 41798 747358
rect 41871 747356 41937 747359
rect 42106 747356 42112 747358
rect 41792 747354 42112 747356
rect 41792 747298 41876 747354
rect 41932 747298 42112 747354
rect 41792 747296 42112 747298
rect 41792 747294 41798 747296
rect 41871 747293 41937 747296
rect 42106 747294 42112 747296
rect 42176 747294 42182 747358
rect 40762 747146 40768 747210
rect 40832 747208 40838 747210
rect 43023 747208 43089 747211
rect 40832 747206 43089 747208
rect 40832 747150 43028 747206
rect 43084 747150 43089 747206
rect 40832 747148 43089 747150
rect 40832 747146 40838 747148
rect 43023 747145 43089 747148
rect 41146 746702 41152 746766
rect 41216 746764 41222 746766
rect 42927 746764 42993 746767
rect 41216 746762 42993 746764
rect 41216 746706 42932 746762
rect 42988 746706 42993 746762
rect 41216 746704 42993 746706
rect 41216 746702 41222 746704
rect 42927 746701 42993 746704
rect 42447 746024 42513 746027
rect 42874 746024 42880 746026
rect 42447 746022 42880 746024
rect 42447 745966 42452 746022
rect 42508 745966 42880 746022
rect 42447 745964 42880 745966
rect 42447 745961 42513 745964
rect 42874 745962 42880 745964
rect 42944 745962 42950 746026
rect 59535 745580 59601 745583
rect 59535 745578 64416 745580
rect 59535 745522 59540 745578
rect 59596 745522 64416 745578
rect 59535 745520 64416 745522
rect 59535 745517 59601 745520
rect 674554 743150 674560 743214
rect 674624 743212 674630 743214
rect 675375 743212 675441 743215
rect 674624 743210 675441 743212
rect 674624 743154 675380 743210
rect 675436 743154 675441 743210
rect 674624 743152 675441 743154
rect 674624 743150 674630 743152
rect 675375 743149 675441 743152
rect 675759 742472 675825 742475
rect 676666 742472 676672 742474
rect 675759 742470 676672 742472
rect 675759 742414 675764 742470
rect 675820 742414 676672 742470
rect 675759 742412 676672 742414
rect 675759 742409 675825 742412
rect 676666 742410 676672 742412
rect 676736 742410 676742 742474
rect 653967 742176 654033 742179
rect 650208 742174 654033 742176
rect 650208 742118 653972 742174
rect 654028 742118 654033 742174
rect 650208 742116 654033 742118
rect 653967 742113 654033 742116
rect 675759 741732 675825 741735
rect 676090 741732 676096 741734
rect 675759 741730 676096 741732
rect 675759 741674 675764 741730
rect 675820 741674 676096 741730
rect 675759 741672 676096 741674
rect 675759 741669 675825 741672
rect 676090 741670 676096 741672
rect 676160 741670 676166 741734
rect 674938 740338 674944 740402
rect 675008 740400 675014 740402
rect 675471 740400 675537 740403
rect 675008 740398 675537 740400
rect 675008 740342 675476 740398
rect 675532 740342 675537 740398
rect 675008 740340 675537 740342
rect 675008 740338 675014 740340
rect 675471 740337 675537 740340
rect 674746 739302 674752 739366
rect 674816 739364 674822 739366
rect 675471 739364 675537 739367
rect 674816 739362 675537 739364
rect 674816 739306 675476 739362
rect 675532 739306 675537 739362
rect 674816 739304 675537 739306
rect 674816 739302 674822 739304
rect 675471 739301 675537 739304
rect 675375 738626 675441 738627
rect 675322 738624 675328 738626
rect 675284 738564 675328 738624
rect 675392 738622 675441 738626
rect 675436 738566 675441 738622
rect 675322 738562 675328 738564
rect 675392 738562 675441 738566
rect 675375 738561 675441 738562
rect 42831 737292 42897 737295
rect 42336 737290 42897 737292
rect 42336 737234 42836 737290
rect 42892 737234 42897 737290
rect 42336 737232 42897 737234
rect 42831 737229 42897 737232
rect 42159 736700 42225 736703
rect 42114 736698 42225 736700
rect 42114 736642 42164 736698
rect 42220 736642 42225 736698
rect 42114 736637 42225 736642
rect 42114 736522 42174 736637
rect 42831 735664 42897 735667
rect 42336 735662 42897 735664
rect 42336 735606 42836 735662
rect 42892 735606 42897 735662
rect 42336 735604 42897 735606
rect 42831 735601 42897 735604
rect 43215 734924 43281 734927
rect 42336 734922 43281 734924
rect 42336 734866 43220 734922
rect 43276 734866 43281 734922
rect 42336 734864 43281 734866
rect 43215 734861 43281 734864
rect 43311 734036 43377 734039
rect 42336 734034 43377 734036
rect 42336 733978 43316 734034
rect 43372 733978 43377 734034
rect 42336 733976 43377 733978
rect 43311 733973 43377 733976
rect 41530 733826 41536 733890
rect 41600 733826 41606 733890
rect 41538 733340 41598 733826
rect 41338 733086 41344 733150
rect 41408 733086 41414 733150
rect 41346 732556 41406 733086
rect 41346 732526 42144 732556
rect 41376 732496 42174 732526
rect 42114 732262 42174 732496
rect 42106 732198 42112 732262
rect 42176 732198 42182 732262
rect 677050 731754 677056 731818
rect 677120 731754 677126 731818
rect 42306 731668 42366 731712
rect 43119 731668 43185 731671
rect 42306 731666 43185 731668
rect 42306 731610 43124 731666
rect 43180 731610 43185 731666
rect 42306 731608 43185 731610
rect 43119 731605 43185 731608
rect 59535 731076 59601 731079
rect 59535 731074 64416 731076
rect 59535 731018 59540 731074
rect 59596 731018 64416 731074
rect 59535 731016 64416 731018
rect 59535 731013 59601 731016
rect 40194 730339 40254 730898
rect 655215 730484 655281 730487
rect 650208 730482 655281 730484
rect 650208 730426 655220 730482
rect 655276 730426 655281 730482
rect 650208 730424 655281 730426
rect 655215 730421 655281 730424
rect 40194 730334 40305 730339
rect 40194 730278 40244 730334
rect 40300 730278 40305 730334
rect 40194 730276 40305 730278
rect 40239 730273 40305 730276
rect 42306 729596 42366 730084
rect 43066 729596 43072 729598
rect 42306 729536 43072 729596
rect 43066 729534 43072 729536
rect 43136 729534 43142 729598
rect 41730 728859 41790 729270
rect 41679 728854 41790 728859
rect 41679 728798 41684 728854
rect 41740 728798 41790 728854
rect 41679 728796 41790 728798
rect 41679 728793 41745 728796
rect 41730 727971 41790 728530
rect 677058 728116 677118 731754
rect 677818 728116 677824 728118
rect 677058 728056 677824 728116
rect 677818 728054 677824 728056
rect 677888 728054 677894 728118
rect 41730 727966 41841 727971
rect 41730 727910 41780 727966
rect 41836 727910 41841 727966
rect 41730 727908 41841 727910
rect 41775 727905 41841 727908
rect 674703 727968 674769 727971
rect 677050 727968 677056 727970
rect 674703 727966 677056 727968
rect 674703 727910 674708 727966
rect 674764 727910 677056 727966
rect 674703 727908 677056 727910
rect 674703 727905 674769 727908
rect 677050 727906 677056 727908
rect 677120 727906 677126 727970
rect 41922 727231 41982 727790
rect 41871 727226 41982 727231
rect 41871 727170 41876 727226
rect 41932 727170 41982 727226
rect 41871 727168 41982 727170
rect 41871 727165 41937 727168
rect 41154 726342 41214 726902
rect 41146 726278 41152 726342
rect 41216 726278 41222 726342
rect 41538 725899 41598 726162
rect 41538 725894 41649 725899
rect 41538 725838 41588 725894
rect 41644 725838 41649 725894
rect 41538 725836 41649 725838
rect 41583 725833 41649 725836
rect 42106 725538 42112 725602
rect 42176 725600 42182 725602
rect 43450 725600 43456 725602
rect 42176 725540 43456 725600
rect 42176 725538 42182 725540
rect 43450 725538 43456 725540
rect 43520 725538 43526 725602
rect 42114 724715 42174 725274
rect 42114 724710 42225 724715
rect 42114 724654 42164 724710
rect 42220 724654 42225 724710
rect 42114 724652 42225 724654
rect 42159 724649 42225 724652
rect 41922 724123 41982 724534
rect 41922 724118 42033 724123
rect 41922 724062 41972 724118
rect 42028 724062 42033 724118
rect 41922 724060 42033 724062
rect 41967 724057 42033 724060
rect 41538 723235 41598 723794
rect 41487 723230 41598 723235
rect 41487 723174 41492 723230
rect 41548 723174 41598 723230
rect 41487 723172 41598 723174
rect 41487 723169 41553 723172
rect 41346 722791 41406 723054
rect 41346 722786 41457 722791
rect 41346 722730 41396 722786
rect 41452 722730 41457 722786
rect 41346 722728 41457 722730
rect 41391 722725 41457 722728
rect 41914 722430 41920 722494
rect 41984 722492 41990 722494
rect 42490 722492 42496 722494
rect 41984 722432 42496 722492
rect 41984 722430 41990 722432
rect 42490 722430 42496 722432
rect 42560 722430 42566 722494
rect 674415 722492 674481 722495
rect 674415 722490 674784 722492
rect 674415 722434 674420 722490
rect 674476 722434 674784 722490
rect 674415 722432 674784 722434
rect 674415 722429 674481 722432
rect 42114 722051 42174 722166
rect 42063 722046 42174 722051
rect 42063 721990 42068 722046
rect 42124 721990 42174 722046
rect 42063 721988 42174 721990
rect 42063 721985 42129 721988
rect 674703 721900 674769 721903
rect 674703 721898 674814 721900
rect 674703 721842 674708 721898
rect 674764 721842 674814 721898
rect 674703 721837 674814 721842
rect 674754 721722 674814 721837
rect 43258 721456 43264 721458
rect 42336 721396 43264 721456
rect 43258 721394 43264 721396
rect 43328 721394 43334 721458
rect 674415 720864 674481 720867
rect 674415 720862 674784 720864
rect 674415 720806 674420 720862
rect 674476 720806 674784 720862
rect 674415 720804 674784 720806
rect 674415 720801 674481 720804
rect 42306 720420 42366 720538
rect 42447 720420 42513 720423
rect 42306 720418 42513 720420
rect 42306 720362 42452 720418
rect 42508 720362 42513 720418
rect 42306 720360 42513 720362
rect 42447 720357 42513 720360
rect 674703 720272 674769 720275
rect 674703 720270 674814 720272
rect 674703 720214 674708 720270
rect 674764 720214 674814 720270
rect 674703 720209 674814 720214
rect 674754 720094 674814 720209
rect 674754 719091 674814 719206
rect 674703 719086 674814 719091
rect 42306 718792 42366 719058
rect 674703 719030 674708 719086
rect 674764 719030 674814 719086
rect 674703 719028 674814 719030
rect 674703 719025 674769 719028
rect 42447 718792 42513 718795
rect 42306 718790 42513 718792
rect 42306 718734 42452 718790
rect 42508 718734 42513 718790
rect 42306 718732 42513 718734
rect 42447 718729 42513 718732
rect 654255 718644 654321 718647
rect 650208 718642 654321 718644
rect 650208 718586 654260 718642
rect 654316 718586 654321 718642
rect 650208 718584 654321 718586
rect 654255 718581 654321 718584
rect 672111 718496 672177 718499
rect 674754 718496 674814 718540
rect 672111 718494 674814 718496
rect 672111 718438 672116 718494
rect 672172 718438 674814 718494
rect 672111 718436 674814 718438
rect 672111 718433 672177 718436
rect 674754 717164 674814 717726
rect 674370 717104 674814 717164
rect 673935 717018 674001 717019
rect 673935 717016 673984 717018
rect 673856 717014 673984 717016
rect 674048 717016 674054 717018
rect 674370 717016 674430 717104
rect 676474 717102 676480 717166
rect 676544 717102 676550 717166
rect 673856 716958 673940 717014
rect 673856 716956 673984 716958
rect 673935 716954 673984 716956
rect 674048 716956 674430 717016
rect 674048 716954 674054 716956
rect 673935 716953 674001 716954
rect 676482 716912 676542 717102
rect 59535 716720 59601 716723
rect 59535 716718 64416 716720
rect 59535 716662 59540 716718
rect 59596 716662 64416 716718
rect 59535 716660 64416 716662
rect 59535 716657 59601 716660
rect 676282 716658 676288 716722
rect 676352 716658 676358 716722
rect 676290 716098 676350 716658
rect 675706 715770 675712 715834
rect 675776 715770 675782 715834
rect 675714 715284 675774 715770
rect 675898 715030 675904 715094
rect 675968 715030 675974 715094
rect 675906 714470 675966 715030
rect 41487 714352 41553 714355
rect 41914 714352 41920 714354
rect 41487 714350 41920 714352
rect 41487 714294 41492 714350
rect 41548 714294 41920 714350
rect 41487 714292 41920 714294
rect 41487 714289 41553 714292
rect 41914 714290 41920 714292
rect 41984 714290 41990 714354
rect 41391 714206 41457 714207
rect 41338 714204 41344 714206
rect 41300 714144 41344 714204
rect 41408 714202 41457 714206
rect 41452 714146 41457 714202
rect 41338 714142 41344 714144
rect 41408 714142 41457 714146
rect 41391 714141 41457 714142
rect 41679 714204 41745 714207
rect 42874 714204 42880 714206
rect 41679 714202 42880 714204
rect 41679 714146 41684 714202
rect 41740 714146 42880 714202
rect 41679 714144 42880 714146
rect 41679 714141 41745 714144
rect 42874 714142 42880 714144
rect 42944 714142 42950 714206
rect 41775 713910 41841 713911
rect 41722 713908 41728 713910
rect 41684 713848 41728 713908
rect 41792 713906 41841 713910
rect 41836 713850 41841 713906
rect 41722 713846 41728 713848
rect 41792 713846 41841 713850
rect 41775 713845 41841 713846
rect 42159 713908 42225 713911
rect 42682 713908 42688 713910
rect 42159 713906 42688 713908
rect 42159 713850 42164 713906
rect 42220 713850 42688 713906
rect 42159 713848 42688 713850
rect 42159 713845 42225 713848
rect 42682 713846 42688 713848
rect 42752 713846 42758 713910
rect 674362 713698 674368 713762
rect 674432 713760 674438 713762
rect 674432 713700 674784 713760
rect 674432 713698 674438 713700
rect 675130 713550 675136 713614
rect 675200 713550 675206 713614
rect 675138 712990 675198 713550
rect 675514 712662 675520 712726
rect 675584 712662 675590 712726
rect 675522 712102 675582 712662
rect 43407 711540 43473 711543
rect 43122 711538 43473 711540
rect 43122 711482 43412 711538
rect 43468 711482 43473 711538
rect 43122 711480 43473 711482
rect 43122 711395 43182 711480
rect 43407 711477 43473 711480
rect 674703 711540 674769 711543
rect 674703 711538 674814 711540
rect 674703 711482 674708 711538
rect 674764 711482 674814 711538
rect 674703 711477 674814 711482
rect 43119 711390 43185 711395
rect 43119 711334 43124 711390
rect 43180 711334 43185 711390
rect 674754 711362 674814 711477
rect 43119 711329 43185 711334
rect 41338 711034 41344 711098
rect 41408 711096 41414 711098
rect 43023 711096 43089 711099
rect 41408 711094 43089 711096
rect 41408 711038 43028 711094
rect 43084 711038 43089 711094
rect 41408 711036 43089 711038
rect 41408 711034 41414 711036
rect 43023 711033 43089 711036
rect 674415 710504 674481 710507
rect 674415 710502 674784 710504
rect 674415 710446 674420 710502
rect 674476 710446 674784 710502
rect 674415 710444 674784 710446
rect 674415 710441 674481 710444
rect 677818 710294 677824 710358
rect 677888 710294 677894 710358
rect 42682 709702 42688 709766
rect 42752 709764 42758 709766
rect 43119 709764 43185 709767
rect 42752 709762 43185 709764
rect 42752 709706 43124 709762
rect 43180 709706 43185 709762
rect 677826 709734 677886 710294
rect 42752 709704 43185 709706
rect 42752 709702 42758 709704
rect 43119 709701 43185 709704
rect 676858 709406 676864 709470
rect 676928 709406 676934 709470
rect 676866 708994 676926 709406
rect 42063 708580 42129 708583
rect 43258 708580 43264 708582
rect 42063 708578 43264 708580
rect 42063 708522 42068 708578
rect 42124 708522 43264 708578
rect 42063 708520 43264 708522
rect 42063 708517 42129 708520
rect 43258 708518 43264 708520
rect 43328 708518 43334 708582
rect 674703 708432 674769 708435
rect 674703 708430 674814 708432
rect 674703 708374 674708 708430
rect 674764 708374 674814 708430
rect 674703 708369 674814 708374
rect 674754 708254 674814 708369
rect 41871 707990 41937 707991
rect 41871 707988 41920 707990
rect 41828 707986 41920 707988
rect 41828 707930 41876 707986
rect 41828 707928 41920 707930
rect 41871 707926 41920 707928
rect 41984 707926 41990 707990
rect 42735 707988 42801 707991
rect 42874 707988 42880 707990
rect 42735 707986 42880 707988
rect 42735 707930 42740 707986
rect 42796 707930 42880 707986
rect 42735 707928 42880 707930
rect 41871 707925 41937 707926
rect 42735 707925 42801 707928
rect 42874 707926 42880 707928
rect 42944 707926 42950 707990
rect 649743 707544 649809 707547
rect 649743 707542 649854 707544
rect 649743 707486 649748 707542
rect 649804 707486 649854 707542
rect 649743 707481 649854 707486
rect 649794 706922 649854 707481
rect 674415 707396 674481 707399
rect 674415 707394 674784 707396
rect 674415 707338 674420 707394
rect 674476 707338 674784 707394
rect 674415 707336 674784 707338
rect 674415 707333 674481 707336
rect 41775 706806 41841 706807
rect 41722 706804 41728 706806
rect 41684 706744 41728 706804
rect 41792 706802 41841 706806
rect 41836 706746 41841 706802
rect 41722 706742 41728 706744
rect 41792 706742 41841 706746
rect 41775 706741 41841 706742
rect 674703 706804 674769 706807
rect 674703 706802 674814 706804
rect 674703 706746 674708 706802
rect 674764 706746 674814 706802
rect 674703 706741 674814 706746
rect 674754 706626 674814 706741
rect 43450 705916 43456 705918
rect 42306 705856 43456 705916
rect 42306 705770 42366 705856
rect 43450 705854 43456 705856
rect 43520 705854 43526 705918
rect 42298 705706 42304 705770
rect 42368 705706 42374 705770
rect 41146 705410 41152 705474
rect 41216 705472 41222 705474
rect 42447 705472 42513 705475
rect 41216 705470 42513 705472
rect 41216 705414 42452 705470
rect 42508 705414 42513 705470
rect 41216 705412 42513 705414
rect 41216 705410 41222 705412
rect 42447 705409 42513 705412
rect 679746 705179 679806 705738
rect 679746 705174 679857 705179
rect 679746 705118 679796 705174
rect 679852 705118 679857 705174
rect 679746 705116 679857 705118
rect 679791 705113 679857 705116
rect 42063 704734 42129 704735
rect 42063 704732 42112 704734
rect 42020 704730 42112 704732
rect 42176 704732 42182 704734
rect 42490 704732 42496 704734
rect 42020 704674 42068 704730
rect 42020 704672 42112 704674
rect 42063 704670 42112 704672
rect 42176 704672 42496 704732
rect 42176 704670 42182 704672
rect 42490 704670 42496 704672
rect 42560 704670 42566 704734
rect 42063 704669 42129 704670
rect 679791 704584 679857 704587
rect 679746 704582 679857 704584
rect 679746 704526 679796 704582
rect 679852 704526 679857 704582
rect 679746 704521 679857 704526
rect 679746 704258 679806 704521
rect 41775 704142 41841 704143
rect 41722 704078 41728 704142
rect 41792 704140 41841 704142
rect 41792 704138 41884 704140
rect 41836 704082 41884 704138
rect 41792 704080 41884 704082
rect 41792 704078 41841 704080
rect 41775 704077 41841 704078
rect 43023 702810 43089 702811
rect 43023 702808 43072 702810
rect 42980 702806 43072 702808
rect 42980 702750 43028 702806
rect 42980 702748 43072 702750
rect 43023 702746 43072 702748
rect 43136 702746 43142 702810
rect 43023 702745 43089 702746
rect 59535 702364 59601 702367
rect 59535 702362 64416 702364
rect 59535 702306 59540 702362
rect 59596 702306 64416 702362
rect 59535 702304 64416 702306
rect 59535 702301 59601 702304
rect 675471 697926 675537 697927
rect 675471 697922 675520 697926
rect 675584 697924 675590 697926
rect 675471 697866 675476 697922
rect 675471 697862 675520 697866
rect 675584 697864 675628 697924
rect 675584 697862 675590 697864
rect 675471 697861 675537 697862
rect 675759 697332 675825 697335
rect 676474 697332 676480 697334
rect 675759 697330 676480 697332
rect 675759 697274 675764 697330
rect 675820 697274 676480 697330
rect 675759 697272 676480 697274
rect 675759 697269 675825 697272
rect 676474 697270 676480 697272
rect 676544 697270 676550 697334
rect 675759 697184 675825 697187
rect 675898 697184 675904 697186
rect 675759 697182 675904 697184
rect 675759 697126 675764 697182
rect 675820 697126 675904 697182
rect 675759 697124 675904 697126
rect 675759 697121 675825 697124
rect 675898 697122 675904 697124
rect 675968 697122 675974 697186
rect 654447 695260 654513 695263
rect 650208 695258 654513 695260
rect 650208 695202 654452 695258
rect 654508 695202 654513 695258
rect 650208 695200 654513 695202
rect 654447 695197 654513 695200
rect 675663 694818 675729 694819
rect 675663 694814 675712 694818
rect 675776 694816 675782 694818
rect 675663 694758 675668 694814
rect 675663 694754 675712 694758
rect 675776 694756 675820 694816
rect 675776 694754 675782 694756
rect 675663 694753 675729 694754
rect 674170 694310 674176 694374
rect 674240 694372 674246 694374
rect 675471 694372 675537 694375
rect 674240 694370 675537 694372
rect 674240 694314 675476 694370
rect 675532 694314 675537 694370
rect 674240 694312 675537 694314
rect 674240 694310 674246 694312
rect 675471 694309 675537 694312
rect 42831 694076 42897 694079
rect 42336 694074 42897 694076
rect 42336 694018 42836 694074
rect 42892 694018 42897 694074
rect 42336 694016 42897 694018
rect 42831 694013 42897 694016
rect 42447 693484 42513 693487
rect 42306 693482 42513 693484
rect 42306 693426 42452 693482
rect 42508 693426 42513 693482
rect 42306 693424 42513 693426
rect 42306 693306 42366 693424
rect 42447 693421 42513 693424
rect 674362 693422 674368 693486
rect 674432 693484 674438 693486
rect 675471 693484 675537 693487
rect 674432 693482 675537 693484
rect 674432 693426 675476 693482
rect 675532 693426 675537 693482
rect 674432 693424 675537 693426
rect 674432 693422 674438 693424
rect 675471 693421 675537 693424
rect 42447 692744 42513 692747
rect 42306 692742 42513 692744
rect 42306 692686 42452 692742
rect 42508 692686 42513 692742
rect 42306 692684 42513 692686
rect 42306 692418 42366 692684
rect 42447 692681 42513 692684
rect 43503 691708 43569 691711
rect 42336 691706 43569 691708
rect 42336 691650 43508 691706
rect 43564 691650 43569 691706
rect 42336 691648 43569 691650
rect 43503 691645 43569 691648
rect 675759 691708 675825 691711
rect 676282 691708 676288 691710
rect 675759 691706 676288 691708
rect 675759 691650 675764 691706
rect 675820 691650 676288 691706
rect 675759 691648 676288 691650
rect 675759 691645 675825 691648
rect 676282 691646 676288 691648
rect 676352 691646 676358 691710
rect 43215 690820 43281 690823
rect 42336 690818 43281 690820
rect 42336 690762 43220 690818
rect 43276 690762 43281 690818
rect 42336 690760 43281 690762
rect 43215 690757 43281 690760
rect 41530 690314 41536 690378
rect 41600 690314 41606 690378
rect 41538 690228 41598 690314
rect 41538 690198 42144 690228
rect 41568 690168 42174 690198
rect 42114 689638 42174 690168
rect 42106 689574 42112 689638
rect 42176 689574 42182 689638
rect 42306 688750 42366 689310
rect 675130 689130 675136 689194
rect 675200 689192 675206 689194
rect 675375 689192 675441 689195
rect 675200 689190 675441 689192
rect 675200 689134 675380 689190
rect 675436 689134 675441 689190
rect 675200 689132 675441 689134
rect 675200 689130 675206 689132
rect 675375 689129 675441 689132
rect 42298 688686 42304 688750
rect 42368 688686 42374 688750
rect 41730 688307 41790 688496
rect 41679 688302 41790 688307
rect 41679 688246 41684 688302
rect 41740 688246 41790 688302
rect 41679 688244 41790 688246
rect 41679 688241 41745 688244
rect 59535 688008 59601 688011
rect 59535 688006 64416 688008
rect 59535 687950 59540 688006
rect 59596 687950 64416 688006
rect 59535 687948 64416 687950
rect 59535 687945 59601 687948
rect 40194 687123 40254 687682
rect 674895 687564 674961 687567
rect 676858 687564 676864 687566
rect 674895 687562 676864 687564
rect 674895 687506 674900 687562
rect 674956 687506 676864 687562
rect 674895 687504 676864 687506
rect 674895 687501 674961 687504
rect 676858 687502 676864 687504
rect 676928 687502 676934 687566
rect 40143 687118 40254 687123
rect 40143 687062 40148 687118
rect 40204 687062 40254 687118
rect 40143 687060 40254 687062
rect 40143 687057 40209 687060
rect 40194 686383 40254 686868
rect 40194 686378 40305 686383
rect 40194 686322 40244 686378
rect 40300 686322 40305 686378
rect 40194 686320 40305 686322
rect 40239 686317 40305 686320
rect 41730 685643 41790 686054
rect 41730 685638 41841 685643
rect 41730 685582 41780 685638
rect 41836 685582 41841 685638
rect 41730 685580 41841 685582
rect 41775 685577 41841 685580
rect 40962 684903 41022 685388
rect 40911 684898 41022 684903
rect 40911 684842 40916 684898
rect 40972 684842 41022 684898
rect 40911 684840 41022 684842
rect 40911 684837 40977 684840
rect 41922 684015 41982 684574
rect 41922 684010 42033 684015
rect 41922 683954 41972 684010
rect 42028 683954 42033 684010
rect 41922 683952 42033 683954
rect 41967 683949 42033 683952
rect 37314 683275 37374 683760
rect 655407 683568 655473 683571
rect 650208 683566 655473 683568
rect 650208 683510 655412 683566
rect 655468 683510 655473 683566
rect 650208 683508 655473 683510
rect 655407 683505 655473 683508
rect 37314 683270 37425 683275
rect 37314 683214 37364 683270
rect 37420 683214 37425 683270
rect 37314 683212 37425 683214
rect 37359 683209 37425 683212
rect 42114 682683 42174 682946
rect 42063 682678 42174 682683
rect 42063 682622 42068 682678
rect 42124 682622 42174 682678
rect 42063 682620 42174 682622
rect 42063 682617 42129 682620
rect 41346 681499 41406 682058
rect 41295 681494 41406 681499
rect 41295 681438 41300 681494
rect 41356 681438 41406 681494
rect 41295 681436 41406 681438
rect 41295 681433 41361 681436
rect 43023 681348 43089 681351
rect 42336 681346 43089 681348
rect 42336 681290 43028 681346
rect 43084 681290 43089 681346
rect 42336 681288 43089 681290
rect 43023 681285 43089 681288
rect 43887 680608 43953 680611
rect 42336 680606 43953 680608
rect 42336 680550 43892 680606
rect 43948 680550 43953 680606
rect 42336 680548 43953 680550
rect 43887 680545 43953 680548
rect 41922 679575 41982 679838
rect 41871 679570 41982 679575
rect 41871 679514 41876 679570
rect 41932 679514 41982 679570
rect 41871 679512 41982 679514
rect 41871 679509 41937 679512
rect 42114 678835 42174 678950
rect 42114 678830 42225 678835
rect 42114 678774 42164 678830
rect 42220 678774 42225 678830
rect 42114 678772 42225 678774
rect 42159 678769 42225 678772
rect 43119 678240 43185 678243
rect 42336 678238 43185 678240
rect 42336 678182 43124 678238
rect 43180 678182 43185 678238
rect 42336 678180 43185 678182
rect 43119 678177 43185 678180
rect 674703 677500 674769 677503
rect 674703 677498 674814 677500
rect 674703 677442 674708 677498
rect 674764 677442 674814 677498
rect 674703 677437 674814 677442
rect 674754 677322 674814 677437
rect 42306 676760 42366 677322
rect 42447 676760 42513 676763
rect 42306 676758 42513 676760
rect 42306 676702 42452 676758
rect 42508 676702 42513 676758
rect 42306 676700 42513 676702
rect 42447 676697 42513 676700
rect 674703 676760 674769 676763
rect 674703 676758 674814 676760
rect 674703 676702 674708 676758
rect 674764 676702 674814 676758
rect 674703 676697 674814 676702
rect 674754 676434 674814 676697
rect 674703 675872 674769 675875
rect 674703 675870 674814 675872
rect 42306 675724 42366 675842
rect 674703 675814 674708 675870
rect 674764 675814 674814 675870
rect 674703 675809 674814 675814
rect 42447 675724 42513 675727
rect 42306 675722 42513 675724
rect 42306 675666 42452 675722
rect 42508 675666 42513 675722
rect 674754 675694 674814 675809
rect 42306 675664 42513 675666
rect 42447 675661 42513 675664
rect 41914 675366 41920 675430
rect 41984 675428 41990 675430
rect 42874 675428 42880 675430
rect 41984 675368 42880 675428
rect 41984 675366 41990 675368
rect 42874 675366 42880 675368
rect 42944 675366 42950 675430
rect 673839 674836 673905 674839
rect 673839 674834 674784 674836
rect 673839 674778 673844 674834
rect 673900 674778 674784 674834
rect 673839 674776 674784 674778
rect 673839 674773 673905 674776
rect 673263 674096 673329 674099
rect 673263 674094 674784 674096
rect 673263 674038 673268 674094
rect 673324 674038 674784 674094
rect 673263 674036 674784 674038
rect 673263 674033 673329 674036
rect 40239 673948 40305 673951
rect 40762 673948 40768 673950
rect 40239 673946 40768 673948
rect 40239 673890 40244 673946
rect 40300 673890 40768 673946
rect 40239 673888 40768 673890
rect 40239 673885 40305 673888
rect 40762 673886 40768 673888
rect 40832 673886 40838 673950
rect 59535 673652 59601 673655
rect 59535 673650 64416 673652
rect 59535 673594 59540 673650
rect 59596 673594 64416 673650
rect 59535 673592 64416 673594
rect 59535 673589 59601 673592
rect 673743 673356 673809 673359
rect 673743 673354 674784 673356
rect 673743 673298 673748 673354
rect 673804 673298 674784 673354
rect 673743 673296 674784 673298
rect 673743 673293 673809 673296
rect 673978 672998 673984 673062
rect 674048 673060 674054 673062
rect 674048 673000 674814 673060
rect 674048 672998 674054 673000
rect 37359 672616 37425 672619
rect 40570 672616 40576 672618
rect 37359 672614 40576 672616
rect 37359 672558 37364 672614
rect 37420 672558 40576 672614
rect 37359 672556 40576 672558
rect 37359 672553 37425 672556
rect 40570 672554 40576 672556
rect 40640 672554 40646 672618
rect 674754 672323 674814 673000
rect 674703 672318 674814 672323
rect 674703 672262 674708 672318
rect 674764 672262 674814 672318
rect 674703 672260 674814 672262
rect 674703 672257 674769 672260
rect 676090 672258 676096 672322
rect 676160 672258 676166 672322
rect 654447 671728 654513 671731
rect 650208 671726 654513 671728
rect 650208 671670 654452 671726
rect 654508 671670 654513 671726
rect 676098 671698 676158 672258
rect 650208 671668 654513 671670
rect 654447 671665 654513 671668
rect 674511 671136 674577 671139
rect 674511 671134 674814 671136
rect 674511 671078 674516 671134
rect 674572 671078 674814 671134
rect 674511 671076 674814 671078
rect 674511 671073 674577 671076
rect 41295 670988 41361 670991
rect 41722 670988 41728 670990
rect 41295 670986 41728 670988
rect 41295 670930 41300 670986
rect 41356 670930 41728 670986
rect 41295 670928 41728 670930
rect 41295 670925 41361 670928
rect 41722 670926 41728 670928
rect 41792 670926 41798 670990
rect 42159 670988 42225 670991
rect 43119 670990 43185 670991
rect 42682 670988 42688 670990
rect 42159 670986 42688 670988
rect 42159 670930 42164 670986
rect 42220 670930 42688 670986
rect 42159 670928 42688 670930
rect 42159 670925 42225 670928
rect 42682 670926 42688 670928
rect 42752 670926 42758 670990
rect 43066 670988 43072 670990
rect 43028 670928 43072 670988
rect 43136 670986 43185 670990
rect 43180 670930 43185 670986
rect 43066 670926 43072 670928
rect 43136 670926 43185 670930
rect 43119 670925 43185 670926
rect 674754 670884 674814 671076
rect 41967 670842 42033 670843
rect 41914 670778 41920 670842
rect 41984 670840 42033 670842
rect 42159 670840 42225 670843
rect 42490 670840 42496 670842
rect 41984 670838 42076 670840
rect 42028 670782 42076 670838
rect 41984 670780 42076 670782
rect 42159 670838 42496 670840
rect 42159 670782 42164 670838
rect 42220 670782 42496 670838
rect 42159 670780 42496 670782
rect 41984 670778 42033 670780
rect 41967 670777 42033 670778
rect 42159 670777 42225 670780
rect 42490 670778 42496 670780
rect 42560 670778 42566 670842
rect 42063 670692 42129 670695
rect 42063 670690 42174 670692
rect 42063 670634 42068 670690
rect 42124 670634 42174 670690
rect 42063 670629 42174 670634
rect 42114 670399 42174 670629
rect 674554 670482 674560 670546
rect 674624 670544 674630 670546
rect 674624 670484 674814 670544
rect 674624 670482 674630 670484
rect 42114 670394 42225 670399
rect 42114 670338 42164 670394
rect 42220 670338 42225 670394
rect 42114 670336 42225 670338
rect 42159 670333 42225 670336
rect 674754 670070 674814 670484
rect 674938 669742 674944 669806
rect 675008 669742 675014 669806
rect 674946 669256 675006 669742
rect 674319 668620 674385 668623
rect 674319 668618 674784 668620
rect 674319 668562 674324 668618
rect 674380 668562 674784 668618
rect 674319 668560 674784 668562
rect 674319 668557 674385 668560
rect 674223 667806 674289 667809
rect 674223 667804 674784 667806
rect 674223 667748 674228 667804
rect 674284 667748 674784 667804
rect 674223 667746 674784 667748
rect 674223 667743 674289 667746
rect 676666 667522 676672 667586
rect 676736 667522 676742 667586
rect 676674 666962 676734 667522
rect 674746 666634 674752 666698
rect 674816 666634 674822 666698
rect 674754 666074 674814 666634
rect 675322 665894 675328 665958
rect 675392 665894 675398 665958
rect 42159 665364 42225 665367
rect 43066 665364 43072 665366
rect 42159 665362 43072 665364
rect 42159 665306 42164 665362
rect 42220 665306 43072 665362
rect 42159 665304 43072 665306
rect 42159 665301 42225 665304
rect 43066 665302 43072 665304
rect 43136 665302 43142 665366
rect 675330 665334 675390 665894
rect 673839 664476 673905 664479
rect 673839 664474 674784 664476
rect 673839 664418 673844 664474
rect 673900 664418 674784 664474
rect 673839 664416 674784 664418
rect 673839 664413 673905 664416
rect 673839 663884 673905 663887
rect 673839 663882 674784 663884
rect 673839 663826 673844 663882
rect 673900 663826 674784 663882
rect 673839 663824 674784 663826
rect 673839 663821 673905 663824
rect 677050 663526 677056 663590
rect 677120 663526 677126 663590
rect 42682 663378 42688 663442
rect 42752 663440 42758 663442
rect 42831 663440 42897 663443
rect 42752 663438 42897 663440
rect 42752 663382 42836 663438
rect 42892 663382 42897 663438
rect 42752 663380 42897 663382
rect 42752 663378 42758 663380
rect 42831 663377 42897 663380
rect 677058 662966 677118 663526
rect 42447 662850 42513 662851
rect 42447 662846 42496 662850
rect 42560 662848 42566 662850
rect 42447 662790 42452 662846
rect 42447 662786 42496 662790
rect 42560 662788 42604 662848
rect 42560 662786 42566 662788
rect 42447 662785 42513 662786
rect 40762 662342 40768 662406
rect 40832 662404 40838 662406
rect 43119 662404 43185 662407
rect 40832 662402 43185 662404
rect 40832 662346 43124 662402
rect 43180 662346 43185 662402
rect 40832 662344 43185 662346
rect 40832 662342 40838 662344
rect 43119 662341 43185 662344
rect 673359 662256 673425 662259
rect 673359 662254 674784 662256
rect 673359 662198 673364 662254
rect 673420 662198 674784 662254
rect 673359 662196 674784 662198
rect 673359 662193 673425 662196
rect 42159 661516 42225 661519
rect 42490 661516 42496 661518
rect 42159 661514 42496 661516
rect 42159 661458 42164 661514
rect 42220 661458 42496 661514
rect 42159 661456 42496 661458
rect 42159 661453 42225 661456
rect 42490 661454 42496 661456
rect 42560 661454 42566 661518
rect 673167 661368 673233 661371
rect 673167 661366 674784 661368
rect 673167 661310 673172 661366
rect 673228 661310 674784 661366
rect 673167 661308 674784 661310
rect 673167 661305 673233 661308
rect 41146 660714 41152 660778
rect 41216 660776 41222 660778
rect 42159 660776 42225 660779
rect 41216 660774 42225 660776
rect 41216 660718 42164 660774
rect 42220 660718 42225 660774
rect 41216 660716 42225 660718
rect 41216 660714 41222 660716
rect 41775 660334 41841 660335
rect 41722 660332 41728 660334
rect 41684 660272 41728 660332
rect 41792 660330 41841 660334
rect 41836 660274 41841 660330
rect 41722 660270 41728 660272
rect 41792 660270 41841 660274
rect 41775 660269 41841 660270
rect 41722 660122 41728 660186
rect 41792 660184 41798 660186
rect 41922 660184 41982 660716
rect 42159 660713 42225 660716
rect 649839 660628 649905 660631
rect 41792 660124 41982 660184
rect 649794 660626 649905 660628
rect 649794 660570 649844 660626
rect 649900 660570 649905 660626
rect 649794 660565 649905 660570
rect 41792 660122 41798 660124
rect 649794 660006 649854 660565
rect 679746 660039 679806 660598
rect 679695 660034 679806 660039
rect 679695 659978 679700 660034
rect 679756 659978 679806 660034
rect 679695 659976 679806 659978
rect 679695 659973 679761 659976
rect 59535 659296 59601 659299
rect 679695 659296 679761 659299
rect 59535 659294 64416 659296
rect 59535 659238 59540 659294
rect 59596 659238 64416 659294
rect 59535 659236 64416 659238
rect 679695 659294 679806 659296
rect 679695 659238 679700 659294
rect 679756 659238 679806 659294
rect 59535 659233 59601 659236
rect 679695 659233 679806 659238
rect 41871 659150 41937 659151
rect 41871 659146 41920 659150
rect 41984 659148 41990 659150
rect 41871 659090 41876 659146
rect 41871 659086 41920 659090
rect 41984 659088 42028 659148
rect 679746 659118 679806 659233
rect 41984 659086 41990 659088
rect 41871 659085 41937 659086
rect 41914 658938 41920 659002
rect 41984 659000 41990 659002
rect 42490 659000 42496 659002
rect 41984 658940 42496 659000
rect 41984 658938 41990 658940
rect 42490 658938 42496 658940
rect 42560 658938 42566 659002
rect 40570 656570 40576 656634
rect 40640 656632 40646 656634
rect 41775 656632 41841 656635
rect 40640 656630 41841 656632
rect 40640 656574 41780 656630
rect 41836 656574 41841 656630
rect 40640 656572 41841 656574
rect 40640 656570 40646 656572
rect 41775 656569 41841 656572
rect 674799 653672 674865 653675
rect 676282 653672 676288 653674
rect 674799 653670 676288 653672
rect 674799 653614 674804 653670
rect 674860 653614 676288 653670
rect 674799 653612 676288 653614
rect 674799 653609 674865 653612
rect 676282 653610 676288 653612
rect 676352 653610 676358 653674
rect 675375 652638 675441 652639
rect 675322 652636 675328 652638
rect 675284 652576 675328 652636
rect 675392 652634 675441 652638
rect 675436 652578 675441 652634
rect 675322 652574 675328 652576
rect 675392 652574 675441 652578
rect 675375 652573 675441 652574
rect 674554 652130 674560 652194
rect 674624 652192 674630 652194
rect 675471 652192 675537 652195
rect 674624 652190 675537 652192
rect 674624 652134 675476 652190
rect 675532 652134 675537 652190
rect 674624 652132 675537 652134
rect 674624 652130 674630 652132
rect 675471 652129 675537 652132
rect 674938 651390 674944 651454
rect 675008 651452 675014 651454
rect 675471 651452 675537 651455
rect 675008 651450 675537 651452
rect 675008 651394 675476 651450
rect 675532 651394 675537 651450
rect 675008 651392 675537 651394
rect 675008 651390 675014 651392
rect 675471 651389 675537 651392
rect 42447 651156 42513 651159
rect 42306 651154 42513 651156
rect 42306 651098 42452 651154
rect 42508 651098 42513 651154
rect 42306 651096 42513 651098
rect 42306 650830 42366 651096
rect 42447 651093 42513 651096
rect 42306 649824 42366 650090
rect 42447 649824 42513 649827
rect 42306 649822 42513 649824
rect 42306 649766 42452 649822
rect 42508 649766 42513 649822
rect 42306 649764 42513 649766
rect 42447 649761 42513 649764
rect 675759 649824 675825 649827
rect 676666 649824 676672 649826
rect 675759 649822 676672 649824
rect 675759 649766 675764 649822
rect 675820 649766 676672 649822
rect 675759 649764 676672 649766
rect 675759 649761 675825 649764
rect 676666 649762 676672 649764
rect 676736 649762 676742 649826
rect 42447 649528 42513 649531
rect 42306 649526 42513 649528
rect 42306 649470 42452 649526
rect 42508 649470 42513 649526
rect 42306 649468 42513 649470
rect 42306 649202 42366 649468
rect 42447 649465 42513 649468
rect 674746 648874 674752 648938
rect 674816 648936 674822 648938
rect 675471 648936 675537 648939
rect 674816 648934 675537 648936
rect 674816 648878 675476 648934
rect 675532 648878 675537 648934
rect 674816 648876 675537 648878
rect 674816 648874 674822 648876
rect 675471 648873 675537 648876
rect 43215 648492 43281 648495
rect 42336 648490 43281 648492
rect 42336 648434 43220 648490
rect 43276 648434 43281 648490
rect 42336 648432 43281 648434
rect 43215 648429 43281 648432
rect 654255 648344 654321 648347
rect 650208 648342 654321 648344
rect 650208 648286 654260 648342
rect 654316 648286 654321 648342
rect 650208 648284 654321 648286
rect 654255 648281 654321 648284
rect 43503 647604 43569 647607
rect 42336 647602 43569 647604
rect 42336 647546 43508 647602
rect 43564 647546 43569 647602
rect 42336 647544 43569 647546
rect 43503 647541 43569 647544
rect 42106 647394 42112 647458
rect 42176 647394 42182 647458
rect 42114 647012 42174 647394
rect 43599 647012 43665 647015
rect 42114 647010 43665 647012
rect 42114 646982 43604 647010
rect 42144 646954 43604 646982
rect 43660 646954 43665 647010
rect 42144 646952 43665 646954
rect 43599 646949 43665 646952
rect 42298 646654 42304 646718
rect 42368 646654 42374 646718
rect 42306 646124 42366 646654
rect 43791 646124 43857 646127
rect 42306 646122 43857 646124
rect 42306 646094 43796 646122
rect 42336 646066 43796 646094
rect 43852 646066 43857 646122
rect 42336 646064 43857 646066
rect 43791 646061 43857 646064
rect 43119 645384 43185 645387
rect 42336 645382 43185 645384
rect 42336 645326 43124 645382
rect 43180 645326 43185 645382
rect 42336 645324 43185 645326
rect 43119 645321 43185 645324
rect 675759 645384 675825 645387
rect 676090 645384 676096 645386
rect 675759 645382 676096 645384
rect 675759 645326 675764 645382
rect 675820 645326 676096 645382
rect 675759 645324 676096 645326
rect 675759 645321 675825 645324
rect 676090 645322 676096 645324
rect 676160 645322 676166 645386
rect 59247 644940 59313 644943
rect 59247 644938 64416 644940
rect 59247 644882 59252 644938
rect 59308 644882 64416 644938
rect 59247 644880 64416 644882
rect 59247 644877 59313 644880
rect 39810 643907 39870 644466
rect 39810 643902 39921 643907
rect 39810 643846 39860 643902
rect 39916 643846 39921 643902
rect 39810 643844 39921 643846
rect 39855 643841 39921 643844
rect 40002 643167 40062 643726
rect 39951 643162 40062 643167
rect 39951 643106 39956 643162
rect 40012 643106 40062 643162
rect 39951 643104 40062 643106
rect 39951 643101 40017 643104
rect 41538 642427 41598 642838
rect 41487 642422 41598 642427
rect 41487 642366 41492 642422
rect 41548 642366 41598 642422
rect 41487 642364 41598 642366
rect 41487 642361 41553 642364
rect 41730 641687 41790 642172
rect 41679 641682 41790 641687
rect 41679 641626 41684 641682
rect 41740 641626 41790 641682
rect 41679 641624 41790 641626
rect 41679 641621 41745 641624
rect 41922 640799 41982 641358
rect 41871 640794 41982 640799
rect 41871 640738 41876 640794
rect 41932 640738 41982 640794
rect 41871 640736 41982 640738
rect 41871 640733 41937 640736
rect 37314 640059 37374 640544
rect 673978 640290 673984 640354
rect 674048 640352 674054 640354
rect 675375 640352 675441 640355
rect 674048 640350 675441 640352
rect 674048 640294 675380 640350
rect 675436 640294 675441 640350
rect 674048 640292 675441 640294
rect 674048 640290 674054 640292
rect 675375 640289 675441 640292
rect 37314 640054 37425 640059
rect 37314 639998 37364 640054
rect 37420 639998 37425 640054
rect 37314 639996 37425 639998
rect 37359 639993 37425 639996
rect 675898 639846 675904 639910
rect 675968 639846 675974 639910
rect 41346 639467 41406 639730
rect 41295 639462 41406 639467
rect 41295 639406 41300 639462
rect 41356 639406 41406 639462
rect 41295 639404 41406 639406
rect 41295 639401 41361 639404
rect 675706 639402 675712 639466
rect 675776 639464 675782 639466
rect 675906 639464 675966 639846
rect 675776 639404 675966 639464
rect 675776 639402 675782 639404
rect 42682 638946 42688 638948
rect 42336 638886 42688 638946
rect 42682 638884 42688 638886
rect 42752 638884 42758 638948
rect 675514 638662 675520 638726
rect 675584 638724 675590 638726
rect 675584 638664 675774 638724
rect 675584 638662 675590 638664
rect 675471 638578 675537 638579
rect 675471 638574 675520 638578
rect 675584 638576 675590 638578
rect 675471 638518 675476 638574
rect 675471 638514 675520 638518
rect 675584 638516 675628 638576
rect 675584 638514 675590 638516
rect 675471 638513 675537 638514
rect 675714 638135 675774 638664
rect 675714 638130 675825 638135
rect 41922 637691 41982 638102
rect 675714 638074 675764 638130
rect 675820 638074 675825 638130
rect 675714 638072 675825 638074
rect 675759 638069 675825 638072
rect 41922 637686 42033 637691
rect 41922 637630 41972 637686
rect 42028 637630 42033 637686
rect 41922 637628 42033 637630
rect 41967 637625 42033 637628
rect 42114 636803 42174 637362
rect 42063 636798 42174 636803
rect 42063 636742 42068 636798
rect 42124 636742 42174 636798
rect 42063 636740 42174 636742
rect 42063 636737 42129 636740
rect 655311 636652 655377 636655
rect 650208 636650 655377 636652
rect 41538 636359 41598 636622
rect 650208 636594 655316 636650
rect 655372 636594 655377 636650
rect 650208 636592 655377 636594
rect 655311 636589 655377 636592
rect 41538 636354 41649 636359
rect 41538 636298 41588 636354
rect 41644 636298 41649 636354
rect 41538 636296 41649 636298
rect 41583 636293 41649 636296
rect 42114 635619 42174 635734
rect 42114 635614 42225 635619
rect 42114 635558 42164 635614
rect 42220 635558 42225 635614
rect 42114 635556 42225 635558
rect 42159 635553 42225 635556
rect 43023 635024 43089 635027
rect 42336 635022 43089 635024
rect 42336 634966 43028 635022
rect 43084 634966 43089 635022
rect 42336 634964 43089 634966
rect 43023 634961 43089 634964
rect 42306 633544 42366 634106
rect 42447 633544 42513 633547
rect 42306 633542 42513 633544
rect 42306 633486 42452 633542
rect 42508 633486 42513 633542
rect 42306 633484 42513 633486
rect 42447 633481 42513 633484
rect 42306 632360 42366 632626
rect 674511 632508 674577 632511
rect 674511 632506 674814 632508
rect 674511 632450 674516 632506
rect 674572 632450 674814 632506
rect 674511 632448 674814 632450
rect 674511 632445 674577 632448
rect 42447 632360 42513 632363
rect 42306 632358 42513 632360
rect 42306 632302 42452 632358
rect 42508 632302 42513 632358
rect 674754 632330 674814 632448
rect 42306 632300 42513 632302
rect 42447 632297 42513 632300
rect 674511 631768 674577 631771
rect 674511 631766 674814 631768
rect 674511 631710 674516 631766
rect 674572 631710 674814 631766
rect 674511 631708 674814 631710
rect 674511 631705 674577 631708
rect 674754 631442 674814 631708
rect 675759 631028 675825 631031
rect 675759 631026 675966 631028
rect 675759 630970 675764 631026
rect 675820 630970 675966 631026
rect 675759 630968 675966 630970
rect 675759 630965 675825 630968
rect 675759 630882 675825 630883
rect 675906 630882 675966 630968
rect 675706 630880 675712 630882
rect 675668 630820 675712 630880
rect 675776 630878 675825 630882
rect 675820 630822 675825 630878
rect 675706 630818 675712 630820
rect 675776 630818 675825 630822
rect 675898 630818 675904 630882
rect 675968 630818 675974 630882
rect 675759 630817 675825 630818
rect 674127 630732 674193 630735
rect 674127 630730 674784 630732
rect 674127 630674 674132 630730
rect 674188 630674 674784 630730
rect 674127 630672 674784 630674
rect 674127 630669 674193 630672
rect 59535 630584 59601 630587
rect 59535 630582 64416 630584
rect 59535 630526 59540 630582
rect 59596 630526 64416 630582
rect 59535 630524 64416 630526
rect 59535 630521 59601 630524
rect 675759 630438 675825 630439
rect 675706 630374 675712 630438
rect 675776 630436 675825 630438
rect 675776 630434 675868 630436
rect 675820 630378 675868 630434
rect 675776 630376 675868 630378
rect 675776 630374 675825 630376
rect 675759 630373 675825 630374
rect 673263 629844 673329 629847
rect 673263 629842 674784 629844
rect 673263 629786 673268 629842
rect 673324 629786 674784 629842
rect 673263 629784 674784 629786
rect 673263 629781 673329 629784
rect 673839 629104 673905 629107
rect 673839 629102 674784 629104
rect 673839 629046 673844 629102
rect 673900 629046 674784 629102
rect 673839 629044 674784 629046
rect 673839 629041 673905 629044
rect 673743 628364 673809 628367
rect 673743 628362 674784 628364
rect 673743 628306 673748 628362
rect 673804 628306 674784 628362
rect 673743 628304 674784 628306
rect 673743 628301 673809 628304
rect 37359 628216 37425 628219
rect 40762 628216 40768 628218
rect 37359 628214 40768 628216
rect 37359 628158 37364 628214
rect 37420 628158 40768 628214
rect 37359 628156 40768 628158
rect 37359 628153 37425 628156
rect 40762 628154 40768 628156
rect 40832 628154 40838 628218
rect 675375 628068 675441 628071
rect 675330 628066 675441 628068
rect 675330 628010 675380 628066
rect 675436 628010 675441 628066
rect 675330 628005 675441 628010
rect 39951 627920 40017 627923
rect 40570 627920 40576 627922
rect 39951 627918 40576 627920
rect 39951 627862 39956 627918
rect 40012 627862 40576 627918
rect 39951 627860 40576 627862
rect 39951 627857 40017 627860
rect 40570 627858 40576 627860
rect 40640 627858 40646 627922
rect 41295 627774 41361 627775
rect 41295 627772 41344 627774
rect 41252 627770 41344 627772
rect 41252 627714 41300 627770
rect 41252 627712 41344 627714
rect 41295 627710 41344 627712
rect 41408 627710 41414 627774
rect 41583 627772 41649 627775
rect 41722 627772 41728 627774
rect 41583 627770 41728 627772
rect 41583 627714 41588 627770
rect 41644 627714 41728 627770
rect 41583 627712 41728 627714
rect 41295 627709 41361 627710
rect 41583 627709 41649 627712
rect 41722 627710 41728 627712
rect 41792 627710 41798 627774
rect 41914 627562 41920 627626
rect 41984 627624 41990 627626
rect 42159 627624 42225 627627
rect 41984 627622 42225 627624
rect 41984 627566 42164 627622
rect 42220 627566 42225 627622
rect 41984 627564 42225 627566
rect 41984 627562 41990 627564
rect 42159 627561 42225 627564
rect 675330 627520 675390 628005
rect 42063 627478 42129 627479
rect 42063 627476 42112 627478
rect 42020 627474 42112 627476
rect 42020 627418 42068 627474
rect 42020 627416 42112 627418
rect 42063 627414 42112 627416
rect 42176 627414 42182 627478
rect 42063 627413 42129 627414
rect 676282 627266 676288 627330
rect 676352 627266 676358 627330
rect 676290 626706 676350 627266
rect 674415 625922 674481 625925
rect 674415 625920 674784 625922
rect 674415 625864 674420 625920
rect 674476 625864 674784 625920
rect 674415 625862 674784 625864
rect 674415 625859 674481 625862
rect 675898 625638 675904 625702
rect 675968 625638 675974 625702
rect 42682 625046 42688 625110
rect 42752 625108 42758 625110
rect 43311 625108 43377 625111
rect 42752 625106 43377 625108
rect 42752 625050 43316 625106
rect 43372 625050 43377 625106
rect 675906 625078 675966 625638
rect 42752 625048 43377 625050
rect 42752 625046 42758 625048
rect 43311 625045 43377 625048
rect 42298 624898 42304 624962
rect 42368 624898 42374 624962
rect 42306 624812 42366 624898
rect 42490 624812 42496 624814
rect 42306 624752 42496 624812
rect 42490 624750 42496 624752
rect 42560 624750 42566 624814
rect 654351 624812 654417 624815
rect 650208 624810 654417 624812
rect 650208 624754 654356 624810
rect 654412 624754 654417 624810
rect 650208 624752 654417 624754
rect 654351 624749 654417 624752
rect 675706 624750 675712 624814
rect 675776 624750 675782 624814
rect 675714 624264 675774 624750
rect 674607 623776 674673 623779
rect 674607 623774 674814 623776
rect 674607 623718 674612 623774
rect 674668 623718 674814 623774
rect 674607 623716 674814 623718
rect 674607 623713 674673 623716
rect 674754 623598 674814 623716
rect 674319 622740 674385 622743
rect 674319 622738 674784 622740
rect 674319 622682 674324 622738
rect 674380 622682 674784 622738
rect 674319 622680 674784 622682
rect 674319 622677 674385 622680
rect 676474 622086 676480 622150
rect 676544 622086 676550 622150
rect 676482 621970 676542 622086
rect 42063 621706 42129 621707
rect 42063 621702 42112 621706
rect 42176 621704 42182 621706
rect 42063 621646 42068 621702
rect 42063 621642 42112 621646
rect 42176 621644 42220 621704
rect 42176 621642 42182 621644
rect 42063 621641 42129 621642
rect 674170 621050 674176 621114
rect 674240 621112 674246 621114
rect 674240 621052 674784 621112
rect 674240 621050 674246 621052
rect 41967 620818 42033 620819
rect 41914 620754 41920 620818
rect 41984 620816 42033 620818
rect 41984 620814 42076 620816
rect 42028 620758 42076 620814
rect 41984 620756 42076 620758
rect 41984 620754 42033 620756
rect 41967 620753 42033 620754
rect 674362 620310 674368 620374
rect 674432 620372 674438 620374
rect 674432 620312 674784 620372
rect 674432 620310 674438 620312
rect 675375 620076 675441 620079
rect 675330 620074 675441 620076
rect 675330 620018 675380 620074
rect 675436 620018 675441 620074
rect 675330 620013 675441 620018
rect 675330 619454 675390 620013
rect 675130 619126 675136 619190
rect 675200 619126 675206 619190
rect 675138 618862 675198 619126
rect 41530 618238 41536 618302
rect 41600 618300 41606 618302
rect 41775 618300 41841 618303
rect 41600 618298 41841 618300
rect 41600 618242 41780 618298
rect 41836 618242 41841 618298
rect 41600 618240 41841 618242
rect 41600 618238 41606 618240
rect 41775 618237 41841 618240
rect 41967 618154 42033 618155
rect 41914 618090 41920 618154
rect 41984 618152 42033 618154
rect 42490 618152 42496 618154
rect 41984 618150 42496 618152
rect 42028 618094 42496 618150
rect 41984 618092 42496 618094
rect 41984 618090 42033 618092
rect 42490 618090 42496 618092
rect 42560 618090 42566 618154
rect 41967 618089 42033 618090
rect 674415 618004 674481 618007
rect 674415 618002 674784 618004
rect 674415 617946 674420 618002
rect 674476 617946 674784 618002
rect 674415 617944 674784 617946
rect 674415 617941 674481 617944
rect 41775 617858 41841 617859
rect 41722 617856 41728 617858
rect 41684 617796 41728 617856
rect 41792 617854 41841 617858
rect 41836 617798 41841 617854
rect 41722 617794 41728 617796
rect 41792 617794 41841 617798
rect 676858 617794 676864 617858
rect 676928 617794 676934 617858
rect 41775 617793 41841 617794
rect 676866 617234 676926 617794
rect 41338 616462 41344 616526
rect 41408 616524 41414 616526
rect 41775 616524 41841 616527
rect 41408 616522 41841 616524
rect 41408 616466 41780 616522
rect 41836 616466 41841 616522
rect 41408 616464 41841 616466
rect 41408 616462 41414 616464
rect 41775 616461 41841 616464
rect 673071 616376 673137 616379
rect 673071 616374 674784 616376
rect 673071 616318 673076 616374
rect 673132 616318 674784 616374
rect 673071 616316 674784 616318
rect 673071 616313 673137 616316
rect 59535 616228 59601 616231
rect 59535 616226 64416 616228
rect 59535 616170 59540 616226
rect 59596 616170 64416 616226
rect 59535 616168 64416 616170
rect 59535 616165 59601 616168
rect 679746 615047 679806 615606
rect 679695 615042 679806 615047
rect 679695 614986 679700 615042
rect 679756 614986 679806 615042
rect 679695 614984 679806 614986
rect 679695 614981 679761 614984
rect 679695 614452 679761 614455
rect 679695 614450 679806 614452
rect 679695 614394 679700 614450
rect 679756 614394 679806 614450
rect 679695 614389 679806 614394
rect 679746 614052 679806 614389
rect 40762 613354 40768 613418
rect 40832 613416 40838 613418
rect 41775 613416 41841 613419
rect 40832 613414 41841 613416
rect 40832 613358 41780 613414
rect 41836 613358 41841 613414
rect 40832 613356 41841 613358
rect 40832 613354 40838 613356
rect 41775 613353 41841 613356
rect 673978 613354 673984 613418
rect 674048 613416 674054 613418
rect 676282 613416 676288 613418
rect 674048 613356 676288 613416
rect 674048 613354 674054 613356
rect 676282 613354 676288 613356
rect 676352 613354 676358 613418
rect 654351 613120 654417 613123
rect 650208 613118 654417 613120
rect 650208 613062 654356 613118
rect 654412 613062 654417 613118
rect 650208 613060 654417 613062
rect 654351 613057 654417 613060
rect 40570 612762 40576 612826
rect 40640 612824 40646 612826
rect 41775 612824 41841 612827
rect 40640 612822 41841 612824
rect 40640 612766 41780 612822
rect 41836 612766 41841 612822
rect 40640 612764 41841 612766
rect 40640 612762 40646 612764
rect 41775 612761 41841 612764
rect 673978 607730 673984 607794
rect 674048 607792 674054 607794
rect 675375 607792 675441 607795
rect 674048 607790 675441 607792
rect 674048 607734 675380 607790
rect 675436 607734 675441 607790
rect 674048 607732 675441 607734
rect 674048 607730 674054 607732
rect 675375 607729 675441 607732
rect 42735 607718 42801 607721
rect 42336 607716 42801 607718
rect 42336 607660 42740 607716
rect 42796 607660 42801 607716
rect 42336 607658 42801 607660
rect 42735 607655 42801 607658
rect 674362 607138 674368 607202
rect 674432 607200 674438 607202
rect 675471 607200 675537 607203
rect 674432 607198 675537 607200
rect 674432 607142 675476 607198
rect 675532 607142 675537 607198
rect 674432 607140 675537 607142
rect 674432 607138 674438 607140
rect 675471 607137 675537 607140
rect 42735 606904 42801 606907
rect 42336 606902 42801 606904
rect 42336 606846 42740 606902
rect 42796 606846 42801 606902
rect 42336 606844 42801 606846
rect 42735 606841 42801 606844
rect 675663 606462 675729 606463
rect 675663 606458 675712 606462
rect 675776 606460 675782 606462
rect 675663 606402 675668 606458
rect 675663 606398 675712 606402
rect 675776 606400 675820 606460
rect 675776 606398 675782 606400
rect 675663 606397 675729 606398
rect 42159 606312 42225 606315
rect 42114 606310 42225 606312
rect 42114 606254 42164 606310
rect 42220 606254 42225 606310
rect 42114 606249 42225 606254
rect 42114 606060 42174 606249
rect 43503 605276 43569 605279
rect 42336 605274 43569 605276
rect 42336 605218 43508 605274
rect 43564 605218 43569 605274
rect 42336 605216 43569 605218
rect 43503 605213 43569 605216
rect 41914 604918 41920 604982
rect 41984 604980 41990 604982
rect 41984 604918 42030 604980
rect 41970 604832 42030 604918
rect 42106 604832 42112 604834
rect 41970 604772 42112 604832
rect 42106 604770 42112 604772
rect 42176 604770 42182 604834
rect 675130 604770 675136 604834
rect 675200 604832 675206 604834
rect 675375 604832 675441 604835
rect 675200 604830 675441 604832
rect 675200 604774 675380 604830
rect 675436 604774 675441 604830
rect 675200 604772 675441 604774
rect 675200 604770 675206 604772
rect 675375 604769 675441 604772
rect 43215 604684 43281 604687
rect 42306 604682 43281 604684
rect 42306 604626 43220 604682
rect 43276 604626 43281 604682
rect 42306 604624 43281 604626
rect 42306 604432 42366 604624
rect 43215 604621 43281 604624
rect 43599 603796 43665 603799
rect 42336 603794 43665 603796
rect 42336 603738 43604 603794
rect 43660 603738 43665 603794
rect 42336 603736 43665 603738
rect 43599 603733 43665 603736
rect 43407 602908 43473 602911
rect 43791 602908 43857 602911
rect 42336 602906 43857 602908
rect 42336 602850 43412 602906
rect 43468 602850 43796 602906
rect 43852 602850 43857 602906
rect 42336 602848 43857 602850
rect 43407 602845 43473 602848
rect 43791 602845 43857 602848
rect 41538 601875 41598 602138
rect 41538 601870 41649 601875
rect 41538 601814 41588 601870
rect 41644 601814 41649 601870
rect 41538 601812 41649 601814
rect 41583 601809 41649 601812
rect 59535 601872 59601 601875
rect 59535 601870 64416 601872
rect 59535 601814 59540 601870
rect 59596 601814 64416 601870
rect 59535 601812 64416 601814
rect 59535 601809 59601 601812
rect 654447 601428 654513 601431
rect 650208 601426 654513 601428
rect 650208 601370 654452 601426
rect 654508 601370 654513 601426
rect 650208 601368 654513 601370
rect 654447 601365 654513 601368
rect 40002 600691 40062 601250
rect 40002 600686 40113 600691
rect 40002 600630 40052 600686
rect 40108 600630 40113 600686
rect 40002 600628 40113 600630
rect 40047 600625 40113 600628
rect 40962 599950 41022 600510
rect 674170 600182 674176 600246
rect 674240 600244 674246 600246
rect 675471 600244 675537 600247
rect 674240 600242 675537 600244
rect 674240 600186 675476 600242
rect 675532 600186 675537 600242
rect 674240 600184 675537 600186
rect 674240 600182 674246 600184
rect 675471 600181 675537 600184
rect 40954 599886 40960 599950
rect 41024 599886 41030 599950
rect 41922 599211 41982 599622
rect 41871 599206 41982 599211
rect 41871 599150 41876 599206
rect 41932 599150 41982 599206
rect 41871 599148 41982 599150
rect 41871 599145 41937 599148
rect 41346 598471 41406 599030
rect 41346 598466 41457 598471
rect 41346 598410 41396 598466
rect 41452 598410 41457 598466
rect 41346 598408 41457 598410
rect 41391 598405 41457 598408
rect 41922 597583 41982 598142
rect 41922 597578 42033 597583
rect 41922 597522 41972 597578
rect 42028 597522 42033 597578
rect 41922 597520 42033 597522
rect 41967 597517 42033 597520
rect 40770 596842 40830 597402
rect 40762 596778 40768 596842
rect 40832 596778 40838 596842
rect 41538 596251 41598 596514
rect 41487 596246 41598 596251
rect 41487 596190 41492 596246
rect 41548 596190 41598 596246
rect 41487 596188 41598 596190
rect 41487 596185 41553 596188
rect 41730 595215 41790 595774
rect 41730 595210 41841 595215
rect 41730 595154 41780 595210
rect 41836 595154 41841 595210
rect 41730 595152 41841 595154
rect 41775 595149 41841 595152
rect 41154 594474 41214 594886
rect 41146 594410 41152 594474
rect 41216 594410 41222 594474
rect 42306 593732 42366 594220
rect 43066 593732 43072 593734
rect 42306 593672 43072 593732
rect 43066 593670 43072 593672
rect 43136 593670 43142 593734
rect 675898 593522 675904 593586
rect 675968 593584 675974 593586
rect 676666 593584 676672 593586
rect 675968 593524 676672 593584
rect 675968 593522 675974 593524
rect 676666 593522 676672 593524
rect 676736 593522 676742 593586
rect 675759 593436 675825 593439
rect 676858 593436 676864 593438
rect 675759 593434 676864 593436
rect 42114 593143 42174 593406
rect 675759 593378 675764 593434
rect 675820 593378 676864 593434
rect 675759 593376 676864 593378
rect 675759 593373 675825 593376
rect 676858 593374 676864 593376
rect 676928 593374 676934 593438
rect 42063 593138 42174 593143
rect 42063 593082 42068 593138
rect 42124 593082 42174 593138
rect 42063 593080 42174 593082
rect 42063 593077 42129 593080
rect 42114 592403 42174 592592
rect 42114 592398 42225 592403
rect 42114 592342 42164 592398
rect 42220 592342 42225 592398
rect 42114 592340 42225 592342
rect 42159 592337 42225 592340
rect 42831 591808 42897 591811
rect 42336 591806 42897 591808
rect 42336 591750 42836 591806
rect 42892 591750 42897 591806
rect 42336 591748 42897 591750
rect 42831 591745 42897 591748
rect 42306 590476 42366 590964
rect 42735 590476 42801 590479
rect 42306 590474 42801 590476
rect 42306 590418 42740 590474
rect 42796 590418 42801 590474
rect 42306 590416 42801 590418
rect 42735 590413 42801 590416
rect 655119 589588 655185 589591
rect 650208 589586 655185 589588
rect 650208 589530 655124 589586
rect 655180 589530 655185 589586
rect 650208 589528 655185 589530
rect 655119 589525 655185 589528
rect 42735 589440 42801 589443
rect 53775 589440 53841 589443
rect 42336 589438 53841 589440
rect 42336 589382 42740 589438
rect 42796 589382 53780 589438
rect 53836 589382 53841 589438
rect 42336 589380 53841 589382
rect 42735 589377 42801 589380
rect 53775 589377 53841 589380
rect 58191 587516 58257 587519
rect 58191 587514 64416 587516
rect 58191 587458 58196 587514
rect 58252 587458 64416 587514
rect 58191 587456 64416 587458
rect 58191 587453 58257 587456
rect 674607 586776 674673 586779
rect 674754 586776 674814 587042
rect 674607 586774 674814 586776
rect 674607 586718 674612 586774
rect 674668 586718 674814 586774
rect 674607 586716 674814 586718
rect 674607 586713 674673 586716
rect 673839 586332 673905 586335
rect 673839 586330 674784 586332
rect 673839 586274 673844 586330
rect 673900 586274 674784 586330
rect 673839 586272 674784 586274
rect 673839 586269 673905 586272
rect 41338 585974 41344 586038
rect 41408 586036 41414 586038
rect 42106 586036 42112 586038
rect 41408 585976 42112 586036
rect 41408 585974 41414 585976
rect 42106 585974 42112 585976
rect 42176 585974 42182 586038
rect 674415 585444 674481 585447
rect 674415 585442 674784 585444
rect 674415 585386 674420 585442
rect 674476 585386 674784 585442
rect 674415 585384 674784 585386
rect 674415 585381 674481 585384
rect 41583 584852 41649 584855
rect 42490 584852 42496 584854
rect 41583 584850 42496 584852
rect 41583 584794 41588 584850
rect 41644 584794 42496 584850
rect 41583 584792 42496 584794
rect 41583 584789 41649 584792
rect 42490 584790 42496 584792
rect 42560 584790 42566 584854
rect 41487 584704 41553 584707
rect 42298 584704 42304 584706
rect 41487 584702 42304 584704
rect 41487 584646 41492 584702
rect 41548 584646 42304 584702
rect 41487 584644 42304 584646
rect 41487 584641 41553 584644
rect 42298 584642 42304 584644
rect 42368 584642 42374 584706
rect 42735 584704 42801 584707
rect 42874 584704 42880 584706
rect 42735 584702 42880 584704
rect 42735 584646 42740 584702
rect 42796 584646 42880 584702
rect 42735 584644 42880 584646
rect 42735 584641 42801 584644
rect 42874 584642 42880 584644
rect 42944 584642 42950 584706
rect 673839 584704 673905 584707
rect 673839 584702 674784 584704
rect 673839 584646 673844 584702
rect 673900 584646 674784 584702
rect 673839 584644 674784 584646
rect 673839 584641 673905 584644
rect 41391 584556 41457 584559
rect 41722 584556 41728 584558
rect 41391 584554 41728 584556
rect 41391 584498 41396 584554
rect 41452 584498 41728 584554
rect 41391 584496 41728 584498
rect 41391 584493 41457 584496
rect 41722 584494 41728 584496
rect 41792 584494 41798 584558
rect 41871 584410 41937 584411
rect 41871 584408 41920 584410
rect 41828 584406 41920 584408
rect 41828 584350 41876 584406
rect 41828 584348 41920 584350
rect 41871 584346 41920 584348
rect 41984 584346 41990 584410
rect 41871 584345 41937 584346
rect 42063 584262 42129 584263
rect 42063 584260 42112 584262
rect 42020 584258 42112 584260
rect 42020 584202 42068 584258
rect 42020 584200 42112 584202
rect 42063 584198 42112 584200
rect 42176 584198 42182 584262
rect 42063 584197 42129 584198
rect 42682 583754 42688 583818
rect 42752 583816 42758 583818
rect 42831 583816 42897 583819
rect 42752 583814 42897 583816
rect 42752 583758 42836 583814
rect 42892 583758 42897 583814
rect 42752 583756 42897 583758
rect 42752 583754 42758 583756
rect 42831 583753 42897 583756
rect 673839 583816 673905 583819
rect 673839 583814 674784 583816
rect 673839 583758 673844 583814
rect 673900 583758 674784 583814
rect 673839 583756 674784 583758
rect 673839 583753 673905 583756
rect 674607 583372 674673 583375
rect 674607 583370 674814 583372
rect 674607 583314 674612 583370
rect 674668 583314 674814 583370
rect 674607 583312 674814 583314
rect 674607 583309 674673 583312
rect 674754 583194 674814 583312
rect 673263 582336 673329 582339
rect 673263 582334 674784 582336
rect 673263 582278 673268 582334
rect 673324 582278 674784 582334
rect 673263 582276 674784 582278
rect 673263 582273 673329 582276
rect 41967 582042 42033 582043
rect 41914 582040 41920 582042
rect 41876 581980 41920 582040
rect 41984 582038 42033 582042
rect 42028 581982 42033 582038
rect 41914 581978 41920 581980
rect 41984 581978 42033 581982
rect 41967 581977 42033 581978
rect 674938 581682 674944 581746
rect 675008 581682 675014 581746
rect 674946 581566 675006 581682
rect 42927 581448 42993 581451
rect 43066 581448 43072 581450
rect 42927 581446 43072 581448
rect 42927 581390 42932 581446
rect 42988 581390 43072 581446
rect 42927 581388 43072 581390
rect 42927 581385 42993 581388
rect 43066 581386 43072 581388
rect 43136 581386 43142 581450
rect 676474 581238 676480 581302
rect 676544 581238 676550 581302
rect 676482 580678 676542 581238
rect 675322 580350 675328 580414
rect 675392 580350 675398 580414
rect 41146 580202 41152 580266
rect 41216 580264 41222 580266
rect 41775 580264 41841 580267
rect 41216 580262 41841 580264
rect 41216 580206 41780 580262
rect 41836 580206 41841 580262
rect 41216 580204 41841 580206
rect 41216 580202 41222 580204
rect 41775 580201 41841 580204
rect 675330 579864 675390 580350
rect 675898 579610 675904 579674
rect 675968 579610 675974 579674
rect 675906 579050 675966 579610
rect 42159 578932 42225 578935
rect 42682 578932 42688 578934
rect 42159 578930 42688 578932
rect 42159 578874 42164 578930
rect 42220 578874 42688 578930
rect 42159 578872 42688 578874
rect 42159 578869 42225 578872
rect 42682 578870 42688 578872
rect 42752 578870 42758 578934
rect 674170 578870 674176 578934
rect 674240 578932 674246 578934
rect 675898 578932 675904 578934
rect 674240 578872 675904 578932
rect 674240 578870 674246 578872
rect 675898 578870 675904 578872
rect 675968 578870 675974 578934
rect 676282 578722 676288 578786
rect 676352 578722 676358 578786
rect 676290 578384 676350 578722
rect 42927 578342 42993 578343
rect 42874 578340 42880 578342
rect 42836 578280 42880 578340
rect 42944 578338 42993 578342
rect 42988 578282 42993 578338
rect 42874 578278 42880 578280
rect 42944 578278 42993 578282
rect 42927 578277 42993 578278
rect 675514 578130 675520 578194
rect 675584 578130 675590 578194
rect 654447 577896 654513 577899
rect 650208 577894 654513 577896
rect 650208 577838 654452 577894
rect 654508 577838 654513 577894
rect 650208 577836 654513 577838
rect 654447 577833 654513 577836
rect 42490 577538 42496 577602
rect 42560 577600 42566 577602
rect 43023 577600 43089 577603
rect 42560 577598 43089 577600
rect 42560 577542 43028 577598
rect 43084 577542 43089 577598
rect 675522 577570 675582 578130
rect 42560 577540 43089 577542
rect 42560 577538 42566 577540
rect 43023 577537 43089 577540
rect 674554 577242 674560 577306
rect 674624 577304 674630 577306
rect 674624 577244 674814 577304
rect 674624 577242 674630 577244
rect 41775 577010 41841 577011
rect 41722 577008 41728 577010
rect 41684 576948 41728 577008
rect 41792 577006 41841 577010
rect 41836 576950 41841 577006
rect 41722 576946 41728 576948
rect 41792 576946 41841 576950
rect 41775 576945 41841 576946
rect 674754 576756 674814 577244
rect 42298 576354 42304 576418
rect 42368 576416 42374 576418
rect 42447 576416 42513 576419
rect 42368 576414 42513 576416
rect 42368 576358 42452 576414
rect 42508 576358 42513 576414
rect 42368 576356 42513 576358
rect 42368 576354 42374 576356
rect 42447 576353 42513 576356
rect 674746 576058 674752 576122
rect 674816 576058 674822 576122
rect 41338 575910 41344 575974
rect 41408 575972 41414 575974
rect 41775 575972 41841 575975
rect 41914 575972 41920 575974
rect 41408 575970 41920 575972
rect 41408 575914 41780 575970
rect 41836 575914 41920 575970
rect 41408 575912 41920 575914
rect 41408 575910 41414 575912
rect 41775 575909 41841 575912
rect 41914 575910 41920 575912
rect 41984 575910 41990 575974
rect 674754 575942 674814 576058
rect 673359 575232 673425 575235
rect 673359 575230 674814 575232
rect 673359 575174 673364 575230
rect 673420 575174 674814 575230
rect 673359 575172 674814 575174
rect 673359 575169 673425 575172
rect 674754 575128 674814 575172
rect 41530 575022 41536 575086
rect 41600 575084 41606 575086
rect 41775 575084 41841 575087
rect 41600 575082 41841 575084
rect 41600 575026 41780 575082
rect 41836 575026 41841 575082
rect 41600 575024 41841 575026
rect 41600 575022 41606 575024
rect 41775 575021 41841 575024
rect 42159 574642 42225 574643
rect 42106 574640 42112 574642
rect 42068 574580 42112 574640
rect 42176 574638 42225 574642
rect 42220 574582 42225 574638
rect 42106 574578 42112 574580
rect 42176 574578 42225 574582
rect 42159 574577 42225 574578
rect 674415 574344 674481 574347
rect 674415 574342 674784 574344
rect 674415 574286 674420 574342
rect 674476 574286 674784 574342
rect 674415 574284 674784 574286
rect 674415 574281 674481 574284
rect 40762 573986 40768 574050
rect 40832 574048 40838 574050
rect 43119 574048 43185 574051
rect 40832 574046 43185 574048
rect 40832 573990 43124 574046
rect 43180 573990 43185 574046
rect 40832 573988 43185 573990
rect 40832 573986 40838 573988
rect 43119 573985 43185 573988
rect 673839 573604 673905 573607
rect 673839 573602 674784 573604
rect 673839 573546 673844 573602
rect 673900 573546 674784 573602
rect 673839 573544 674784 573546
rect 673839 573541 673905 573544
rect 40954 573098 40960 573162
rect 41024 573160 41030 573162
rect 42447 573160 42513 573163
rect 41024 573158 42513 573160
rect 41024 573102 42452 573158
rect 42508 573102 42513 573158
rect 41024 573100 42513 573102
rect 41024 573098 41030 573100
rect 42447 573097 42513 573100
rect 41914 572950 41920 573014
rect 41984 573012 41990 573014
rect 43066 573012 43072 573014
rect 41984 572952 43072 573012
rect 41984 572950 41990 572952
rect 43066 572950 43072 572952
rect 43136 572950 43142 573014
rect 59535 573012 59601 573015
rect 59535 573010 64416 573012
rect 59535 572954 59540 573010
rect 59596 572954 64416 573010
rect 59535 572952 64416 572954
rect 59535 572949 59601 572952
rect 674415 572864 674481 572867
rect 674415 572862 674784 572864
rect 674415 572806 674420 572862
rect 674476 572806 674784 572862
rect 674415 572804 674784 572806
rect 674415 572801 674481 572804
rect 674415 571976 674481 571979
rect 674415 571974 674784 571976
rect 674415 571918 674420 571974
rect 674476 571918 674784 571974
rect 674415 571916 674784 571918
rect 674415 571913 674481 571916
rect 673839 571236 673905 571239
rect 673839 571234 674784 571236
rect 673839 571178 673844 571234
rect 673900 571178 674784 571234
rect 673839 571176 674784 571178
rect 673839 571173 673905 571176
rect 679746 570203 679806 570318
rect 679746 570198 679857 570203
rect 679746 570142 679796 570198
rect 679852 570142 679857 570198
rect 679746 570140 679857 570142
rect 679791 570137 679857 570140
rect 679791 569312 679857 569315
rect 679746 569310 679857 569312
rect 679746 569254 679796 569310
rect 679852 569254 679857 569310
rect 679746 569249 679857 569254
rect 679746 568838 679806 569249
rect 674895 568722 674961 568723
rect 674895 568720 674944 568722
rect 674852 568718 674944 568720
rect 674852 568662 674900 568718
rect 674852 568660 674944 568662
rect 674895 568658 674944 568660
rect 675008 568658 675014 568722
rect 674895 568657 674961 568658
rect 654351 566204 654417 566207
rect 650208 566202 654417 566204
rect 650208 566146 654356 566202
rect 654412 566146 654417 566202
rect 650208 566144 654417 566146
rect 654351 566141 654417 566144
rect 34479 564724 34545 564727
rect 34434 564722 34545 564724
rect 34434 564666 34484 564722
rect 34540 564666 34545 564722
rect 34434 564661 34545 564666
rect 34434 564472 34494 564661
rect 42114 563543 42174 563658
rect 42114 563538 42225 563543
rect 42114 563482 42164 563538
rect 42220 563482 42225 563538
rect 42114 563480 42225 563482
rect 42159 563477 42225 563480
rect 42831 562874 42897 562877
rect 42336 562872 42897 562874
rect 42336 562816 42836 562872
rect 42892 562816 42897 562872
rect 42336 562814 42897 562816
rect 42831 562811 42897 562814
rect 675322 562442 675328 562506
rect 675392 562504 675398 562506
rect 675471 562504 675537 562507
rect 675392 562502 675537 562504
rect 675392 562446 675476 562502
rect 675532 562446 675537 562502
rect 675392 562444 675537 562446
rect 675392 562442 675398 562444
rect 675471 562441 675537 562444
rect 43215 562060 43281 562063
rect 42336 562058 43281 562060
rect 42336 562002 43220 562058
rect 43276 562002 43281 562058
rect 42336 562000 43281 562002
rect 43215 561997 43281 562000
rect 674170 561998 674176 562062
rect 674240 562060 674246 562062
rect 675471 562060 675537 562063
rect 674240 562058 675537 562060
rect 674240 562002 675476 562058
rect 675532 562002 675537 562058
rect 674240 562000 675537 562002
rect 674240 561998 674246 562000
rect 675471 561997 675537 562000
rect 675471 561766 675537 561767
rect 675471 561762 675520 561766
rect 675584 561764 675590 561766
rect 675471 561706 675476 561762
rect 675471 561702 675520 561706
rect 675584 561704 675628 561764
rect 675584 561702 675590 561704
rect 675471 561701 675537 561702
rect 43503 561616 43569 561619
rect 42306 561614 43569 561616
rect 42306 561558 43508 561614
rect 43564 561558 43569 561614
rect 42306 561556 43569 561558
rect 42306 561216 42366 561556
rect 43503 561553 43569 561556
rect 43599 560580 43665 560583
rect 42336 560578 43665 560580
rect 42336 560522 43604 560578
rect 43660 560522 43665 560578
rect 42336 560520 43665 560522
rect 43599 560517 43665 560520
rect 43407 559840 43473 559843
rect 42306 559838 43473 559840
rect 42306 559782 43412 559838
rect 43468 559782 43473 559838
rect 42306 559780 43473 559782
rect 42306 559736 42366 559780
rect 43407 559777 43473 559780
rect 42927 558952 42993 558955
rect 42336 558950 42993 558952
rect 42336 558894 42932 558950
rect 42988 558894 42993 558950
rect 42336 558892 42993 558894
rect 42927 558889 42993 558892
rect 59439 558952 59505 558955
rect 59439 558950 64416 558952
rect 59439 558894 59444 558950
rect 59500 558894 64416 558950
rect 59439 558892 64416 558894
rect 59439 558889 59505 558892
rect 674938 558890 674944 558954
rect 675008 558952 675014 558954
rect 675008 558892 675774 558952
rect 675008 558890 675014 558892
rect 674938 558742 674944 558806
rect 675008 558804 675014 558806
rect 675471 558804 675537 558807
rect 675008 558802 675537 558804
rect 675008 558746 675476 558802
rect 675532 558746 675537 558802
rect 675008 558744 675537 558746
rect 675714 558804 675774 558892
rect 676282 558804 676288 558806
rect 675714 558744 676288 558804
rect 675008 558742 675014 558744
rect 675471 558741 675537 558744
rect 676282 558742 676288 558744
rect 676352 558742 676358 558806
rect 674554 558150 674560 558214
rect 674624 558212 674630 558214
rect 675375 558212 675441 558215
rect 674624 558210 675441 558212
rect 674624 558154 675380 558210
rect 675436 558154 675441 558210
rect 674624 558152 675441 558154
rect 674624 558150 674630 558152
rect 675375 558149 675441 558152
rect 40194 557475 40254 558034
rect 675759 557620 675825 557623
rect 676858 557620 676864 557622
rect 675759 557618 676864 557620
rect 675759 557562 675764 557618
rect 675820 557562 676864 557618
rect 675759 557560 676864 557562
rect 675759 557557 675825 557560
rect 676858 557558 676864 557560
rect 676928 557558 676934 557622
rect 40194 557470 40305 557475
rect 40194 557414 40244 557470
rect 40300 557414 40305 557470
rect 40194 557412 40305 557414
rect 40239 557409 40305 557412
rect 40770 556734 40830 557294
rect 40762 556670 40768 556734
rect 40832 556670 40838 556734
rect 41730 555995 41790 556406
rect 41391 555994 41457 555995
rect 41338 555930 41344 555994
rect 41408 555992 41457 555994
rect 41408 555990 41500 555992
rect 41452 555934 41500 555990
rect 41408 555932 41500 555934
rect 41679 555990 41790 555995
rect 41679 555934 41684 555990
rect 41740 555934 41790 555990
rect 41679 555932 41790 555934
rect 41408 555930 41457 555932
rect 41391 555929 41457 555930
rect 41679 555929 41745 555932
rect 42114 555255 42174 555814
rect 42114 555250 42225 555255
rect 42114 555194 42164 555250
rect 42220 555194 42225 555250
rect 42114 555192 42225 555194
rect 42159 555189 42225 555192
rect 41922 554367 41982 554926
rect 654447 554512 654513 554515
rect 650208 554510 654513 554512
rect 650208 554454 654452 554510
rect 654508 554454 654513 554510
rect 650208 554452 654513 554454
rect 654447 554449 654513 554452
rect 674746 554450 674752 554514
rect 674816 554512 674822 554514
rect 675375 554512 675441 554515
rect 674816 554510 675441 554512
rect 674816 554454 675380 554510
rect 675436 554454 675441 554510
rect 674816 554452 675441 554454
rect 674816 554450 674822 554452
rect 675375 554449 675441 554452
rect 41922 554362 42033 554367
rect 41922 554306 41972 554362
rect 42028 554306 42033 554362
rect 41922 554304 42033 554306
rect 41967 554301 42033 554304
rect 40962 553626 41022 554186
rect 40954 553562 40960 553626
rect 41024 553562 41030 553626
rect 41730 553035 41790 553298
rect 41391 553034 41457 553035
rect 41338 553032 41344 553034
rect 41300 552972 41344 553032
rect 41408 553030 41457 553034
rect 41452 552974 41457 553030
rect 41338 552970 41344 552972
rect 41408 552970 41457 552974
rect 41730 553030 41841 553035
rect 41730 552974 41780 553030
rect 41836 552974 41841 553030
rect 41730 552972 41841 552974
rect 41391 552969 41457 552970
rect 41775 552969 41841 552972
rect 41538 551999 41598 552558
rect 41538 551994 41649 551999
rect 41538 551938 41588 551994
rect 41644 551938 41649 551994
rect 41538 551936 41649 551938
rect 41583 551933 41649 551936
rect 42306 551256 42366 551670
rect 42447 551404 42513 551407
rect 42447 551402 42750 551404
rect 42447 551346 42452 551402
rect 42508 551346 42750 551402
rect 42447 551344 42750 551346
rect 42447 551341 42513 551344
rect 42447 551256 42513 551259
rect 42306 551254 42513 551256
rect 42306 551198 42452 551254
rect 42508 551198 42513 551254
rect 42306 551196 42513 551198
rect 42447 551193 42513 551196
rect 42690 551108 42750 551344
rect 42336 551048 42750 551108
rect 41922 550072 41982 550190
rect 676474 550158 676480 550222
rect 676544 550158 676550 550222
rect 42063 550072 42129 550075
rect 41922 550070 42129 550072
rect 41922 550014 42068 550070
rect 42124 550014 42129 550070
rect 41922 550012 42129 550014
rect 42063 550009 42129 550012
rect 676482 549924 676542 550158
rect 676666 549924 676672 549926
rect 676482 549864 676672 549924
rect 676666 549862 676672 549864
rect 676736 549862 676742 549926
rect 42306 549332 42366 549376
rect 42927 549332 42993 549335
rect 42306 549330 42993 549332
rect 42306 549274 42932 549330
rect 42988 549274 42993 549330
rect 42306 549272 42993 549274
rect 42927 549269 42993 549272
rect 43023 548592 43089 548595
rect 42336 548590 43089 548592
rect 42336 548534 43028 548590
rect 43084 548534 43089 548590
rect 42336 548532 43089 548534
rect 43023 548529 43089 548532
rect 42306 547704 42366 547748
rect 43311 547704 43377 547707
rect 42306 547702 43377 547704
rect 42306 547646 43316 547702
rect 43372 547646 43377 547702
rect 42306 547644 43377 547646
rect 43311 547641 43377 547644
rect 42306 546224 42366 546268
rect 43311 546224 43377 546227
rect 42306 546222 43377 546224
rect 42306 546166 43316 546222
rect 43372 546166 43377 546222
rect 42306 546164 43377 546166
rect 43311 546161 43377 546164
rect 40570 544830 40576 544894
rect 40640 544892 40646 544894
rect 41338 544892 41344 544894
rect 40640 544832 41344 544892
rect 40640 544830 40646 544832
rect 41338 544830 41344 544832
rect 41408 544830 41414 544894
rect 59535 544448 59601 544451
rect 59535 544446 64416 544448
rect 59535 544390 59540 544446
rect 59596 544390 64416 544446
rect 59535 544388 64416 544390
rect 59535 544385 59601 544388
rect 41007 544152 41073 544155
rect 41146 544152 41152 544154
rect 41007 544150 41152 544152
rect 41007 544094 41012 544150
rect 41068 544094 41152 544150
rect 41007 544092 41152 544094
rect 41007 544089 41073 544092
rect 41146 544090 41152 544092
rect 41216 544090 41222 544154
rect 654159 542672 654225 542675
rect 650208 542670 654225 542672
rect 650208 542614 654164 542670
rect 654220 542614 654225 542670
rect 650208 542612 654225 542614
rect 654159 542609 654225 542612
rect 674319 542080 674385 542083
rect 674319 542078 674784 542080
rect 674319 542022 674324 542078
rect 674380 542022 674784 542078
rect 674319 542020 674784 542022
rect 674319 542017 674385 542020
rect 673935 541488 674001 541491
rect 674415 541488 674481 541491
rect 673935 541486 674481 541488
rect 673935 541430 673940 541486
rect 673996 541430 674420 541486
rect 674476 541430 674481 541486
rect 673935 541428 674481 541430
rect 673935 541425 674001 541428
rect 674415 541425 674481 541428
rect 674607 541488 674673 541491
rect 674607 541486 674814 541488
rect 674607 541430 674612 541486
rect 674668 541430 674814 541486
rect 674607 541428 674814 541430
rect 674607 541425 674673 541428
rect 41338 541278 41344 541342
rect 41408 541340 41414 541342
rect 41487 541340 41553 541343
rect 41408 541338 41553 541340
rect 41408 541282 41492 541338
rect 41548 541282 41553 541338
rect 41408 541280 41553 541282
rect 41408 541278 41414 541280
rect 41487 541277 41553 541280
rect 41679 541340 41745 541343
rect 42298 541340 42304 541342
rect 41679 541338 42304 541340
rect 41679 541282 41684 541338
rect 41740 541282 42304 541338
rect 41679 541280 42304 541282
rect 41679 541277 41745 541280
rect 42298 541278 42304 541280
rect 42368 541278 42374 541342
rect 674754 541310 674814 541428
rect 42447 541192 42513 541195
rect 42874 541192 42880 541194
rect 42447 541190 42880 541192
rect 42447 541134 42452 541190
rect 42508 541134 42880 541190
rect 42447 541132 42880 541134
rect 42447 541129 42513 541132
rect 42874 541130 42880 541132
rect 42944 541130 42950 541194
rect 41871 541046 41937 541047
rect 42159 541046 42225 541047
rect 41871 541044 41920 541046
rect 41828 541042 41920 541044
rect 41828 540986 41876 541042
rect 41828 540984 41920 540986
rect 41871 540982 41920 540984
rect 41984 540982 41990 541046
rect 42106 541044 42112 541046
rect 42068 540984 42112 541044
rect 42176 541042 42225 541046
rect 42220 540986 42225 541042
rect 42106 540982 42112 540984
rect 42176 540982 42225 540986
rect 41871 540981 41937 540982
rect 42159 540981 42225 540982
rect 674607 540748 674673 540751
rect 674607 540746 674814 540748
rect 674607 540690 674612 540746
rect 674668 540690 674814 540746
rect 674607 540688 674814 540690
rect 674607 540685 674673 540688
rect 674754 540422 674814 540688
rect 674607 539860 674673 539863
rect 674607 539858 674814 539860
rect 674607 539802 674612 539858
rect 674668 539802 674814 539858
rect 674607 539800 674814 539802
rect 674607 539797 674673 539800
rect 674754 539682 674814 539800
rect 41146 538910 41152 538974
rect 41216 538972 41222 538974
rect 41871 538972 41937 538975
rect 41216 538970 41937 538972
rect 41216 538914 41876 538970
rect 41932 538914 41937 538970
rect 41216 538912 41937 538914
rect 41216 538910 41222 538912
rect 41871 538909 41937 538912
rect 676674 538679 676734 538794
rect 676674 538674 676785 538679
rect 676674 538618 676724 538674
rect 676780 538618 676785 538674
rect 676674 538616 676785 538618
rect 676719 538613 676785 538616
rect 676482 537643 676542 538128
rect 676482 537638 676593 537643
rect 676482 537582 676532 537638
rect 676588 537582 676593 537638
rect 676482 537580 676593 537582
rect 676527 537577 676593 537580
rect 676674 537051 676734 537314
rect 42063 537050 42129 537051
rect 42063 537048 42112 537050
rect 42020 537046 42112 537048
rect 42020 536990 42068 537046
rect 42020 536988 42112 536990
rect 42063 536986 42112 536988
rect 42176 536986 42182 537050
rect 675706 536986 675712 537050
rect 675776 536986 675782 537050
rect 676623 537046 676734 537051
rect 676623 536990 676628 537046
rect 676684 536990 676734 537046
rect 676623 536988 676734 536990
rect 42063 536985 42129 536986
rect 675714 536500 675774 536986
rect 676623 536985 676689 536988
rect 676282 536246 676288 536310
rect 676352 536246 676358 536310
rect 40570 535654 40576 535718
rect 40640 535716 40646 535718
rect 41530 535716 41536 535718
rect 40640 535656 41536 535716
rect 40640 535654 40646 535656
rect 41530 535654 41536 535656
rect 41600 535654 41606 535718
rect 676290 535686 676350 536246
rect 673978 535358 673984 535422
rect 674048 535420 674054 535422
rect 674048 535360 674814 535420
rect 674048 535358 674054 535360
rect 42159 535272 42225 535275
rect 42874 535272 42880 535274
rect 42159 535270 42880 535272
rect 42159 535214 42164 535270
rect 42220 535214 42880 535270
rect 42159 535212 42880 535214
rect 42159 535209 42225 535212
rect 42874 535210 42880 535212
rect 42944 535210 42950 535274
rect 674754 534872 674814 535360
rect 675130 534618 675136 534682
rect 675200 534618 675206 534682
rect 42298 534470 42304 534534
rect 42368 534532 42374 534534
rect 42927 534532 42993 534535
rect 42368 534530 42993 534532
rect 42368 534474 42932 534530
rect 42988 534474 42993 534530
rect 42368 534472 42993 534474
rect 42368 534470 42374 534472
rect 42927 534469 42993 534472
rect 675138 534058 675198 534618
rect 41967 533794 42033 533795
rect 41914 533730 41920 533794
rect 41984 533792 42033 533794
rect 41984 533790 42076 533792
rect 42028 533734 42076 533790
rect 41984 533732 42076 533734
rect 41984 533730 42033 533732
rect 675898 533730 675904 533794
rect 675968 533730 675974 533794
rect 41967 533729 42033 533730
rect 675906 533392 675966 533730
rect 42159 532758 42225 532759
rect 42106 532756 42112 532758
rect 42032 532696 42112 532756
rect 42176 532756 42225 532758
rect 43066 532756 43072 532758
rect 42176 532754 43072 532756
rect 42220 532698 43072 532754
rect 42106 532694 42112 532696
rect 42176 532696 43072 532698
rect 42176 532694 42225 532696
rect 43066 532694 43072 532696
rect 43136 532694 43142 532758
rect 676666 532694 676672 532758
rect 676736 532694 676742 532758
rect 42159 532693 42225 532694
rect 676674 532578 676734 532694
rect 41530 531806 41536 531870
rect 41600 531868 41606 531870
rect 41775 531868 41841 531871
rect 41600 531866 41841 531868
rect 41600 531810 41780 531866
rect 41836 531810 41841 531866
rect 41600 531808 41841 531810
rect 41600 531806 41606 531808
rect 41775 531805 41841 531808
rect 674362 531658 674368 531722
rect 674432 531720 674438 531722
rect 674432 531660 674784 531720
rect 674432 531658 674438 531660
rect 41338 531362 41344 531426
rect 41408 531424 41414 531426
rect 42447 531424 42513 531427
rect 41408 531422 42513 531424
rect 41408 531366 42452 531422
rect 42508 531366 42513 531422
rect 41408 531364 42513 531366
rect 41408 531362 41414 531364
rect 42447 531361 42513 531364
rect 674799 531128 674865 531131
rect 674754 531126 674865 531128
rect 674754 531070 674804 531126
rect 674860 531070 674865 531126
rect 674754 531065 674865 531070
rect 654063 530980 654129 530983
rect 650208 530978 654129 530980
rect 650208 530922 654068 530978
rect 654124 530922 654129 530978
rect 674754 530950 674814 531065
rect 650208 530920 654129 530922
rect 654063 530917 654129 530920
rect 40954 530030 40960 530094
rect 41024 530092 41030 530094
rect 42927 530092 42993 530095
rect 41024 530090 42993 530092
rect 41024 530034 42932 530090
rect 42988 530034 42993 530090
rect 41024 530032 42993 530034
rect 41024 530030 41030 530032
rect 42927 530029 42993 530032
rect 59535 530092 59601 530095
rect 673071 530092 673137 530095
rect 59535 530090 64416 530092
rect 59535 530034 59540 530090
rect 59596 530034 64416 530090
rect 59535 530032 64416 530034
rect 673071 530090 674784 530092
rect 673071 530034 673076 530090
rect 673132 530034 674784 530090
rect 673071 530032 674784 530034
rect 59535 530029 59601 530032
rect 673071 530029 673137 530032
rect 674799 529500 674865 529503
rect 674754 529498 674865 529500
rect 674754 529442 674804 529498
rect 674860 529442 674865 529498
rect 674754 529437 674865 529442
rect 674754 529322 674814 529437
rect 674799 528908 674865 528911
rect 674754 528906 674865 528908
rect 674754 528850 674804 528906
rect 674860 528850 674865 528906
rect 674754 528845 674865 528850
rect 674754 528582 674814 528845
rect 674799 528020 674865 528023
rect 674754 528018 674865 528020
rect 674754 527962 674804 528018
rect 674860 527962 674865 528018
rect 674754 527957 674865 527962
rect 674754 527842 674814 527957
rect 673551 526984 673617 526987
rect 673551 526982 674784 526984
rect 673551 526926 673556 526982
rect 673612 526926 674784 526982
rect 673551 526924 674784 526926
rect 673551 526921 673617 526924
rect 40762 526478 40768 526542
rect 40832 526540 40838 526542
rect 41775 526540 41841 526543
rect 40832 526538 41841 526540
rect 40832 526482 41780 526538
rect 41836 526482 41841 526538
rect 40832 526480 41841 526482
rect 40832 526478 40838 526480
rect 41775 526477 41841 526480
rect 673167 526244 673233 526247
rect 673167 526242 674784 526244
rect 673167 526186 673172 526242
rect 673228 526186 674784 526242
rect 673167 526184 674784 526186
rect 673167 526181 673233 526184
rect 679746 524767 679806 525326
rect 679746 524762 679857 524767
rect 679746 524706 679796 524762
rect 679852 524706 679857 524762
rect 679746 524704 679857 524706
rect 679791 524701 679857 524704
rect 41583 524174 41649 524175
rect 41530 524172 41536 524174
rect 41492 524112 41536 524172
rect 41600 524170 41649 524174
rect 679791 524172 679857 524175
rect 41644 524114 41649 524170
rect 41530 524110 41536 524112
rect 41600 524110 41649 524114
rect 41583 524109 41649 524110
rect 679746 524170 679857 524172
rect 679746 524114 679796 524170
rect 679852 524114 679857 524170
rect 679746 524109 679857 524114
rect 679746 523846 679806 524109
rect 654063 519288 654129 519291
rect 650208 519286 654129 519288
rect 650208 519230 654068 519286
rect 654124 519230 654129 519286
rect 650208 519228 654129 519230
rect 654063 519225 654129 519228
rect 59535 515736 59601 515739
rect 59535 515734 64416 515736
rect 59535 515678 59540 515734
rect 59596 515678 64416 515734
rect 59535 515676 64416 515678
rect 59535 515673 59601 515676
rect 42159 510114 42225 510115
rect 42106 510050 42112 510114
rect 42176 510112 42225 510114
rect 42176 510110 42268 510112
rect 42220 510054 42268 510110
rect 42176 510052 42268 510054
rect 42176 510050 42225 510052
rect 42159 510049 42225 510050
rect 656367 507448 656433 507451
rect 650208 507446 656433 507448
rect 650208 507390 656372 507446
rect 656428 507390 656433 507446
rect 650208 507388 656433 507390
rect 656367 507385 656433 507388
rect 41583 504044 41649 504047
rect 42159 504046 42225 504047
rect 41722 504044 41728 504046
rect 41583 504042 41728 504044
rect 41583 503986 41588 504042
rect 41644 503986 41728 504042
rect 41583 503984 41728 503986
rect 41583 503981 41649 503984
rect 41722 503982 41728 503984
rect 41792 503982 41798 504046
rect 42106 504044 42112 504046
rect 42068 503984 42112 504044
rect 42176 504042 42225 504046
rect 42220 503986 42225 504042
rect 42106 503982 42112 503984
rect 42176 503982 42225 503986
rect 42159 503981 42225 503982
rect 59535 501232 59601 501235
rect 59535 501230 64416 501232
rect 59535 501174 59540 501230
rect 59596 501174 64416 501230
rect 59535 501172 64416 501174
rect 59535 501169 59601 501172
rect 674754 497831 674814 498094
rect 674703 497826 674814 497831
rect 674703 497770 674708 497826
rect 674764 497770 674814 497826
rect 674703 497768 674814 497770
rect 674703 497765 674769 497768
rect 674415 497310 674481 497313
rect 674415 497308 674784 497310
rect 674415 497252 674420 497308
rect 674476 497252 674784 497308
rect 674415 497250 674784 497252
rect 674415 497247 674481 497250
rect 674415 496496 674481 496499
rect 674415 496494 674784 496496
rect 674415 496438 674420 496494
rect 674476 496438 674784 496494
rect 674415 496436 674784 496438
rect 674415 496433 674481 496436
rect 676719 495904 676785 495907
rect 676674 495902 676785 495904
rect 676674 495846 676724 495902
rect 676780 495846 676785 495902
rect 676674 495841 676785 495846
rect 655215 495756 655281 495759
rect 650208 495754 655281 495756
rect 650208 495698 655220 495754
rect 655276 495698 655281 495754
rect 650208 495696 655281 495698
rect 655215 495693 655281 495696
rect 676674 495578 676734 495841
rect 676674 494575 676734 494838
rect 676674 494570 676785 494575
rect 676674 494514 676724 494570
rect 676780 494514 676785 494570
rect 676674 494512 676785 494514
rect 676719 494509 676785 494512
rect 676482 493983 676542 494098
rect 676482 493978 676593 493983
rect 676482 493922 676532 493978
rect 676588 493922 676593 493978
rect 676482 493920 676593 493922
rect 676527 493917 676593 493920
rect 676674 493095 676734 493358
rect 676623 493090 676734 493095
rect 676623 493034 676628 493090
rect 676684 493034 676734 493090
rect 676623 493032 676734 493034
rect 676623 493029 676689 493032
rect 675514 492734 675520 492798
rect 675584 492734 675590 492798
rect 675522 492470 675582 492734
rect 674511 491908 674577 491911
rect 674511 491906 674814 491908
rect 674511 491850 674516 491906
rect 674572 491850 674814 491906
rect 674511 491848 674814 491850
rect 674511 491845 674577 491848
rect 674754 491730 674814 491848
rect 675322 491402 675328 491466
rect 675392 491402 675398 491466
rect 41775 491022 41841 491023
rect 41722 491020 41728 491022
rect 41684 490960 41728 491020
rect 41792 491018 41841 491022
rect 41836 490962 41841 491018
rect 41722 490958 41728 490960
rect 41792 490958 41841 490962
rect 41775 490957 41841 490958
rect 675330 490842 675390 491402
rect 674991 490280 675057 490283
rect 674946 490278 675057 490280
rect 674946 490222 674996 490278
rect 675052 490222 675057 490278
rect 674946 490217 675057 490222
rect 674946 490102 675006 490217
rect 42106 489626 42112 489690
rect 42176 489626 42182 489690
rect 42114 489392 42174 489626
rect 42298 489392 42304 489394
rect 42114 489332 42304 489392
rect 42298 489330 42304 489332
rect 42368 489330 42374 489394
rect 674319 489392 674385 489395
rect 674319 489390 674784 489392
rect 674319 489334 674324 489390
rect 674380 489334 674784 489390
rect 674319 489332 674784 489334
rect 674319 489329 674385 489332
rect 674607 488800 674673 488803
rect 674607 488798 674814 488800
rect 674607 488742 674612 488798
rect 674668 488742 674814 488798
rect 674607 488740 674814 488742
rect 674607 488737 674673 488740
rect 674754 488622 674814 488740
rect 674170 487702 674176 487766
rect 674240 487764 674246 487766
rect 674240 487704 674784 487764
rect 674240 487702 674246 487704
rect 674938 487406 674944 487470
rect 675008 487406 675014 487470
rect 674946 486920 675006 487406
rect 58575 486876 58641 486879
rect 58575 486874 64416 486876
rect 58575 486818 58580 486874
rect 58636 486818 64416 486874
rect 58575 486816 64416 486818
rect 58575 486813 58641 486816
rect 674554 486666 674560 486730
rect 674624 486728 674630 486730
rect 674624 486668 674814 486728
rect 674624 486666 674630 486668
rect 674754 486106 674814 486668
rect 674895 485544 674961 485547
rect 674895 485542 675006 485544
rect 674895 485486 674900 485542
rect 674956 485486 675006 485542
rect 674895 485481 675006 485486
rect 674946 485292 675006 485481
rect 674223 484656 674289 484659
rect 674223 484654 674784 484656
rect 674223 484598 674228 484654
rect 674284 484598 674784 484654
rect 674223 484596 674784 484598
rect 674223 484593 674289 484596
rect 654255 484064 654321 484067
rect 650208 484062 654321 484064
rect 650208 484006 654260 484062
rect 654316 484006 654321 484062
rect 650208 484004 654321 484006
rect 654255 484001 654321 484004
rect 676858 484002 676864 484066
rect 676928 484002 676934 484066
rect 676866 483812 676926 484002
rect 42298 483706 42304 483770
rect 42368 483768 42374 483770
rect 42682 483768 42688 483770
rect 42368 483708 42688 483768
rect 42368 483706 42374 483708
rect 42682 483706 42688 483708
rect 42752 483706 42758 483770
rect 674746 483558 674752 483622
rect 674816 483558 674822 483622
rect 674754 482998 674814 483558
rect 673743 482288 673809 482291
rect 673743 482286 674814 482288
rect 673743 482230 673748 482286
rect 673804 482230 674814 482286
rect 673743 482228 674814 482230
rect 673743 482225 673809 482228
rect 674754 482184 674814 482228
rect 41775 481104 41841 481107
rect 41914 481104 41920 481106
rect 41775 481102 41920 481104
rect 41775 481046 41780 481102
rect 41836 481046 41920 481102
rect 41775 481044 41920 481046
rect 41775 481041 41841 481044
rect 41914 481042 41920 481044
rect 41984 481042 41990 481106
rect 679746 480811 679806 481370
rect 679746 480806 679857 480811
rect 679746 480750 679796 480806
rect 679852 480750 679857 480806
rect 679746 480748 679857 480750
rect 679791 480745 679857 480748
rect 679791 480068 679857 480071
rect 679746 480066 679857 480068
rect 679746 480010 679796 480066
rect 679852 480010 679857 480066
rect 679746 480005 679857 480010
rect 679746 479890 679806 480005
rect 59535 472520 59601 472523
rect 59535 472518 64416 472520
rect 59535 472462 59540 472518
rect 59596 472462 64416 472518
rect 59535 472460 64416 472462
rect 59535 472457 59601 472460
rect 654447 472224 654513 472227
rect 650208 472222 654513 472224
rect 650208 472166 654452 472222
rect 654508 472166 654513 472222
rect 650208 472164 654513 472166
rect 654447 472161 654513 472164
rect 41914 463936 41920 463938
rect 41730 463876 41920 463936
rect 41730 463790 41790 463876
rect 41914 463874 41920 463876
rect 41984 463874 41990 463938
rect 41722 463726 41728 463790
rect 41792 463726 41798 463790
rect 654447 460532 654513 460535
rect 650208 460530 654513 460532
rect 650208 460474 654452 460530
rect 654508 460474 654513 460530
rect 650208 460472 654513 460474
rect 654447 460469 654513 460472
rect 59535 458164 59601 458167
rect 59535 458162 64416 458164
rect 59535 458106 59540 458162
rect 59596 458106 64416 458162
rect 59535 458104 64416 458106
rect 59535 458101 59601 458104
rect 654351 448840 654417 448843
rect 650208 448838 654417 448840
rect 650208 448782 654356 448838
rect 654412 448782 654417 448838
rect 650208 448780 654417 448782
rect 654351 448777 654417 448780
rect 59535 443808 59601 443811
rect 59535 443806 64416 443808
rect 59535 443750 59540 443806
rect 59596 443750 64416 443806
rect 59535 443748 64416 443750
rect 59535 443745 59601 443748
rect 42255 437148 42321 437151
rect 42255 437146 42366 437148
rect 42255 437090 42260 437146
rect 42316 437090 42366 437146
rect 42255 437085 42366 437090
rect 42306 436896 42366 437085
rect 654447 437000 654513 437003
rect 650208 436998 654513 437000
rect 650208 436942 654452 436998
rect 654508 436942 654513 436998
rect 650208 436940 654513 436942
rect 654447 436937 654513 436940
rect 42255 436260 42321 436263
rect 42255 436258 42366 436260
rect 42255 436202 42260 436258
rect 42316 436202 42366 436258
rect 42255 436197 42366 436202
rect 42306 436082 42366 436197
rect 41871 435520 41937 435523
rect 41871 435518 41982 435520
rect 41871 435462 41876 435518
rect 41932 435462 41982 435518
rect 41871 435457 41982 435462
rect 41922 435194 41982 435457
rect 43311 434484 43377 434487
rect 42336 434482 43377 434484
rect 42336 434426 43316 434482
rect 43372 434426 43377 434482
rect 42336 434424 43377 434426
rect 43311 434421 43377 434424
rect 43215 433596 43281 433599
rect 42336 433594 43281 433596
rect 42336 433538 43220 433594
rect 43276 433538 43281 433594
rect 42336 433536 43281 433538
rect 43215 433533 43281 433536
rect 43599 433004 43665 433007
rect 40416 433002 43665 433004
rect 40416 432974 43604 433002
rect 40386 432946 43604 432974
rect 43660 432946 43665 433002
rect 40386 432944 43665 432946
rect 40386 432710 40446 432944
rect 43599 432941 43665 432944
rect 40378 432646 40384 432710
rect 40448 432646 40454 432710
rect 43407 432116 43473 432119
rect 40608 432114 43473 432116
rect 40608 432086 43412 432114
rect 40578 432058 43412 432086
rect 43468 432058 43473 432114
rect 40578 432056 43473 432058
rect 40578 431970 40638 432056
rect 43407 432053 43473 432056
rect 40570 431906 40576 431970
rect 40640 431906 40646 431970
rect 40770 430786 40830 431346
rect 40762 430722 40768 430786
rect 40832 430722 40838 430786
rect 41922 429899 41982 430458
rect 41922 429894 42033 429899
rect 41922 429838 41972 429894
rect 42028 429838 42033 429894
rect 41922 429836 42033 429838
rect 41967 429833 42033 429836
rect 40962 429454 41022 429718
rect 40954 429390 40960 429454
rect 41024 429390 41030 429454
rect 59535 429452 59601 429455
rect 59535 429450 64416 429452
rect 59535 429394 59540 429450
rect 59596 429394 64416 429450
rect 59535 429392 64416 429394
rect 59535 429389 59601 429392
rect 41346 428418 41406 428830
rect 41338 428354 41344 428418
rect 41408 428354 41414 428418
rect 42114 427678 42174 428238
rect 42106 427614 42112 427678
rect 42176 427614 42182 427678
rect 41730 426939 41790 427350
rect 41730 426934 41841 426939
rect 41730 426878 41780 426934
rect 41836 426878 41841 426934
rect 41730 426876 41841 426878
rect 41775 426873 41841 426876
rect 41154 426346 41214 426536
rect 41146 426282 41152 426346
rect 41216 426282 41222 426346
rect 41538 425162 41598 425722
rect 654447 425456 654513 425459
rect 650208 425454 654513 425456
rect 650208 425398 654452 425454
rect 654508 425398 654513 425454
rect 650208 425396 654513 425398
rect 654447 425393 654513 425396
rect 41530 425098 41536 425162
rect 41600 425098 41606 425162
rect 42306 424420 42366 424908
rect 42543 424420 42609 424423
rect 42306 424418 42609 424420
rect 42306 424362 42548 424418
rect 42604 424362 42609 424418
rect 42306 424360 42609 424362
rect 42543 424357 42609 424360
rect 37314 423683 37374 424094
rect 37314 423678 37425 423683
rect 37314 423622 37364 423678
rect 37420 423622 37425 423678
rect 37314 423620 37425 423622
rect 37359 423617 37425 423620
rect 40194 423239 40254 423428
rect 40143 423234 40254 423239
rect 40143 423178 40148 423234
rect 40204 423178 40254 423234
rect 40143 423176 40254 423178
rect 40143 423173 40209 423176
rect 42106 423174 42112 423238
rect 42176 423174 42182 423238
rect 42114 423090 42174 423174
rect 42106 423026 42112 423090
rect 42176 423026 42182 423090
rect 37314 422055 37374 422614
rect 37263 422050 37374 422055
rect 37263 421994 37268 422050
rect 37324 421994 37374 422050
rect 37263 421992 37374 421994
rect 37263 421989 37329 421992
rect 40194 421315 40254 421800
rect 40194 421310 40305 421315
rect 40194 421254 40244 421310
rect 40300 421254 40305 421310
rect 40194 421252 40305 421254
rect 40239 421249 40305 421252
rect 43119 421016 43185 421019
rect 42336 421014 43185 421016
rect 42336 420958 43124 421014
rect 43180 420958 43185 421014
rect 42336 420956 43185 420958
rect 43119 420953 43185 420956
rect 42306 419983 42366 420098
rect 42306 419978 42417 419983
rect 42306 419922 42356 419978
rect 42412 419922 42417 419978
rect 42306 419920 42417 419922
rect 42351 419917 42417 419920
rect 42306 418503 42366 418618
rect 42306 418498 42417 418503
rect 42306 418442 42356 418498
rect 42412 418442 42417 418498
rect 42306 418440 42417 418442
rect 42351 418437 42417 418440
rect 58383 415096 58449 415099
rect 58383 415094 64416 415096
rect 58383 415038 58388 415094
rect 58444 415038 64416 415094
rect 58383 415036 64416 415038
rect 58383 415033 58449 415036
rect 653871 413616 653937 413619
rect 650208 413614 653937 413616
rect 650208 413558 653876 413614
rect 653932 413558 653937 413614
rect 650208 413556 653937 413558
rect 653871 413553 653937 413556
rect 676527 412138 676593 412139
rect 676474 412136 676480 412138
rect 676436 412076 676480 412136
rect 676544 412134 676593 412138
rect 676588 412078 676593 412134
rect 676474 412074 676480 412076
rect 676544 412074 676593 412078
rect 676527 412073 676593 412074
rect 676623 411990 676689 411991
rect 676623 411986 676672 411990
rect 676736 411988 676742 411990
rect 676623 411930 676628 411986
rect 676623 411926 676672 411930
rect 676736 411928 676780 411988
rect 676736 411926 676742 411928
rect 676623 411925 676689 411926
rect 674754 409327 674814 409886
rect 674703 409322 674814 409327
rect 674703 409266 674708 409322
rect 674764 409266 674814 409322
rect 674703 409264 674814 409266
rect 674703 409261 674769 409264
rect 42298 409114 42304 409178
rect 42368 409176 42374 409178
rect 42368 409116 42558 409176
rect 42368 409114 42374 409116
rect 42498 408882 42558 409116
rect 674415 409102 674481 409105
rect 674415 409100 674784 409102
rect 674415 409044 674420 409100
rect 674476 409044 674784 409100
rect 674415 409042 674784 409044
rect 674415 409039 674481 409042
rect 42490 408818 42496 408882
rect 42560 408818 42566 408882
rect 674703 408436 674769 408439
rect 674703 408434 674814 408436
rect 674703 408378 674708 408434
rect 674764 408378 674814 408434
rect 674703 408373 674814 408378
rect 674754 408258 674814 408373
rect 676719 407696 676785 407699
rect 676674 407694 676785 407696
rect 676674 407638 676724 407694
rect 676780 407638 676785 407694
rect 676674 407633 676785 407638
rect 676674 407444 676734 407633
rect 673839 406660 673905 406663
rect 673839 406658 674784 406660
rect 673839 406602 673844 406658
rect 673900 406602 674784 406658
rect 673839 406600 674784 406602
rect 673839 406597 673905 406600
rect 42063 406366 42129 406367
rect 42063 406362 42112 406366
rect 42176 406364 42182 406366
rect 42063 406306 42068 406362
rect 42063 406302 42112 406306
rect 42176 406304 42220 406364
rect 42176 406302 42182 406304
rect 42063 406301 42129 406302
rect 676474 406154 676480 406218
rect 676544 406154 676550 406218
rect 674170 405858 674176 405922
rect 674240 405920 674246 405922
rect 676482 405920 676542 406154
rect 674240 405890 676542 405920
rect 674240 405860 676512 405890
rect 674240 405858 674246 405860
rect 675322 405266 675328 405330
rect 675392 405328 675398 405330
rect 676666 405328 676672 405330
rect 675392 405268 676672 405328
rect 675392 405266 675398 405268
rect 676666 405266 676672 405268
rect 676736 405266 676742 405330
rect 42159 405180 42225 405183
rect 42490 405180 42496 405182
rect 42159 405178 42496 405180
rect 42159 405122 42164 405178
rect 42220 405122 42496 405178
rect 42159 405120 42496 405122
rect 42159 405117 42225 405120
rect 42490 405118 42496 405120
rect 42560 405118 42566 405182
rect 676674 405150 676734 405266
rect 674031 404292 674097 404295
rect 674031 404290 674784 404292
rect 674031 404234 674036 404290
rect 674092 404234 674784 404290
rect 674031 404232 674784 404234
rect 674031 404229 674097 404232
rect 41775 403702 41841 403703
rect 41722 403638 41728 403702
rect 41792 403700 41841 403702
rect 41792 403698 41884 403700
rect 41836 403642 41884 403698
rect 41792 403640 41884 403642
rect 41792 403638 41841 403640
rect 41775 403637 41841 403638
rect 41914 403194 41920 403258
rect 41984 403256 41990 403258
rect 42255 403256 42321 403259
rect 41984 403254 42321 403256
rect 41984 403198 42260 403254
rect 42316 403198 42321 403254
rect 41984 403196 42321 403198
rect 41984 403194 41990 403196
rect 42255 403193 42321 403196
rect 43503 403256 43569 403259
rect 43695 403256 43761 403259
rect 674946 403258 675006 403522
rect 43503 403254 43761 403256
rect 43503 403198 43508 403254
rect 43564 403198 43700 403254
rect 43756 403198 43761 403254
rect 43503 403196 43761 403198
rect 43503 403193 43569 403196
rect 43695 403193 43761 403196
rect 674938 403194 674944 403258
rect 675008 403194 675014 403258
rect 41530 402602 41536 402666
rect 41600 402664 41606 402666
rect 41775 402664 41841 402667
rect 41600 402662 41841 402664
rect 41600 402606 41780 402662
rect 41836 402606 41841 402662
rect 41600 402604 41841 402606
rect 41600 402602 41606 402604
rect 41775 402601 41841 402604
rect 675330 402075 675390 402634
rect 675330 402070 675441 402075
rect 675330 402014 675380 402070
rect 675436 402014 675441 402070
rect 675330 402012 675441 402014
rect 675375 402009 675441 402012
rect 41338 401862 41344 401926
rect 41408 401924 41414 401926
rect 41775 401924 41841 401927
rect 41408 401922 41841 401924
rect 41408 401866 41780 401922
rect 41836 401866 41841 401922
rect 41408 401864 41841 401866
rect 41408 401862 41414 401864
rect 41775 401861 41841 401864
rect 673935 401924 674001 401927
rect 673935 401922 674784 401924
rect 673935 401866 673940 401922
rect 673996 401866 674784 401922
rect 673935 401864 674784 401866
rect 673935 401861 674001 401864
rect 654447 401776 654513 401779
rect 650208 401774 654513 401776
rect 650208 401718 654452 401774
rect 654508 401718 654513 401774
rect 650208 401716 654513 401718
rect 654447 401713 654513 401716
rect 57615 400740 57681 400743
rect 57615 400738 64416 400740
rect 57615 400682 57620 400738
rect 57676 400682 64416 400738
rect 57615 400680 64416 400682
rect 57615 400677 57681 400680
rect 674554 400530 674560 400594
rect 674624 400592 674630 400594
rect 674754 400592 674814 401154
rect 674624 400532 674814 400592
rect 674624 400530 674630 400532
rect 674362 400382 674368 400446
rect 674432 400444 674438 400446
rect 674432 400384 674784 400444
rect 674432 400382 674438 400384
rect 40762 400086 40768 400150
rect 40832 400148 40838 400150
rect 41775 400148 41841 400151
rect 40832 400146 41841 400148
rect 40832 400090 41780 400146
rect 41836 400090 41841 400146
rect 40832 400088 41841 400090
rect 40832 400086 40838 400088
rect 41775 400085 41841 400088
rect 41146 399494 41152 399558
rect 41216 399556 41222 399558
rect 41775 399556 41841 399559
rect 41216 399554 41841 399556
rect 41216 399498 41780 399554
rect 41836 399498 41841 399554
rect 41216 399496 41841 399498
rect 41216 399494 41222 399496
rect 41775 399493 41841 399496
rect 675138 399411 675198 399526
rect 675138 399406 675249 399411
rect 675138 399350 675188 399406
rect 675244 399350 675249 399406
rect 675138 399348 675249 399350
rect 675183 399345 675249 399348
rect 40954 398754 40960 398818
rect 41024 398816 41030 398818
rect 41775 398816 41841 398819
rect 41024 398814 41841 398816
rect 41024 398758 41780 398814
rect 41836 398758 41841 398814
rect 41024 398756 41841 398758
rect 41024 398754 41030 398756
rect 41775 398753 41841 398756
rect 674607 398520 674673 398523
rect 674754 398520 674814 398786
rect 674607 398518 674814 398520
rect 674607 398462 674612 398518
rect 674668 398462 674814 398518
rect 674607 398460 674814 398462
rect 674607 398457 674673 398460
rect 674319 397928 674385 397931
rect 674319 397926 674784 397928
rect 674319 397870 674324 397926
rect 674380 397870 674784 397926
rect 674319 397868 674784 397870
rect 674319 397865 674385 397868
rect 674127 397188 674193 397191
rect 674127 397186 674784 397188
rect 674127 397130 674132 397186
rect 674188 397130 674784 397186
rect 674127 397128 674784 397130
rect 674127 397125 674193 397128
rect 674946 396155 675006 396418
rect 674895 396150 675006 396155
rect 674895 396094 674900 396150
rect 674956 396094 675006 396150
rect 674895 396092 675006 396094
rect 674895 396089 674961 396092
rect 675138 395415 675198 395604
rect 675087 395410 675198 395415
rect 675087 395354 675092 395410
rect 675148 395354 675198 395410
rect 675087 395352 675198 395354
rect 675087 395349 675153 395352
rect 674946 394527 675006 394790
rect 674946 394522 675057 394527
rect 674946 394466 674996 394522
rect 675052 394466 675057 394522
rect 674946 394464 675057 394466
rect 674991 394461 675057 394464
rect 42351 393932 42417 393935
rect 42306 393930 42417 393932
rect 42306 393874 42356 393930
rect 42412 393874 42417 393930
rect 42306 393869 42417 393874
rect 42306 393680 42366 393869
rect 674754 393787 674814 393976
rect 674703 393782 674814 393787
rect 674703 393726 674708 393782
rect 674764 393726 674814 393782
rect 674703 393724 674814 393726
rect 674703 393721 674769 393724
rect 42639 392896 42705 392899
rect 42336 392894 42705 392896
rect 42336 392838 42644 392894
rect 42700 392838 42705 392894
rect 42336 392836 42705 392838
rect 42639 392833 42705 392836
rect 679746 392603 679806 393162
rect 679695 392598 679806 392603
rect 679695 392542 679700 392598
rect 679756 392542 679806 392598
rect 679695 392540 679806 392542
rect 679695 392537 679761 392540
rect 42351 392304 42417 392307
rect 42306 392302 42417 392304
rect 42306 392246 42356 392302
rect 42412 392246 42417 392302
rect 42306 392241 42417 392246
rect 42306 392052 42366 392241
rect 679695 392156 679761 392159
rect 679695 392154 679806 392156
rect 679695 392098 679700 392154
rect 679756 392098 679806 392154
rect 679695 392093 679806 392098
rect 679746 391682 679806 392093
rect 43215 391268 43281 391271
rect 42336 391266 43281 391268
rect 42336 391210 43220 391266
rect 43276 391210 43281 391266
rect 42336 391208 43281 391210
rect 43215 391205 43281 391208
rect 43503 390972 43569 390975
rect 42306 390970 43569 390972
rect 42306 390914 43508 390970
rect 43564 390914 43569 390970
rect 42306 390912 43569 390914
rect 42306 390424 42366 390912
rect 43503 390909 43569 390912
rect 40378 390170 40384 390234
rect 40448 390170 40454 390234
rect 40386 389758 40446 390170
rect 654447 390084 654513 390087
rect 650208 390082 654513 390084
rect 650208 390026 654452 390082
rect 654508 390026 654513 390082
rect 650208 390024 654513 390026
rect 654447 390021 654513 390024
rect 40570 389134 40576 389198
rect 40640 389134 40646 389198
rect 40578 388870 40638 389134
rect 40770 387570 40830 388130
rect 40762 387506 40768 387570
rect 40832 387506 40838 387570
rect 41922 386683 41982 387242
rect 41922 386678 42033 386683
rect 41922 386622 41972 386678
rect 42028 386622 42033 386678
rect 41922 386620 42033 386622
rect 41967 386617 42033 386620
rect 40962 386090 41022 386502
rect 59247 386384 59313 386387
rect 59247 386382 64416 386384
rect 59247 386326 59252 386382
rect 59308 386326 64416 386382
rect 59247 386324 64416 386326
rect 59247 386321 59313 386324
rect 40954 386026 40960 386090
rect 41024 386026 41030 386090
rect 41346 385202 41406 385614
rect 41338 385138 41344 385202
rect 41408 385138 41414 385202
rect 42114 384462 42174 385022
rect 42106 384398 42112 384462
rect 42176 384398 42182 384462
rect 42306 383575 42366 384134
rect 42306 383570 42417 383575
rect 42306 383514 42356 383570
rect 42412 383514 42417 383570
rect 42306 383512 42417 383514
rect 42351 383509 42417 383512
rect 41154 383130 41214 383394
rect 41146 383066 41152 383130
rect 41216 383066 41222 383130
rect 41538 381946 41598 382506
rect 41530 381882 41536 381946
rect 41600 381882 41606 381946
rect 37314 381207 37374 381766
rect 37263 381202 37374 381207
rect 37263 381146 37268 381202
rect 37324 381146 37374 381202
rect 37263 381144 37374 381146
rect 37263 381141 37329 381144
rect 40194 380467 40254 380878
rect 40143 380462 40254 380467
rect 40143 380406 40148 380462
rect 40204 380406 40254 380462
rect 40143 380404 40254 380406
rect 40143 380401 40209 380404
rect 40002 380023 40062 380212
rect 40002 380018 40113 380023
rect 40002 379962 40052 380018
rect 40108 379962 40113 380018
rect 40002 379960 40113 379962
rect 40047 379957 40113 379960
rect 37314 378839 37374 379398
rect 37314 378834 37425 378839
rect 37314 378778 37364 378834
rect 37420 378778 37425 378834
rect 37314 378776 37425 378778
rect 37359 378773 37425 378776
rect 674554 378774 674560 378838
rect 674624 378836 674630 378838
rect 675471 378836 675537 378839
rect 674624 378834 675537 378836
rect 674624 378778 675476 378834
rect 675532 378778 675537 378834
rect 674624 378776 675537 378778
rect 674624 378774 674630 378776
rect 675471 378773 675537 378776
rect 40194 378099 40254 378584
rect 654447 378540 654513 378543
rect 650208 378538 654513 378540
rect 650208 378482 654452 378538
rect 654508 378482 654513 378538
rect 650208 378480 654513 378482
rect 654447 378477 654513 378480
rect 40194 378094 40305 378099
rect 40194 378038 40244 378094
rect 40300 378038 40305 378094
rect 40194 378036 40305 378038
rect 40239 378033 40305 378036
rect 43119 377800 43185 377803
rect 42336 377798 43185 377800
rect 42336 377742 43124 377798
rect 43180 377742 43185 377798
rect 42336 377740 43185 377742
rect 43119 377737 43185 377740
rect 42306 376619 42366 376956
rect 42255 376614 42366 376619
rect 42255 376558 42260 376614
rect 42316 376558 42366 376614
rect 42255 376556 42366 376558
rect 42255 376553 42321 376556
rect 42306 375287 42366 375402
rect 42255 375282 42366 375287
rect 42255 375226 42260 375282
rect 42316 375226 42366 375282
rect 42255 375224 42366 375226
rect 42255 375221 42321 375224
rect 675183 374544 675249 374547
rect 675514 374544 675520 374546
rect 675183 374542 675520 374544
rect 675183 374486 675188 374542
rect 675244 374486 675520 374542
rect 675183 374484 675520 374486
rect 675183 374481 675249 374484
rect 675514 374482 675520 374484
rect 675584 374482 675590 374546
rect 675087 374100 675153 374103
rect 675706 374100 675712 374102
rect 675087 374098 675712 374100
rect 675087 374042 675092 374098
rect 675148 374042 675712 374098
rect 675087 374040 675712 374042
rect 675087 374037 675153 374040
rect 675706 374038 675712 374040
rect 675776 374038 675782 374102
rect 674938 373890 674944 373954
rect 675008 373952 675014 373954
rect 675471 373952 675537 373955
rect 675008 373950 675537 373952
rect 675008 373894 675476 373950
rect 675532 373894 675537 373950
rect 675008 373892 675537 373894
rect 675008 373890 675014 373892
rect 675471 373889 675537 373892
rect 674362 371966 674368 372030
rect 674432 372028 674438 372030
rect 675375 372028 675441 372031
rect 674432 372026 675441 372028
rect 674432 371970 675380 372026
rect 675436 371970 675441 372026
rect 674432 371968 675441 371970
rect 674432 371966 674438 371968
rect 675375 371965 675441 371968
rect 59535 371880 59601 371883
rect 59535 371878 64416 371880
rect 59535 371822 59540 371878
rect 59596 371822 64416 371878
rect 59535 371820 64416 371822
rect 59535 371817 59601 371820
rect 38319 370548 38385 370551
rect 42298 370548 42304 370550
rect 38319 370546 42304 370548
rect 38319 370490 38324 370546
rect 38380 370490 42304 370546
rect 38319 370488 42304 370490
rect 38319 370485 38385 370488
rect 42298 370486 42304 370488
rect 42368 370486 42374 370550
rect 654447 366552 654513 366555
rect 650208 366550 654513 366552
rect 650208 366494 654452 366550
rect 654508 366494 654513 366550
rect 650208 366492 654513 366494
rect 654447 366489 654513 366492
rect 674703 364924 674769 364927
rect 674703 364922 674814 364924
rect 674703 364866 674708 364922
rect 674764 364866 674814 364922
rect 674703 364861 674814 364866
rect 674754 364672 674814 364861
rect 674415 363888 674481 363891
rect 674415 363886 674784 363888
rect 674415 363830 674420 363886
rect 674476 363830 674784 363886
rect 674415 363828 674784 363830
rect 674415 363825 674481 363828
rect 674703 363296 674769 363299
rect 674703 363294 674814 363296
rect 674703 363238 674708 363294
rect 674764 363238 674814 363294
rect 674703 363233 674814 363238
rect 674754 363044 674814 363233
rect 42063 362854 42129 362855
rect 42063 362850 42112 362854
rect 42176 362852 42182 362854
rect 42063 362794 42068 362850
rect 42063 362790 42112 362794
rect 42176 362792 42220 362852
rect 42176 362790 42182 362792
rect 42063 362789 42129 362790
rect 673839 362260 673905 362263
rect 673839 362258 674784 362260
rect 673839 362202 673844 362258
rect 673900 362202 674784 362258
rect 673839 362200 674784 362202
rect 673839 362197 673905 362200
rect 41871 361966 41937 361967
rect 41871 361964 41920 361966
rect 41828 361962 41920 361964
rect 41828 361906 41876 361962
rect 41828 361904 41920 361906
rect 41871 361902 41920 361904
rect 41984 361902 41990 361966
rect 41871 361901 41937 361902
rect 674362 361384 674368 361448
rect 674432 361446 674438 361448
rect 674432 361386 674784 361446
rect 674432 361384 674438 361386
rect 674170 360718 674176 360782
rect 674240 360780 674246 360782
rect 674240 360720 674784 360780
rect 674240 360718 674246 360720
rect 41775 360634 41841 360635
rect 41722 360570 41728 360634
rect 41792 360632 41841 360634
rect 41792 360630 41884 360632
rect 41836 360574 41884 360630
rect 41792 360572 41884 360574
rect 41792 360570 41841 360572
rect 41775 360569 41841 360570
rect 42255 360190 42321 360191
rect 42255 360186 42304 360190
rect 42368 360188 42374 360190
rect 42255 360130 42260 360186
rect 42255 360126 42304 360130
rect 42368 360128 42412 360188
rect 42368 360126 42374 360128
rect 675322 360126 675328 360190
rect 675392 360126 675398 360190
rect 42255 360125 42321 360126
rect 673978 359978 673984 360042
rect 674048 360040 674054 360042
rect 675330 360040 675390 360126
rect 674048 359980 675390 360040
rect 674048 359978 674054 359980
rect 675330 359936 675390 359980
rect 41530 359386 41536 359450
rect 41600 359448 41606 359450
rect 41775 359448 41841 359451
rect 41600 359446 41841 359448
rect 41600 359390 41780 359446
rect 41836 359390 41841 359446
rect 41600 359388 41841 359390
rect 41600 359386 41606 359388
rect 41775 359385 41841 359388
rect 673935 359152 674001 359155
rect 673935 359150 674784 359152
rect 673935 359094 673940 359150
rect 673996 359094 674784 359150
rect 673935 359092 674784 359094
rect 673935 359089 674001 359092
rect 41338 358646 41344 358710
rect 41408 358708 41414 358710
rect 41775 358708 41841 358711
rect 41408 358706 41841 358708
rect 41408 358650 41780 358706
rect 41836 358650 41841 358706
rect 41408 358648 41841 358650
rect 41408 358646 41414 358648
rect 41775 358645 41841 358648
rect 677058 358119 677118 358234
rect 677058 358114 677169 358119
rect 677058 358058 677108 358114
rect 677164 358058 677169 358114
rect 677058 358056 677169 358058
rect 677103 358053 677169 358056
rect 60207 357672 60273 357675
rect 60207 357670 64416 357672
rect 60207 357614 60212 357670
rect 60268 357614 64416 357670
rect 60207 357612 64416 357614
rect 60207 357609 60273 357612
rect 674607 357228 674673 357231
rect 674754 357228 674814 357494
rect 674607 357226 674814 357228
rect 674607 357170 674612 357226
rect 674668 357170 674814 357226
rect 674607 357168 674814 357170
rect 674607 357165 674673 357168
rect 40762 356870 40768 356934
rect 40832 356932 40838 356934
rect 41775 356932 41841 356935
rect 40832 356930 41841 356932
rect 40832 356874 41780 356930
rect 41836 356874 41841 356930
rect 40832 356872 41841 356874
rect 40832 356870 40838 356872
rect 41775 356869 41841 356872
rect 675138 356491 675198 356606
rect 41146 356426 41152 356490
rect 41216 356488 41222 356490
rect 41775 356488 41841 356491
rect 41216 356486 41841 356488
rect 41216 356430 41780 356486
rect 41836 356430 41841 356486
rect 41216 356428 41841 356430
rect 675138 356486 675249 356491
rect 675138 356430 675188 356486
rect 675244 356430 675249 356486
rect 675138 356428 675249 356430
rect 41216 356426 41222 356428
rect 41775 356425 41841 356428
rect 675183 356425 675249 356428
rect 676866 355751 676926 356014
rect 676866 355746 676977 355751
rect 676866 355690 676916 355746
rect 676972 355690 676977 355746
rect 676866 355688 676977 355690
rect 676911 355685 676977 355688
rect 40954 355538 40960 355602
rect 41024 355600 41030 355602
rect 41775 355600 41841 355603
rect 41024 355598 41841 355600
rect 41024 355542 41780 355598
rect 41836 355542 41841 355598
rect 41024 355540 41841 355542
rect 41024 355538 41030 355540
rect 41775 355537 41841 355540
rect 677058 355011 677118 355126
rect 677007 355006 677118 355011
rect 677007 354950 677012 355006
rect 677068 354950 677118 355006
rect 677007 354948 677118 354950
rect 677007 354945 677073 354948
rect 655311 354860 655377 354863
rect 650208 354858 655377 354860
rect 650208 354802 655316 354858
rect 655372 354802 655377 354858
rect 650208 354800 655377 354802
rect 655311 354797 655377 354800
rect 675330 354123 675390 354386
rect 675279 354118 675390 354123
rect 675279 354062 675284 354118
rect 675340 354062 675390 354118
rect 675279 354060 675390 354062
rect 675279 354057 675345 354060
rect 675138 353383 675198 353498
rect 675087 353378 675198 353383
rect 675087 353322 675092 353378
rect 675148 353322 675198 353378
rect 675087 353320 675198 353322
rect 675087 353317 675153 353320
rect 674319 352788 674385 352791
rect 674319 352786 674784 352788
rect 674319 352730 674324 352786
rect 674380 352730 674784 352786
rect 674319 352728 674784 352730
rect 674319 352725 674385 352728
rect 676866 351755 676926 351870
rect 676815 351750 676926 351755
rect 676815 351694 676820 351750
rect 676876 351694 676926 351750
rect 676815 351692 676926 351694
rect 676815 351689 676881 351692
rect 674223 351308 674289 351311
rect 674223 351306 674784 351308
rect 674223 351250 674228 351306
rect 674284 351250 674784 351306
rect 674223 351248 674784 351250
rect 674223 351245 674289 351248
rect 42351 350716 42417 350719
rect 42306 350714 42417 350716
rect 42306 350658 42356 350714
rect 42412 350658 42417 350714
rect 42306 350653 42417 350658
rect 42306 350538 42366 350653
rect 674754 350275 674814 350390
rect 674754 350270 674865 350275
rect 674754 350214 674804 350270
rect 674860 350214 674865 350270
rect 674754 350212 674865 350214
rect 674799 350209 674865 350212
rect 42351 349976 42417 349979
rect 42306 349974 42417 349976
rect 42306 349918 42356 349974
rect 42412 349918 42417 349974
rect 42306 349913 42417 349918
rect 42306 349650 42366 349913
rect 674031 349532 674097 349535
rect 674754 349532 674814 349576
rect 674031 349530 674814 349532
rect 674031 349474 674036 349530
rect 674092 349474 674814 349530
rect 674031 349472 674814 349474
rect 674031 349469 674097 349472
rect 42351 349088 42417 349091
rect 42306 349086 42417 349088
rect 42306 349030 42356 349086
rect 42412 349030 42417 349086
rect 42306 349025 42417 349030
rect 42306 348910 42366 349025
rect 674127 348792 674193 348795
rect 674127 348790 674784 348792
rect 674127 348734 674132 348790
rect 674188 348734 674784 348790
rect 674127 348732 674784 348734
rect 674127 348729 674193 348732
rect 42306 347904 42366 348022
rect 42306 347844 43518 347904
rect 43215 347756 43281 347759
rect 42306 347754 43281 347756
rect 42306 347698 43220 347754
rect 43276 347698 43281 347754
rect 42306 347696 43281 347698
rect 42306 347208 42366 347696
rect 43215 347693 43281 347696
rect 43215 347608 43281 347611
rect 43458 347608 43518 347844
rect 43215 347606 43518 347608
rect 43215 347550 43220 347606
rect 43276 347550 43518 347606
rect 43215 347548 43518 347550
rect 43215 347545 43281 347548
rect 679746 347463 679806 347948
rect 679746 347458 679857 347463
rect 679746 347402 679796 347458
rect 679852 347402 679857 347458
rect 679746 347400 679857 347402
rect 679791 347397 679857 347400
rect 40378 346806 40384 346870
rect 40448 346806 40454 346870
rect 40386 346542 40446 346806
rect 679791 346720 679857 346723
rect 679746 346718 679857 346720
rect 679746 346662 679796 346718
rect 679852 346662 679857 346718
rect 679746 346657 679857 346662
rect 679746 346468 679806 346657
rect 40570 346214 40576 346278
rect 40640 346214 40646 346278
rect 40578 345728 40638 346214
rect 676474 345474 676480 345538
rect 676544 345536 676550 345538
rect 677103 345536 677169 345539
rect 676544 345534 677169 345536
rect 676544 345478 677108 345534
rect 677164 345478 677169 345534
rect 676544 345476 677169 345478
rect 676544 345474 676550 345476
rect 677103 345473 677169 345476
rect 676282 345326 676288 345390
rect 676352 345388 676358 345390
rect 676911 345388 676977 345391
rect 676352 345386 676977 345388
rect 676352 345330 676916 345386
rect 676972 345330 676977 345386
rect 676352 345328 676977 345330
rect 676352 345326 676358 345328
rect 676911 345325 676977 345328
rect 676666 345178 676672 345242
rect 676736 345240 676742 345242
rect 677007 345240 677073 345243
rect 676736 345238 677073 345240
rect 676736 345182 677012 345238
rect 677068 345182 677073 345238
rect 676736 345180 677073 345182
rect 676736 345178 676742 345180
rect 677007 345177 677073 345180
rect 40962 344354 41022 344914
rect 40954 344290 40960 344354
rect 41024 344290 41030 344354
rect 41922 343615 41982 344100
rect 41871 343610 41982 343615
rect 41871 343554 41876 343610
rect 41932 343554 41982 343610
rect 41871 343552 41982 343554
rect 41871 343549 41937 343552
rect 40770 342874 40830 343286
rect 58383 343168 58449 343171
rect 654447 343168 654513 343171
rect 58383 343166 64416 343168
rect 58383 343110 58388 343166
rect 58444 343110 64416 343166
rect 58383 343108 64416 343110
rect 650208 343166 654513 343168
rect 650208 343110 654452 343166
rect 654508 343110 654513 343166
rect 650208 343108 654513 343110
rect 58383 343105 58449 343108
rect 654447 343105 654513 343108
rect 40762 342810 40768 342874
rect 40832 342810 40838 342874
rect 41154 341986 41214 342472
rect 41146 341922 41152 341986
rect 41216 341922 41222 341986
rect 42114 341246 42174 341806
rect 42106 341182 42112 341246
rect 42176 341182 42182 341246
rect 41730 340359 41790 340918
rect 41730 340354 41841 340359
rect 41730 340298 41780 340354
rect 41836 340298 41841 340354
rect 41730 340296 41841 340298
rect 41775 340293 41841 340296
rect 37314 339915 37374 340178
rect 37314 339910 37425 339915
rect 37314 339854 37364 339910
rect 37420 339854 37425 339910
rect 37314 339852 37425 339854
rect 37359 339849 37425 339852
rect 41346 338730 41406 339290
rect 41338 338666 41344 338730
rect 41408 338666 41414 338730
rect 40002 337991 40062 338550
rect 39951 337986 40062 337991
rect 39951 337930 39956 337986
rect 40012 337930 40062 337986
rect 39951 337928 40062 337930
rect 39951 337925 40017 337928
rect 37122 337399 37182 337662
rect 37122 337394 37233 337399
rect 37122 337338 37172 337394
rect 37228 337338 37233 337394
rect 37122 337336 37233 337338
rect 37167 337333 37233 337336
rect 40047 337248 40113 337251
rect 40002 337246 40113 337248
rect 40002 337190 40052 337246
rect 40108 337190 40113 337246
rect 40002 337185 40113 337190
rect 40002 337070 40062 337185
rect 37359 336508 37425 336511
rect 41530 336508 41536 336510
rect 37359 336506 41536 336508
rect 37359 336450 37364 336506
rect 37420 336450 41536 336506
rect 37359 336448 41536 336450
rect 37359 336445 37425 336448
rect 41530 336446 41536 336448
rect 41600 336446 41606 336510
rect 37314 335623 37374 336182
rect 37314 335618 37425 335623
rect 37314 335562 37364 335618
rect 37420 335562 37425 335618
rect 37314 335560 37425 335562
rect 37359 335557 37425 335560
rect 40194 334883 40254 335442
rect 675471 335178 675537 335179
rect 675471 335174 675520 335178
rect 675584 335176 675590 335178
rect 675471 335118 675476 335174
rect 675471 335114 675520 335118
rect 675584 335116 675628 335176
rect 675584 335114 675590 335116
rect 675471 335113 675537 335114
rect 40194 334878 40305 334883
rect 40194 334822 40244 334878
rect 40300 334822 40305 334878
rect 40194 334820 40305 334822
rect 40239 334817 40305 334820
rect 42306 334436 42366 334554
rect 42543 334436 42609 334439
rect 42306 334434 42609 334436
rect 42306 334378 42548 334434
rect 42604 334378 42609 334434
rect 42306 334376 42609 334378
rect 42543 334373 42609 334376
rect 42306 333551 42366 333814
rect 675322 333782 675328 333846
rect 675392 333844 675398 333846
rect 675471 333844 675537 333847
rect 675392 333842 675537 333844
rect 675392 333786 675476 333842
rect 675532 333786 675537 333842
rect 675392 333784 675537 333786
rect 675392 333782 675398 333784
rect 675471 333781 675537 333784
rect 42255 333546 42366 333551
rect 42255 333490 42260 333546
rect 42316 333490 42366 333546
rect 42255 333488 42366 333490
rect 675759 333548 675825 333551
rect 676282 333548 676288 333550
rect 675759 333546 676288 333548
rect 675759 333490 675764 333546
rect 675820 333490 676288 333546
rect 675759 333488 676288 333490
rect 42255 333485 42321 333488
rect 675759 333485 675825 333488
rect 676282 333486 676288 333488
rect 676352 333486 676358 333550
rect 42306 332071 42366 332260
rect 42255 332066 42366 332071
rect 42255 332010 42260 332066
rect 42316 332010 42366 332066
rect 42255 332008 42366 332010
rect 42255 332005 42321 332008
rect 654447 331624 654513 331627
rect 650208 331622 654513 331624
rect 650208 331566 654452 331622
rect 654508 331566 654513 331622
rect 650208 331564 654513 331566
rect 654447 331561 654513 331564
rect 675183 329552 675249 329555
rect 675514 329552 675520 329554
rect 675183 329550 675520 329552
rect 675183 329494 675188 329550
rect 675244 329494 675520 329550
rect 675183 329492 675520 329494
rect 675183 329489 675249 329492
rect 675514 329490 675520 329492
rect 675584 329490 675590 329554
rect 57807 328812 57873 328815
rect 57807 328810 64416 328812
rect 57807 328754 57812 328810
rect 57868 328754 64416 328810
rect 57807 328752 64416 328754
rect 57807 328749 57873 328752
rect 675759 328072 675825 328075
rect 676474 328072 676480 328074
rect 675759 328070 676480 328072
rect 675759 328014 675764 328070
rect 675820 328014 676480 328070
rect 675759 328012 676480 328014
rect 675759 328009 675825 328012
rect 676474 328010 676480 328012
rect 676544 328010 676550 328074
rect 675759 326888 675825 326891
rect 676666 326888 676672 326890
rect 675759 326886 676672 326888
rect 675759 326830 675764 326886
rect 675820 326830 676672 326886
rect 675759 326828 676672 326830
rect 675759 326825 675825 326828
rect 676666 326826 676672 326828
rect 676736 326826 676742 326890
rect 42063 319786 42129 319787
rect 42063 319782 42112 319786
rect 42176 319784 42182 319786
rect 655119 319784 655185 319787
rect 42063 319726 42068 319782
rect 42063 319722 42112 319726
rect 42176 319724 42220 319784
rect 650208 319782 655185 319784
rect 650208 319726 655124 319782
rect 655180 319726 655185 319782
rect 650208 319724 655185 319726
rect 42176 319722 42182 319724
rect 42063 319721 42129 319722
rect 655119 319721 655185 319724
rect 674415 319710 674481 319713
rect 674415 319708 674784 319710
rect 674415 319652 674420 319708
rect 674476 319652 674784 319708
rect 674415 319650 674784 319652
rect 674415 319647 674481 319650
rect 674415 318896 674481 318899
rect 674415 318894 674784 318896
rect 674415 318838 674420 318894
rect 674476 318838 674784 318894
rect 674415 318836 674784 318838
rect 674415 318833 674481 318836
rect 41871 318750 41937 318751
rect 41871 318748 41920 318750
rect 41828 318746 41920 318748
rect 41828 318690 41876 318746
rect 41828 318688 41920 318690
rect 41871 318686 41920 318688
rect 41984 318686 41990 318750
rect 41871 318685 41937 318686
rect 674703 318304 674769 318307
rect 674703 318302 674814 318304
rect 674703 318246 674708 318302
rect 674764 318246 674814 318302
rect 674703 318241 674814 318246
rect 674754 318052 674814 318241
rect 41775 317862 41841 317863
rect 41722 317798 41728 317862
rect 41792 317860 41841 317862
rect 41792 317858 41884 317860
rect 41836 317802 41884 317858
rect 41792 317800 41884 317802
rect 41792 317798 41841 317800
rect 41775 317797 41841 317798
rect 674362 317206 674368 317270
rect 674432 317268 674438 317270
rect 674432 317208 674784 317268
rect 674432 317206 674438 317208
rect 41338 316022 41344 316086
rect 41408 316084 41414 316086
rect 41775 316084 41841 316087
rect 41408 316082 41841 316084
rect 41408 316026 41780 316082
rect 41836 316026 41841 316082
rect 41408 316024 41841 316026
rect 41408 316022 41414 316024
rect 41775 316021 41841 316024
rect 674946 315938 675006 316424
rect 674938 315874 674944 315938
rect 675008 315874 675014 315938
rect 674170 315726 674176 315790
rect 674240 315788 674246 315790
rect 674240 315728 674784 315788
rect 674240 315726 674246 315728
rect 41146 315430 41152 315494
rect 41216 315492 41222 315494
rect 41775 315492 41841 315495
rect 41216 315490 41841 315492
rect 41216 315434 41780 315490
rect 41836 315434 41841 315490
rect 41216 315432 41841 315434
rect 41216 315430 41222 315432
rect 41775 315429 41841 315432
rect 673978 314838 673984 314902
rect 674048 314900 674054 314902
rect 674048 314870 674784 314900
rect 674048 314840 674814 314870
rect 674048 314838 674054 314840
rect 57999 314604 58065 314607
rect 57999 314602 64416 314604
rect 57999 314546 58004 314602
rect 58060 314546 64416 314602
rect 57999 314544 64416 314546
rect 57999 314541 58065 314544
rect 674554 314246 674560 314310
rect 674624 314308 674630 314310
rect 674754 314308 674814 314840
rect 674624 314248 674814 314308
rect 674624 314246 674630 314248
rect 674031 314160 674097 314163
rect 674031 314158 674784 314160
rect 674031 314102 674036 314158
rect 674092 314102 674784 314158
rect 674031 314100 674784 314102
rect 674031 314097 674097 314100
rect 40954 313654 40960 313718
rect 41024 313716 41030 313718
rect 41871 313716 41937 313719
rect 41024 313714 41937 313716
rect 41024 313658 41876 313714
rect 41932 313658 41937 313714
rect 41024 313656 41937 313658
rect 41024 313654 41030 313656
rect 41871 313653 41937 313656
rect 41530 313210 41536 313274
rect 41600 313272 41606 313274
rect 41775 313272 41841 313275
rect 41600 313270 41841 313272
rect 41600 313214 41780 313270
rect 41836 313214 41841 313270
rect 41600 313212 41841 313214
rect 41600 313210 41606 313212
rect 41775 313209 41841 313212
rect 674362 313210 674368 313274
rect 674432 313272 674438 313274
rect 674432 313212 674784 313272
rect 674432 313210 674438 313212
rect 40762 312322 40768 312386
rect 40832 312384 40838 312386
rect 41775 312384 41841 312387
rect 40832 312382 41841 312384
rect 40832 312326 41780 312382
rect 41836 312326 41841 312382
rect 40832 312324 41841 312326
rect 40832 312322 40838 312324
rect 41775 312321 41841 312324
rect 675138 312239 675198 312502
rect 675087 312234 675198 312239
rect 675087 312178 675092 312234
rect 675148 312178 675198 312234
rect 675087 312176 675198 312178
rect 675087 312173 675153 312176
rect 673935 311644 674001 311647
rect 673935 311642 674784 311644
rect 673935 311586 673940 311642
rect 673996 311586 674784 311642
rect 673935 311584 674784 311586
rect 673935 311581 674001 311584
rect 676866 310759 676926 311022
rect 676866 310754 676977 310759
rect 676866 310698 676916 310754
rect 676972 310698 676977 310754
rect 676866 310696 676977 310698
rect 676911 310693 676977 310696
rect 677058 310019 677118 310134
rect 677058 310014 677169 310019
rect 677058 309958 677108 310014
rect 677164 309958 677169 310014
rect 677058 309956 677169 309958
rect 677103 309953 677169 309956
rect 674946 309131 675006 309394
rect 674895 309126 675006 309131
rect 674895 309070 674900 309126
rect 674956 309070 675006 309126
rect 674895 309068 675006 309070
rect 674895 309065 674961 309068
rect 674223 308536 674289 308539
rect 674223 308534 674784 308536
rect 674223 308478 674228 308534
rect 674284 308478 674784 308534
rect 674223 308476 674784 308478
rect 674223 308473 674289 308476
rect 655215 307944 655281 307947
rect 650208 307942 655281 307944
rect 650208 307886 655220 307942
rect 655276 307886 655281 307942
rect 650208 307884 655281 307886
rect 655215 307881 655281 307884
rect 42351 307500 42417 307503
rect 42306 307498 42417 307500
rect 42306 307442 42356 307498
rect 42412 307442 42417 307498
rect 42306 307437 42417 307442
rect 674607 307500 674673 307503
rect 674754 307500 674814 307766
rect 674607 307498 674814 307500
rect 674607 307442 674612 307498
rect 674668 307442 674814 307498
rect 674607 307440 674814 307442
rect 674607 307437 674673 307440
rect 42306 307322 42366 307437
rect 677058 306763 677118 306878
rect 42351 306760 42417 306763
rect 42306 306758 42417 306760
rect 42306 306702 42356 306758
rect 42412 306702 42417 306758
rect 42306 306697 42417 306702
rect 677007 306758 677118 306763
rect 677007 306702 677012 306758
rect 677068 306702 677118 306758
rect 677007 306700 677118 306702
rect 677007 306697 677073 306700
rect 42306 306434 42366 306697
rect 676866 306023 676926 306212
rect 676815 306018 676926 306023
rect 676815 305962 676820 306018
rect 676876 305962 676926 306018
rect 676815 305960 676926 305962
rect 676815 305957 676881 305960
rect 42306 305431 42366 305694
rect 42306 305426 42417 305431
rect 42306 305370 42356 305426
rect 42412 305370 42417 305426
rect 42306 305368 42417 305370
rect 42351 305365 42417 305368
rect 674319 305428 674385 305431
rect 674319 305426 674784 305428
rect 674319 305370 674324 305426
rect 674380 305370 674784 305426
rect 674319 305368 674784 305370
rect 674319 305365 674385 305368
rect 42306 304244 42366 304806
rect 674415 304614 674481 304617
rect 674415 304612 674784 304614
rect 674415 304556 674420 304612
rect 674476 304556 674784 304612
rect 674415 304554 674784 304556
rect 674415 304551 674481 304554
rect 42306 304184 43518 304244
rect 43215 304096 43281 304099
rect 42336 304094 43281 304096
rect 42336 304038 43220 304094
rect 43276 304038 43281 304094
rect 42336 304036 43281 304038
rect 43215 304033 43281 304036
rect 43215 303948 43281 303951
rect 43458 303948 43518 304184
rect 43215 303946 43518 303948
rect 43215 303890 43220 303946
rect 43276 303890 43518 303946
rect 43215 303888 43518 303890
rect 43215 303885 43281 303888
rect 40378 303738 40384 303802
rect 40448 303738 40454 303802
rect 674127 303800 674193 303803
rect 674127 303798 674784 303800
rect 674127 303742 674132 303798
rect 674188 303742 674784 303798
rect 674127 303740 674784 303742
rect 40386 303356 40446 303738
rect 674127 303737 674193 303740
rect 40386 303326 42336 303356
rect 40416 303296 42366 303326
rect 42306 303210 42366 303296
rect 42298 303146 42304 303210
rect 42368 303146 42374 303210
rect 40570 302998 40576 303062
rect 40640 302998 40646 303062
rect 40578 302542 40638 302998
rect 40578 302512 42144 302542
rect 40608 302482 42174 302512
rect 42114 302322 42174 302482
rect 679746 302471 679806 302956
rect 679746 302466 679857 302471
rect 679746 302410 679796 302466
rect 679852 302410 679857 302466
rect 679746 302408 679857 302410
rect 679791 302405 679857 302408
rect 42106 302258 42112 302322
rect 42176 302258 42182 302322
rect 679791 301728 679857 301731
rect 679746 301726 679857 301728
rect 40770 301138 40830 301698
rect 679746 301670 679796 301726
rect 679852 301670 679857 301726
rect 679746 301665 679857 301670
rect 679746 301402 679806 301665
rect 40762 301074 40768 301138
rect 40832 301074 40838 301138
rect 41922 300399 41982 300884
rect 41871 300394 41982 300399
rect 41871 300338 41876 300394
rect 41932 300338 41982 300394
rect 41871 300336 41982 300338
rect 41871 300333 41937 300336
rect 59439 300100 59505 300103
rect 59439 300098 64416 300100
rect 40962 299658 41022 300070
rect 59439 300042 59444 300098
rect 59500 300042 64416 300098
rect 59439 300040 64416 300042
rect 59439 300037 59505 300040
rect 40954 299594 40960 299658
rect 41024 299594 41030 299658
rect 675898 299446 675904 299510
rect 675968 299508 675974 299510
rect 677007 299508 677073 299511
rect 675968 299506 677073 299508
rect 675968 299450 677012 299506
rect 677068 299450 677073 299506
rect 675968 299448 677073 299450
rect 675968 299446 675974 299448
rect 677007 299445 677073 299448
rect 676666 299298 676672 299362
rect 676736 299360 676742 299362
rect 677103 299360 677169 299363
rect 676736 299358 677169 299360
rect 676736 299302 677108 299358
rect 677164 299302 677169 299358
rect 676736 299300 677169 299302
rect 676736 299298 676742 299300
rect 677103 299297 677169 299300
rect 41154 298770 41214 299256
rect 41146 298706 41152 298770
rect 41216 298706 41222 298770
rect 40386 298030 40446 298590
rect 40378 297966 40384 298030
rect 40448 297966 40454 298030
rect 42306 297291 42366 297776
rect 42255 297286 42366 297291
rect 42255 297230 42260 297286
rect 42316 297230 42366 297286
rect 42255 297228 42366 297230
rect 42255 297225 42321 297228
rect 37314 296699 37374 296962
rect 37314 296694 37425 296699
rect 37314 296638 37364 296694
rect 37420 296638 37425 296694
rect 37314 296636 37425 296638
rect 37359 296633 37425 296636
rect 655407 296252 655473 296255
rect 650208 296250 655473 296252
rect 650208 296194 655412 296250
rect 655468 296194 655473 296250
rect 650208 296192 655473 296194
rect 655407 296189 655473 296192
rect 41538 295514 41598 296074
rect 41530 295450 41536 295514
rect 41600 295450 41606 295514
rect 40002 294775 40062 295334
rect 40002 294770 40113 294775
rect 40002 294714 40052 294770
rect 40108 294714 40113 294770
rect 40002 294712 40113 294714
rect 40047 294709 40113 294712
rect 37314 294035 37374 294446
rect 37263 294030 37374 294035
rect 37263 293974 37268 294030
rect 37324 293974 37374 294030
rect 37263 293972 37374 293974
rect 40143 294032 40209 294035
rect 40143 294030 40254 294032
rect 40143 293974 40148 294030
rect 40204 293974 40254 294030
rect 37263 293969 37329 293972
rect 40143 293969 40254 293974
rect 40194 293854 40254 293969
rect 37359 292404 37425 292407
rect 41338 292404 41344 292406
rect 37359 292402 41344 292404
rect 37359 292346 37364 292402
rect 37420 292346 41344 292402
rect 37359 292344 41344 292346
rect 37359 292341 37425 292344
rect 41338 292342 41344 292344
rect 41408 292342 41414 292406
rect 42306 292404 42366 292966
rect 42447 292404 42513 292407
rect 42306 292402 42513 292404
rect 42306 292346 42452 292402
rect 42508 292346 42513 292402
rect 42306 292344 42513 292346
rect 42447 292341 42513 292344
rect 40194 291667 40254 292226
rect 40194 291662 40305 291667
rect 40194 291606 40244 291662
rect 40300 291606 40305 291662
rect 40194 291604 40305 291606
rect 40239 291601 40305 291604
rect 42927 291368 42993 291371
rect 42336 291366 42993 291368
rect 42336 291310 42932 291366
rect 42988 291310 42993 291366
rect 42336 291308 42993 291310
rect 42927 291305 42993 291308
rect 42306 290036 42366 290598
rect 42306 289976 42750 290036
rect 42690 289592 42750 289976
rect 675471 289742 675537 289743
rect 675471 289740 675520 289742
rect 675428 289738 675520 289740
rect 675428 289682 675476 289738
rect 675428 289680 675520 289682
rect 675471 289678 675520 289680
rect 675584 289678 675590 289742
rect 675471 289677 675537 289678
rect 675375 289594 675441 289595
rect 675322 289592 675328 289594
rect 42306 289532 42750 289592
rect 675284 289532 675328 289592
rect 675392 289590 675441 289594
rect 675436 289534 675441 289590
rect 42306 288855 42366 289532
rect 675322 289530 675328 289532
rect 675392 289530 675441 289534
rect 675375 289529 675441 289530
rect 42255 288850 42366 288855
rect 42255 288794 42260 288850
rect 42316 288794 42366 288850
rect 42255 288792 42366 288794
rect 42255 288789 42321 288792
rect 58095 285892 58161 285895
rect 58095 285890 64416 285892
rect 58095 285834 58100 285890
rect 58156 285834 64416 285890
rect 58095 285832 64416 285834
rect 58095 285829 58161 285832
rect 674746 284942 674752 285006
rect 674816 285004 674822 285006
rect 675183 285004 675249 285007
rect 674816 285002 675249 285004
rect 674816 284946 675188 285002
rect 675244 284946 675249 285002
rect 674816 284944 675249 284946
rect 674816 284942 674822 284944
rect 675183 284941 675249 284944
rect 675759 284856 675825 284859
rect 675898 284856 675904 284858
rect 675759 284854 675904 284856
rect 675759 284798 675764 284854
rect 675820 284798 675904 284854
rect 675759 284796 675904 284798
rect 675759 284793 675825 284796
rect 675898 284794 675904 284796
rect 675968 284794 675974 284858
rect 654447 284708 654513 284711
rect 650208 284706 654513 284708
rect 650208 284650 654452 284706
rect 654508 284650 654513 284706
rect 650208 284648 654513 284650
rect 654447 284645 654513 284648
rect 40527 284118 40593 284119
rect 40527 284116 40576 284118
rect 40484 284114 40576 284116
rect 40484 284058 40532 284114
rect 40484 284056 40576 284058
rect 40527 284054 40576 284056
rect 40640 284054 40646 284118
rect 40527 284053 40593 284054
rect 674362 283610 674368 283674
rect 674432 283672 674438 283674
rect 675375 283672 675441 283675
rect 674432 283670 675441 283672
rect 674432 283614 675380 283670
rect 675436 283614 675441 283670
rect 674432 283612 675441 283614
rect 674432 283610 674438 283612
rect 675375 283609 675441 283612
rect 42255 283378 42321 283379
rect 42255 283376 42304 283378
rect 42212 283374 42304 283376
rect 42212 283318 42260 283374
rect 42212 283316 42304 283318
rect 42255 283314 42304 283316
rect 42368 283314 42374 283378
rect 42255 283313 42321 283314
rect 42447 282488 42513 282491
rect 42682 282488 42688 282490
rect 42447 282486 42688 282488
rect 42447 282430 42452 282486
rect 42508 282430 42688 282486
rect 42447 282428 42688 282430
rect 42447 282425 42513 282428
rect 42682 282426 42688 282428
rect 42752 282426 42758 282490
rect 675759 281896 675825 281899
rect 676666 281896 676672 281898
rect 675759 281894 676672 281896
rect 675759 281838 675764 281894
rect 675820 281838 676672 281894
rect 675759 281836 676672 281838
rect 675759 281833 675825 281836
rect 676666 281834 676672 281836
rect 676736 281834 676742 281898
rect 40570 279762 40576 279826
rect 40640 279824 40646 279826
rect 41775 279824 41841 279827
rect 40640 279822 41841 279824
rect 40640 279766 41780 279822
rect 41836 279766 41841 279822
rect 40640 279764 41841 279766
rect 40640 279762 40646 279764
rect 41775 279761 41841 279764
rect 372879 278640 372945 278643
rect 84354 278638 372945 278640
rect 84354 278582 372884 278638
rect 372940 278582 372945 278638
rect 84354 278580 372945 278582
rect 82863 278492 82929 278495
rect 84354 278492 84414 278580
rect 372879 278577 372945 278580
rect 374319 278640 374385 278643
rect 395055 278640 395121 278643
rect 374319 278638 395121 278640
rect 374319 278582 374324 278638
rect 374380 278582 395060 278638
rect 395116 278582 395121 278638
rect 374319 278580 395121 278582
rect 374319 278577 374385 278580
rect 395055 278577 395121 278580
rect 82863 278490 84414 278492
rect 82863 278434 82868 278490
rect 82924 278434 84414 278490
rect 82863 278432 84414 278434
rect 304527 278492 304593 278495
rect 474735 278492 474801 278495
rect 304527 278490 474801 278492
rect 304527 278434 304532 278490
rect 304588 278434 474740 278490
rect 474796 278434 474801 278490
rect 304527 278432 474801 278434
rect 82863 278429 82929 278432
rect 304527 278429 304593 278432
rect 474735 278429 474801 278432
rect 305199 278344 305265 278347
rect 481839 278344 481905 278347
rect 305199 278342 481905 278344
rect 305199 278286 305204 278342
rect 305260 278286 481844 278342
rect 481900 278286 481905 278342
rect 305199 278284 481905 278286
rect 305199 278281 305265 278284
rect 481839 278281 481905 278284
rect 305583 278196 305649 278199
rect 485391 278196 485457 278199
rect 305583 278194 485457 278196
rect 305583 278138 305588 278194
rect 305644 278138 485396 278194
rect 485452 278138 485457 278194
rect 305583 278136 485457 278138
rect 305583 278133 305649 278136
rect 485391 278133 485457 278136
rect 306351 278048 306417 278051
rect 488943 278048 489009 278051
rect 306351 278046 489009 278048
rect 306351 277990 306356 278046
rect 306412 277990 488948 278046
rect 489004 277990 489009 278046
rect 306351 277988 489009 277990
rect 306351 277985 306417 277988
rect 488943 277985 489009 277988
rect 307023 277900 307089 277903
rect 496143 277900 496209 277903
rect 307023 277898 496209 277900
rect 307023 277842 307028 277898
rect 307084 277842 496148 277898
rect 496204 277842 496209 277898
rect 307023 277840 496209 277842
rect 307023 277837 307089 277840
rect 496143 277837 496209 277840
rect 307791 277752 307857 277755
rect 503247 277752 503313 277755
rect 307791 277750 503313 277752
rect 307791 277694 307796 277750
rect 307852 277694 503252 277750
rect 503308 277694 503313 277750
rect 307791 277692 503313 277694
rect 307791 277689 307857 277692
rect 503247 277689 503313 277692
rect 309519 277604 309585 277607
rect 517743 277604 517809 277607
rect 309519 277602 517809 277604
rect 309519 277546 309524 277602
rect 309580 277546 517748 277602
rect 517804 277546 517809 277602
rect 309519 277544 517809 277546
rect 309519 277541 309585 277544
rect 517743 277541 517809 277544
rect 310383 277456 310449 277459
rect 524943 277456 525009 277459
rect 310383 277454 525009 277456
rect 310383 277398 310388 277454
rect 310444 277398 524948 277454
rect 525004 277398 525009 277454
rect 310383 277396 525009 277398
rect 310383 277393 310449 277396
rect 524943 277393 525009 277396
rect 311535 277308 311601 277311
rect 532143 277308 532209 277311
rect 311535 277306 532209 277308
rect 311535 277250 311540 277306
rect 311596 277250 532148 277306
rect 532204 277250 532209 277306
rect 311535 277248 532209 277250
rect 311535 277245 311601 277248
rect 532143 277245 532209 277248
rect 311631 277160 311697 277163
rect 535599 277160 535665 277163
rect 311631 277158 535665 277160
rect 311631 277102 311636 277158
rect 311692 277102 535604 277158
rect 535660 277102 535665 277158
rect 311631 277100 535665 277102
rect 311631 277097 311697 277100
rect 535599 277097 535665 277100
rect 313167 277012 313233 277015
rect 546351 277012 546417 277015
rect 313167 277010 546417 277012
rect 313167 276954 313172 277010
rect 313228 276954 546356 277010
rect 546412 276954 546417 277010
rect 313167 276952 546417 276954
rect 313167 276949 313233 276952
rect 546351 276949 546417 276952
rect 120495 276864 120561 276867
rect 375183 276864 375249 276867
rect 120495 276862 375249 276864
rect 120495 276806 120500 276862
rect 120556 276806 375188 276862
rect 375244 276806 375249 276862
rect 120495 276804 375249 276806
rect 120495 276801 120561 276804
rect 375183 276801 375249 276804
rect 375375 276864 375441 276867
rect 393711 276864 393777 276867
rect 375375 276862 393777 276864
rect 375375 276806 375380 276862
rect 375436 276806 393716 276862
rect 393772 276806 393777 276862
rect 375375 276804 393777 276806
rect 375375 276801 375441 276804
rect 393711 276801 393777 276804
rect 113487 276716 113553 276719
rect 375279 276716 375345 276719
rect 113487 276714 375345 276716
rect 113487 276658 113492 276714
rect 113548 276658 375284 276714
rect 375340 276658 375345 276714
rect 113487 276656 375345 276658
rect 113487 276653 113553 276656
rect 375279 276653 375345 276656
rect 375471 276716 375537 276719
rect 388719 276716 388785 276719
rect 375471 276714 388785 276716
rect 375471 276658 375476 276714
rect 375532 276658 388724 276714
rect 388780 276658 388785 276714
rect 375471 276656 388785 276658
rect 375471 276653 375537 276656
rect 388719 276653 388785 276656
rect 40378 276506 40384 276570
rect 40448 276568 40454 276570
rect 41775 276568 41841 276571
rect 40448 276566 41841 276568
rect 40448 276510 41780 276566
rect 41836 276510 41841 276566
rect 40448 276508 41841 276510
rect 40448 276506 40454 276508
rect 41775 276505 41841 276508
rect 303375 276568 303441 276571
rect 467823 276568 467889 276571
rect 303375 276566 467889 276568
rect 303375 276510 303380 276566
rect 303436 276510 467828 276566
rect 467884 276510 467889 276566
rect 303375 276508 467889 276510
rect 303375 276505 303441 276508
rect 467823 276505 467889 276508
rect 262671 276420 262737 276423
rect 320175 276420 320241 276423
rect 603375 276420 603441 276423
rect 262671 276418 268926 276420
rect 262671 276362 262676 276418
rect 262732 276362 268926 276418
rect 262671 276360 268926 276362
rect 262671 276357 262737 276360
rect 262863 276124 262929 276127
rect 268866 276124 268926 276360
rect 320175 276418 603441 276420
rect 320175 276362 320180 276418
rect 320236 276362 603380 276418
rect 603436 276362 603441 276418
rect 320175 276360 603441 276362
rect 320175 276357 320241 276360
rect 603375 276357 603441 276360
rect 299631 276272 299697 276275
rect 322479 276272 322545 276275
rect 299631 276270 322545 276272
rect 299631 276214 299636 276270
rect 299692 276214 322484 276270
rect 322540 276214 322545 276270
rect 299631 276212 322545 276214
rect 299631 276209 299697 276212
rect 322479 276209 322545 276212
rect 322671 276272 322737 276275
rect 624879 276272 624945 276275
rect 322671 276270 624945 276272
rect 322671 276214 322676 276270
rect 322732 276214 624884 276270
rect 624940 276214 624945 276270
rect 322671 276212 624945 276214
rect 322671 276209 322737 276212
rect 624879 276209 624945 276212
rect 429135 276124 429201 276127
rect 262863 276122 268734 276124
rect 262863 276066 262868 276122
rect 262924 276066 268734 276122
rect 262863 276064 268734 276066
rect 268866 276122 429201 276124
rect 268866 276066 429140 276122
rect 429196 276066 429201 276122
rect 268866 276064 429201 276066
rect 262863 276061 262929 276064
rect 263631 275976 263697 275979
rect 268674 275976 268734 276064
rect 429135 276061 429201 276064
rect 449199 276124 449265 276127
rect 469455 276124 469521 276127
rect 449199 276122 469521 276124
rect 449199 276066 449204 276122
rect 449260 276066 469460 276122
rect 469516 276066 469521 276122
rect 449199 276064 469521 276066
rect 449199 276061 449265 276064
rect 469455 276061 469521 276064
rect 489519 276124 489585 276127
rect 509775 276124 509841 276127
rect 489519 276122 509841 276124
rect 489519 276066 489524 276122
rect 489580 276066 509780 276122
rect 509836 276066 509841 276122
rect 489519 276064 509841 276066
rect 489519 276061 489585 276064
rect 509775 276061 509841 276064
rect 529839 276124 529905 276127
rect 545679 276124 545745 276127
rect 529839 276122 545745 276124
rect 529839 276066 529844 276122
rect 529900 276066 545684 276122
rect 545740 276066 545745 276122
rect 529839 276064 545745 276066
rect 529839 276061 529905 276064
rect 545679 276061 545745 276064
rect 570063 276124 570129 276127
rect 587919 276124 587985 276127
rect 570063 276122 587985 276124
rect 570063 276066 570068 276122
rect 570124 276066 587924 276122
rect 587980 276066 587985 276122
rect 570063 276064 587985 276066
rect 570063 276061 570129 276064
rect 587919 276061 587985 276064
rect 591567 275976 591633 275979
rect 263631 275974 268542 275976
rect 263631 275918 263636 275974
rect 263692 275918 268542 275974
rect 263631 275916 268542 275918
rect 268674 275974 591633 275976
rect 268674 275918 591572 275974
rect 591628 275918 591633 275974
rect 268674 275916 591633 275918
rect 263631 275913 263697 275916
rect 263727 275828 263793 275831
rect 268482 275828 268542 275916
rect 591567 275913 591633 275916
rect 595119 275828 595185 275831
rect 263727 275826 268350 275828
rect 263727 275770 263732 275826
rect 263788 275770 268350 275826
rect 263727 275768 268350 275770
rect 268482 275826 595185 275828
rect 268482 275770 595124 275826
rect 595180 275770 595185 275826
rect 268482 275768 595185 275770
rect 263727 275765 263793 275768
rect 264399 275680 264465 275683
rect 268143 275680 268209 275683
rect 264399 275678 268209 275680
rect 264399 275622 264404 275678
rect 264460 275622 268148 275678
rect 268204 275622 268209 275678
rect 264399 275620 268209 275622
rect 268290 275680 268350 275768
rect 595119 275765 595185 275768
rect 598767 275680 598833 275683
rect 268290 275678 598833 275680
rect 268290 275622 598772 275678
rect 598828 275622 598833 275678
rect 268290 275620 598833 275622
rect 264399 275617 264465 275620
rect 268143 275617 268209 275620
rect 598767 275617 598833 275620
rect 41967 275534 42033 275535
rect 41914 275470 41920 275534
rect 41984 275532 42033 275534
rect 42874 275532 42880 275534
rect 41984 275530 42880 275532
rect 42028 275474 42880 275530
rect 41984 275472 42880 275474
rect 41984 275470 42033 275472
rect 42874 275470 42880 275472
rect 42944 275470 42950 275534
rect 265455 275532 265521 275535
rect 268815 275532 268881 275535
rect 602223 275532 602289 275535
rect 265455 275530 268734 275532
rect 265455 275474 265460 275530
rect 265516 275474 268734 275530
rect 265455 275472 268734 275474
rect 41967 275469 42033 275470
rect 265455 275469 265521 275472
rect 267663 275384 267729 275387
rect 267855 275384 267921 275387
rect 267663 275382 267921 275384
rect 267663 275326 267668 275382
rect 267724 275326 267860 275382
rect 267916 275326 267921 275382
rect 267663 275324 267921 275326
rect 268674 275384 268734 275472
rect 268815 275530 602289 275532
rect 268815 275474 268820 275530
rect 268876 275474 602228 275530
rect 602284 275474 602289 275530
rect 268815 275472 602289 275474
rect 268815 275469 268881 275472
rect 602223 275469 602289 275472
rect 612975 275384 613041 275387
rect 268674 275382 613041 275384
rect 268674 275326 612980 275382
rect 613036 275326 613041 275382
rect 268674 275324 613041 275326
rect 267663 275321 267729 275324
rect 267855 275321 267921 275324
rect 612975 275321 613041 275324
rect 265935 275236 266001 275239
rect 616527 275236 616593 275239
rect 265935 275234 616593 275236
rect 265935 275178 265940 275234
rect 265996 275178 616532 275234
rect 616588 275178 616593 275234
rect 265935 275176 616593 275178
rect 265935 275173 266001 275176
rect 616527 275173 616593 275176
rect 620559 275236 620625 275239
rect 637935 275236 638001 275239
rect 620559 275234 638001 275236
rect 620559 275178 620564 275234
rect 620620 275178 637940 275234
rect 637996 275178 638001 275234
rect 620559 275176 638001 275178
rect 620559 275173 620625 275176
rect 637935 275173 638001 275176
rect 266895 275088 266961 275091
rect 623631 275088 623697 275091
rect 266895 275086 623697 275088
rect 266895 275030 266900 275086
rect 266956 275030 623636 275086
rect 623692 275030 623697 275086
rect 266895 275028 623697 275030
rect 266895 275025 266961 275028
rect 623631 275025 623697 275028
rect 41775 274942 41841 274943
rect 41722 274878 41728 274942
rect 41792 274940 41841 274942
rect 261999 274940 262065 274943
rect 369999 274940 370065 274943
rect 378490 274940 378496 274942
rect 41792 274938 41884 274940
rect 41836 274882 41884 274938
rect 41792 274880 41884 274882
rect 261999 274938 370065 274940
rect 261999 274882 262004 274938
rect 262060 274882 370004 274938
rect 370060 274882 370065 274938
rect 261999 274880 370065 274882
rect 41792 274878 41841 274880
rect 41775 274877 41841 274878
rect 261999 274877 262065 274880
rect 369999 274877 370065 274880
rect 370242 274880 378496 274940
rect 259407 274792 259473 274795
rect 368463 274792 368529 274795
rect 259407 274790 368529 274792
rect 259407 274734 259412 274790
rect 259468 274734 368468 274790
rect 368524 274734 368529 274790
rect 259407 274732 368529 274734
rect 259407 274729 259473 274732
rect 368463 274729 368529 274732
rect 253935 274644 254001 274647
rect 370242 274644 370302 274880
rect 378490 274878 378496 274880
rect 378560 274878 378566 274942
rect 378831 274940 378897 274943
rect 645135 274940 645201 274943
rect 378831 274938 645201 274940
rect 378831 274882 378836 274938
rect 378892 274882 645140 274938
rect 645196 274882 645201 274938
rect 378831 274880 645201 274882
rect 378831 274877 378897 274880
rect 645135 274877 645201 274880
rect 674703 274940 674769 274943
rect 674703 274938 674814 274940
rect 674703 274882 674708 274938
rect 674764 274882 674814 274938
rect 674703 274877 674814 274882
rect 370383 274792 370449 274795
rect 620559 274792 620625 274795
rect 370383 274790 620625 274792
rect 370383 274734 370388 274790
rect 370444 274734 620564 274790
rect 620620 274734 620625 274790
rect 370383 274732 620625 274734
rect 370383 274729 370449 274732
rect 620559 274729 620625 274732
rect 674754 274688 674814 274877
rect 253935 274642 370302 274644
rect 253935 274586 253940 274642
rect 253996 274586 370302 274642
rect 253935 274584 370302 274586
rect 372399 274644 372465 274647
rect 409167 274644 409233 274647
rect 372399 274642 409233 274644
rect 372399 274586 372404 274642
rect 372460 274586 409172 274642
rect 409228 274586 409233 274642
rect 372399 274584 409233 274586
rect 253935 274581 254001 274584
rect 372399 274581 372465 274584
rect 409167 274581 409233 274584
rect 429039 274644 429105 274647
rect 429231 274644 429297 274647
rect 429039 274642 429297 274644
rect 429039 274586 429044 274642
rect 429100 274586 429236 274642
rect 429292 274586 429297 274642
rect 429039 274584 429297 274586
rect 429039 274581 429105 274584
rect 429231 274581 429297 274584
rect 449103 274644 449169 274647
rect 469551 274644 469617 274647
rect 449103 274642 469617 274644
rect 449103 274586 449108 274642
rect 449164 274586 469556 274642
rect 469612 274586 469617 274642
rect 449103 274584 469617 274586
rect 449103 274581 449169 274584
rect 469551 274581 469617 274584
rect 489423 274644 489489 274647
rect 504399 274644 504465 274647
rect 489423 274642 504465 274644
rect 489423 274586 489428 274642
rect 489484 274586 504404 274642
rect 504460 274586 504465 274642
rect 489423 274584 504465 274586
rect 489423 274581 489489 274584
rect 504399 274581 504465 274584
rect 252399 274496 252465 274499
rect 505935 274496 506001 274499
rect 252399 274494 506001 274496
rect 252399 274438 252404 274494
rect 252460 274438 505940 274494
rect 505996 274438 506001 274494
rect 252399 274436 506001 274438
rect 252399 274433 252465 274436
rect 505935 274433 506001 274436
rect 509775 274496 509841 274499
rect 529839 274496 529905 274499
rect 509775 274494 529905 274496
rect 509775 274438 509780 274494
rect 509836 274438 529844 274494
rect 529900 274438 529905 274494
rect 509775 274436 529905 274438
rect 509775 274433 509841 274436
rect 529839 274433 529905 274436
rect 545679 274496 545745 274499
rect 570063 274496 570129 274499
rect 545679 274494 570129 274496
rect 545679 274438 545684 274494
rect 545740 274438 570068 274494
rect 570124 274438 570129 274494
rect 545679 274436 570129 274438
rect 545679 274433 545745 274436
rect 570063 274433 570129 274436
rect 584751 274496 584817 274499
rect 593295 274496 593361 274499
rect 584751 274494 593361 274496
rect 584751 274438 584756 274494
rect 584812 274438 593300 274494
rect 593356 274438 593361 274494
rect 584751 274436 593361 274438
rect 584751 274433 584817 274436
rect 593295 274433 593361 274436
rect 613359 274496 613425 274499
rect 613359 274494 616446 274496
rect 613359 274438 613364 274494
rect 613420 274438 616446 274494
rect 613359 274436 616446 274438
rect 613359 274433 613425 274436
rect 251823 274348 251889 274351
rect 573039 274348 573105 274351
rect 584559 274348 584625 274351
rect 251823 274346 492414 274348
rect 251823 274290 251828 274346
rect 251884 274290 492414 274346
rect 251823 274288 492414 274290
rect 251823 274285 251889 274288
rect 42159 274200 42225 274203
rect 42682 274200 42688 274202
rect 42159 274198 42688 274200
rect 42159 274142 42164 274198
rect 42220 274142 42688 274198
rect 42159 274140 42688 274142
rect 42159 274137 42225 274140
rect 42682 274138 42688 274140
rect 42752 274138 42758 274202
rect 250671 274200 250737 274203
rect 491631 274200 491697 274203
rect 250671 274198 491697 274200
rect 250671 274142 250676 274198
rect 250732 274142 491636 274198
rect 491692 274142 491697 274198
rect 250671 274140 491697 274142
rect 492354 274200 492414 274288
rect 573039 274346 584625 274348
rect 573039 274290 573044 274346
rect 573100 274290 584564 274346
rect 584620 274290 584625 274346
rect 573039 274288 584625 274290
rect 616386 274348 616446 274436
rect 619119 274348 619185 274351
rect 616386 274346 619185 274348
rect 616386 274290 619124 274346
rect 619180 274290 619185 274346
rect 616386 274288 619185 274290
rect 573039 274285 573105 274288
rect 584559 274285 584625 274288
rect 619119 274285 619185 274288
rect 498831 274200 498897 274203
rect 492354 274198 498897 274200
rect 492354 274142 498836 274198
rect 498892 274142 498897 274198
rect 492354 274140 498897 274142
rect 250671 274137 250737 274140
rect 491631 274137 491697 274140
rect 498831 274137 498897 274140
rect 504399 274200 504465 274203
rect 552975 274200 553041 274203
rect 504399 274198 545790 274200
rect 504399 274142 504404 274198
rect 504460 274142 545790 274198
rect 504399 274140 545790 274142
rect 504399 274137 504465 274140
rect 249807 274052 249873 274055
rect 484431 274052 484497 274055
rect 249807 274050 484497 274052
rect 249807 273994 249812 274050
rect 249868 273994 484436 274050
rect 484492 273994 484497 274050
rect 249807 273992 484497 273994
rect 545730 274052 545790 274140
rect 550098 274198 553041 274200
rect 550098 274142 552980 274198
rect 553036 274142 553041 274198
rect 550098 274140 553041 274142
rect 550098 274052 550158 274140
rect 552975 274137 553041 274140
rect 545730 273992 550158 274052
rect 674703 274052 674769 274055
rect 674703 274050 674814 274052
rect 674703 273994 674708 274050
rect 674764 273994 674814 274050
rect 249807 273989 249873 273992
rect 484431 273989 484497 273992
rect 674703 273989 674814 273994
rect 249135 273904 249201 273907
rect 477423 273904 477489 273907
rect 249135 273902 477489 273904
rect 249135 273846 249140 273902
rect 249196 273846 477428 273902
rect 477484 273846 477489 273902
rect 249135 273844 477489 273846
rect 249135 273841 249201 273844
rect 477423 273841 477489 273844
rect 477615 273904 477681 273907
rect 489423 273904 489489 273907
rect 477615 273902 489489 273904
rect 477615 273846 477620 273902
rect 477676 273846 489428 273902
rect 489484 273846 489489 273902
rect 674754 273874 674814 273989
rect 477615 273844 489489 273846
rect 477615 273841 477681 273844
rect 489423 273841 489489 273844
rect 42255 273758 42321 273759
rect 42255 273756 42304 273758
rect 42212 273754 42304 273756
rect 42212 273698 42260 273754
rect 42212 273696 42304 273698
rect 42255 273694 42304 273696
rect 42368 273694 42374 273758
rect 255087 273756 255153 273759
rect 381231 273756 381297 273759
rect 383343 273756 383409 273759
rect 255087 273754 378414 273756
rect 255087 273698 255092 273754
rect 255148 273698 378414 273754
rect 255087 273696 378414 273698
rect 42255 273693 42321 273694
rect 255087 273693 255153 273696
rect 116559 273608 116625 273611
rect 146895 273608 146961 273611
rect 116559 273606 146961 273608
rect 116559 273550 116564 273606
rect 116620 273550 146900 273606
rect 146956 273550 146961 273606
rect 116559 273548 146961 273550
rect 116559 273545 116625 273548
rect 146895 273545 146961 273548
rect 187215 273608 187281 273611
rect 207279 273608 207345 273611
rect 187215 273606 207345 273608
rect 187215 273550 187220 273606
rect 187276 273550 207284 273606
rect 207340 273550 207345 273606
rect 187215 273548 207345 273550
rect 187215 273545 187281 273548
rect 207279 273545 207345 273548
rect 248175 273608 248241 273611
rect 368506 273608 368512 273610
rect 248175 273606 368512 273608
rect 248175 273550 248180 273606
rect 248236 273550 368512 273606
rect 248175 273548 368512 273550
rect 248175 273545 248241 273548
rect 368506 273546 368512 273548
rect 368576 273546 368582 273610
rect 377967 273608 378033 273611
rect 378159 273610 378225 273611
rect 368946 273606 378033 273608
rect 368946 273550 377972 273606
rect 378028 273550 378033 273606
rect 368946 273548 378033 273550
rect 88431 273460 88497 273463
rect 156879 273460 156945 273463
rect 88431 273458 156945 273460
rect 88431 273402 88436 273458
rect 88492 273402 156884 273458
rect 156940 273402 156945 273458
rect 88431 273400 156945 273402
rect 88431 273397 88497 273400
rect 156879 273397 156945 273400
rect 177039 273460 177105 273463
rect 194511 273460 194577 273463
rect 177039 273458 194577 273460
rect 177039 273402 177044 273458
rect 177100 273402 194516 273458
rect 194572 273402 194577 273458
rect 177039 273400 194577 273402
rect 177039 273397 177105 273400
rect 194511 273397 194577 273400
rect 212559 273460 212625 273463
rect 237615 273460 237681 273463
rect 212559 273458 237681 273460
rect 212559 273402 212564 273458
rect 212620 273402 237620 273458
rect 237676 273402 237681 273458
rect 212559 273400 237681 273402
rect 212559 273397 212625 273400
rect 237615 273397 237681 273400
rect 257679 273460 257745 273463
rect 368946 273460 369006 273548
rect 377967 273545 378033 273548
rect 378106 273546 378112 273610
rect 378176 273608 378225 273610
rect 378354 273608 378414 273696
rect 379458 273754 381297 273756
rect 379458 273698 381236 273754
rect 381292 273698 381297 273754
rect 379458 273696 381297 273698
rect 379458 273608 379518 273696
rect 381231 273693 381297 273696
rect 383106 273754 383409 273756
rect 383106 273698 383348 273754
rect 383404 273698 383409 273754
rect 383106 273696 383409 273698
rect 378176 273606 378268 273608
rect 378220 273550 378268 273606
rect 378176 273548 378268 273550
rect 378354 273548 379518 273608
rect 379695 273608 379761 273611
rect 383106 273608 383166 273696
rect 383343 273693 383409 273696
rect 383535 273756 383601 273759
rect 389679 273756 389745 273759
rect 383535 273754 389745 273756
rect 383535 273698 383540 273754
rect 383596 273698 389684 273754
rect 389740 273698 389745 273754
rect 383535 273696 389745 273698
rect 383535 273693 383601 273696
rect 389679 273693 389745 273696
rect 409167 273756 409233 273759
rect 428943 273756 429009 273759
rect 409167 273754 429009 273756
rect 409167 273698 409172 273754
rect 409228 273698 428948 273754
rect 429004 273698 429009 273754
rect 409167 273696 429009 273698
rect 409167 273693 409233 273696
rect 428943 273693 429009 273696
rect 429135 273756 429201 273759
rect 449199 273756 449265 273759
rect 429135 273754 449265 273756
rect 429135 273698 429140 273754
rect 429196 273698 449204 273754
rect 449260 273698 449265 273754
rect 429135 273696 449265 273698
rect 429135 273693 429201 273696
rect 449199 273693 449265 273696
rect 469455 273756 469521 273759
rect 489519 273756 489585 273759
rect 469455 273754 489585 273756
rect 469455 273698 469460 273754
rect 469516 273698 489524 273754
rect 489580 273698 489585 273754
rect 469455 273696 489585 273698
rect 469455 273693 469521 273696
rect 489519 273693 489585 273696
rect 379695 273606 383166 273608
rect 379695 273550 379700 273606
rect 379756 273550 383166 273606
rect 379695 273548 383166 273550
rect 383247 273608 383313 273611
rect 648687 273608 648753 273611
rect 383247 273606 648753 273608
rect 383247 273550 383252 273606
rect 383308 273550 648692 273606
rect 648748 273550 648753 273606
rect 383247 273548 648753 273550
rect 378176 273546 378225 273548
rect 378159 273545 378225 273546
rect 379695 273545 379761 273548
rect 383247 273545 383313 273548
rect 648687 273545 648753 273548
rect 257679 273458 369006 273460
rect 257679 273402 257684 273458
rect 257740 273402 369006 273458
rect 257679 273400 369006 273402
rect 369135 273460 369201 273463
rect 379215 273460 379281 273463
rect 369135 273458 379281 273460
rect 369135 273402 369140 273458
rect 369196 273402 379220 273458
rect 379276 273402 379281 273458
rect 369135 273400 379281 273402
rect 257679 273397 257745 273400
rect 369135 273397 369201 273400
rect 379215 273397 379281 273400
rect 379407 273460 379473 273463
rect 381807 273460 381873 273463
rect 379407 273458 381873 273460
rect 379407 273402 379412 273458
rect 379468 273402 381812 273458
rect 381868 273402 381873 273458
rect 379407 273400 381873 273402
rect 379407 273397 379473 273400
rect 381807 273397 381873 273400
rect 383151 273460 383217 273463
rect 605775 273460 605841 273463
rect 383151 273458 605841 273460
rect 383151 273402 383156 273458
rect 383212 273402 605780 273458
rect 605836 273402 605841 273458
rect 383151 273400 605841 273402
rect 383151 273397 383217 273400
rect 605775 273397 605841 273400
rect 83631 273312 83697 273315
rect 156975 273312 157041 273315
rect 83631 273310 157041 273312
rect 83631 273254 83636 273310
rect 83692 273254 156980 273310
rect 157036 273254 157041 273310
rect 83631 273252 157041 273254
rect 83631 273249 83697 273252
rect 156975 273249 157041 273252
rect 157167 273312 157233 273315
rect 177423 273312 177489 273315
rect 157167 273310 177489 273312
rect 157167 273254 157172 273310
rect 157228 273254 177428 273310
rect 177484 273254 177489 273310
rect 157167 273252 177489 273254
rect 157167 273249 157233 273252
rect 177423 273249 177489 273252
rect 177711 273312 177777 273315
rect 197583 273312 197649 273315
rect 177711 273310 197649 273312
rect 177711 273254 177716 273310
rect 177772 273254 197588 273310
rect 197644 273254 197649 273310
rect 177711 273252 197649 273254
rect 177711 273249 177777 273252
rect 197583 273249 197649 273252
rect 217359 273312 217425 273315
rect 237711 273312 237777 273315
rect 217359 273310 237777 273312
rect 217359 273254 217364 273310
rect 217420 273254 237716 273310
rect 237772 273254 237777 273310
rect 217359 273252 237777 273254
rect 217359 273249 217425 273252
rect 237711 273249 237777 273252
rect 250575 273312 250641 273315
rect 378106 273312 378112 273314
rect 250575 273310 378112 273312
rect 250575 273254 250580 273310
rect 250636 273254 378112 273310
rect 250575 273252 378112 273254
rect 250575 273249 250641 273252
rect 378106 273250 378112 273252
rect 378176 273250 378182 273314
rect 379023 273312 379089 273315
rect 584367 273312 584433 273315
rect 379023 273310 584433 273312
rect 379023 273254 379028 273310
rect 379084 273254 584372 273310
rect 584428 273254 584433 273310
rect 379023 273252 584433 273254
rect 379023 273249 379089 273252
rect 584367 273249 584433 273252
rect 674703 273312 674769 273315
rect 674703 273310 674814 273312
rect 674703 273254 674708 273310
rect 674764 273254 674814 273310
rect 674703 273249 674814 273254
rect 86031 273164 86097 273167
rect 376335 273164 376401 273167
rect 86031 273162 376401 273164
rect 86031 273106 86036 273162
rect 86092 273106 376340 273162
rect 376396 273106 376401 273162
rect 86031 273104 376401 273106
rect 86031 273101 86097 273104
rect 376335 273101 376401 273104
rect 376527 273164 376593 273167
rect 379311 273164 379377 273167
rect 384399 273164 384465 273167
rect 376527 273162 379377 273164
rect 376527 273106 376532 273162
rect 376588 273106 379316 273162
rect 379372 273106 379377 273162
rect 376527 273104 379377 273106
rect 376527 273101 376593 273104
rect 379311 273101 379377 273104
rect 379458 273162 384465 273164
rect 379458 273106 384404 273162
rect 384460 273106 384465 273162
rect 379458 273104 384465 273106
rect 41530 272954 41536 273018
rect 41600 273016 41606 273018
rect 41775 273016 41841 273019
rect 41600 273014 41841 273016
rect 41600 272958 41780 273014
rect 41836 272958 41841 273014
rect 41600 272956 41841 272958
rect 41600 272954 41606 272956
rect 41775 272953 41841 272956
rect 81327 273016 81393 273019
rect 378927 273016 378993 273019
rect 81327 273014 378993 273016
rect 81327 272958 81332 273014
rect 81388 272958 378932 273014
rect 378988 272958 378993 273014
rect 81327 272956 378993 272958
rect 81327 272953 81393 272956
rect 378927 272953 378993 272956
rect 379215 273016 379281 273019
rect 379458 273016 379518 273104
rect 384399 273101 384465 273104
rect 384634 273102 384640 273166
rect 384704 273164 384710 273166
rect 384783 273164 384849 273167
rect 384704 273162 384849 273164
rect 384704 273106 384788 273162
rect 384844 273106 384849 273162
rect 384704 273104 384849 273106
rect 384704 273102 384710 273104
rect 384783 273101 384849 273104
rect 389679 273164 389745 273167
rect 394671 273164 394737 273167
rect 389679 273162 394737 273164
rect 389679 273106 389684 273162
rect 389740 273106 394676 273162
rect 394732 273106 394737 273162
rect 389679 273104 394737 273106
rect 389679 273101 389745 273104
rect 394671 273101 394737 273104
rect 674754 273060 674814 273249
rect 379215 273014 379518 273016
rect 379215 272958 379220 273014
rect 379276 272958 379518 273014
rect 379215 272956 379518 272958
rect 379215 272953 379281 272956
rect 379642 272954 379648 273018
rect 379712 273016 379718 273018
rect 395343 273016 395409 273019
rect 379712 273014 395409 273016
rect 379712 272958 395348 273014
rect 395404 272958 395409 273014
rect 379712 272956 395409 272958
rect 379712 272954 379718 272956
rect 395343 272953 395409 272956
rect 71727 272868 71793 272871
rect 213039 272868 213105 272871
rect 71727 272866 213105 272868
rect 71727 272810 71732 272866
rect 71788 272810 213044 272866
rect 213100 272810 213105 272866
rect 71727 272808 213105 272810
rect 71727 272805 71793 272808
rect 213039 272805 213105 272808
rect 237519 272868 237585 272871
rect 260079 272868 260145 272871
rect 566511 272868 566577 272871
rect 237519 272866 248382 272868
rect 237519 272810 237524 272866
rect 237580 272810 248382 272866
rect 237519 272808 248382 272810
rect 237519 272805 237585 272808
rect 78927 272720 78993 272723
rect 156687 272720 156753 272723
rect 78927 272718 156753 272720
rect 78927 272662 78932 272718
rect 78988 272662 156692 272718
rect 156748 272662 156753 272718
rect 78927 272660 156753 272662
rect 78927 272657 78993 272660
rect 156687 272657 156753 272660
rect 156879 272720 156945 272723
rect 177039 272720 177105 272723
rect 156879 272718 177105 272720
rect 156879 272662 156884 272718
rect 156940 272662 177044 272718
rect 177100 272662 177105 272718
rect 156879 272660 177105 272662
rect 156879 272657 156945 272660
rect 177039 272657 177105 272660
rect 177231 272720 177297 272723
rect 197199 272720 197265 272723
rect 177231 272718 197265 272720
rect 177231 272662 177236 272718
rect 177292 272662 197204 272718
rect 197260 272662 197265 272718
rect 177231 272660 197265 272662
rect 177231 272657 177297 272660
rect 197199 272657 197265 272660
rect 197434 272658 197440 272722
rect 197504 272720 197510 272722
rect 248175 272720 248241 272723
rect 197504 272718 248241 272720
rect 197504 272662 248180 272718
rect 248236 272662 248241 272718
rect 197504 272660 248241 272662
rect 248322 272720 248382 272808
rect 260079 272866 566577 272868
rect 260079 272810 260084 272866
rect 260140 272810 566516 272866
rect 566572 272810 566577 272866
rect 260079 272808 566577 272810
rect 260079 272805 260145 272808
rect 566511 272805 566577 272808
rect 674938 272806 674944 272870
rect 675008 272806 675014 272870
rect 368655 272720 368721 272723
rect 248322 272718 368721 272720
rect 248322 272662 368660 272718
rect 368716 272662 368721 272718
rect 248322 272660 368721 272662
rect 197504 272658 197510 272660
rect 248175 272657 248241 272660
rect 368655 272657 368721 272660
rect 368847 272720 368913 272723
rect 563055 272720 563121 272723
rect 368847 272718 563121 272720
rect 368847 272662 368852 272718
rect 368908 272662 563060 272718
rect 563116 272662 563121 272718
rect 368847 272660 563121 272662
rect 368847 272657 368913 272660
rect 563055 272657 563121 272660
rect 76527 272572 76593 272575
rect 383535 272572 383601 272575
rect 76527 272570 383601 272572
rect 76527 272514 76532 272570
rect 76588 272514 383540 272570
rect 383596 272514 383601 272570
rect 76527 272512 383601 272514
rect 76527 272509 76593 272512
rect 383535 272509 383601 272512
rect 383919 272572 383985 272575
rect 387087 272572 387153 272575
rect 383919 272570 387153 272572
rect 383919 272514 383924 272570
rect 383980 272514 387092 272570
rect 387148 272514 387153 272570
rect 383919 272512 387153 272514
rect 383919 272509 383985 272512
rect 387087 272509 387153 272512
rect 389007 272572 389073 272575
rect 389967 272572 390033 272575
rect 389007 272570 390033 272572
rect 389007 272514 389012 272570
rect 389068 272514 389972 272570
rect 390028 272514 390033 272570
rect 389007 272512 390033 272514
rect 389007 272509 389073 272512
rect 389967 272509 390033 272512
rect 70575 272424 70641 272427
rect 381615 272424 381681 272427
rect 70575 272422 381681 272424
rect 70575 272366 70580 272422
rect 70636 272366 381620 272422
rect 381676 272366 381681 272422
rect 70575 272364 381681 272366
rect 70575 272361 70641 272364
rect 381615 272361 381681 272364
rect 381807 272424 381873 272427
rect 386127 272424 386193 272427
rect 381807 272422 386193 272424
rect 381807 272366 381812 272422
rect 381868 272366 386132 272422
rect 386188 272366 386193 272422
rect 381807 272364 386193 272366
rect 381807 272361 381873 272364
rect 386127 272361 386193 272364
rect 386607 272424 386673 272427
rect 405370 272424 405376 272426
rect 386607 272422 405376 272424
rect 386607 272366 386612 272422
rect 386668 272366 405376 272422
rect 386607 272364 405376 272366
rect 386607 272361 386673 272364
rect 405370 272362 405376 272364
rect 405440 272362 405446 272426
rect 41146 272214 41152 272278
rect 41216 272276 41222 272278
rect 41775 272276 41841 272279
rect 41216 272274 41841 272276
rect 41216 272218 41780 272274
rect 41836 272218 41841 272274
rect 41216 272216 41841 272218
rect 41216 272214 41222 272216
rect 41775 272213 41841 272216
rect 69423 272276 69489 272279
rect 374991 272276 375057 272279
rect 379311 272276 379377 272279
rect 69423 272274 374910 272276
rect 69423 272218 69428 272274
rect 69484 272218 374910 272274
rect 69423 272216 374910 272218
rect 69423 272213 69489 272216
rect 74127 272128 74193 272131
rect 374850 272128 374910 272216
rect 374991 272274 379377 272276
rect 374991 272218 374996 272274
rect 375052 272218 379316 272274
rect 379372 272218 379377 272274
rect 374991 272216 379377 272218
rect 374991 272213 375057 272216
rect 379311 272213 379377 272216
rect 379450 272214 379456 272278
rect 379520 272276 379526 272278
rect 379791 272276 379857 272279
rect 379520 272274 379857 272276
rect 379520 272218 379796 272274
rect 379852 272218 379857 272274
rect 379520 272216 379857 272218
rect 379520 272214 379526 272216
rect 379791 272213 379857 272216
rect 380175 272276 380241 272279
rect 573711 272276 573777 272279
rect 380175 272274 573777 272276
rect 380175 272218 380180 272274
rect 380236 272218 573716 272274
rect 573772 272218 573777 272274
rect 674946 272246 675006 272806
rect 380175 272216 573777 272218
rect 380175 272213 380241 272216
rect 573711 272213 573777 272216
rect 381807 272128 381873 272131
rect 74127 272126 374718 272128
rect 74127 272070 74132 272126
rect 74188 272070 374718 272126
rect 74127 272068 374718 272070
rect 374850 272126 381873 272128
rect 374850 272070 381812 272126
rect 381868 272070 381873 272126
rect 374850 272068 381873 272070
rect 74127 272065 74193 272068
rect 93231 271980 93297 271983
rect 374511 271980 374577 271983
rect 93231 271978 374577 271980
rect 93231 271922 93236 271978
rect 93292 271922 374516 271978
rect 374572 271922 374577 271978
rect 93231 271920 374577 271922
rect 374658 271980 374718 272068
rect 381807 272065 381873 272068
rect 383343 272128 383409 272131
rect 384879 272128 384945 272131
rect 383343 272126 384945 272128
rect 383343 272070 383348 272126
rect 383404 272070 384884 272126
rect 384940 272070 384945 272126
rect 383343 272068 384945 272070
rect 383343 272065 383409 272068
rect 384879 272065 384945 272068
rect 383439 271980 383505 271983
rect 374658 271978 383505 271980
rect 374658 271922 383444 271978
rect 383500 271922 383505 271978
rect 374658 271920 383505 271922
rect 93231 271917 93297 271920
rect 374511 271917 374577 271920
rect 383439 271917 383505 271920
rect 383631 271980 383697 271983
rect 385551 271980 385617 271983
rect 383631 271978 385617 271980
rect 383631 271922 383636 271978
rect 383692 271922 385556 271978
rect 385612 271922 385617 271978
rect 383631 271920 385617 271922
rect 383631 271917 383697 271920
rect 385551 271917 385617 271920
rect 96783 271832 96849 271835
rect 389199 271832 389265 271835
rect 96783 271830 389265 271832
rect 96783 271774 96788 271830
rect 96844 271774 389204 271830
rect 389260 271774 389265 271830
rect 96783 271772 389265 271774
rect 96783 271769 96849 271772
rect 389199 271769 389265 271772
rect 391407 271832 391473 271835
rect 404218 271832 404224 271834
rect 391407 271830 404224 271832
rect 391407 271774 391412 271830
rect 391468 271774 404224 271830
rect 391407 271772 404224 271774
rect 391407 271769 391473 271772
rect 404218 271770 404224 271772
rect 404288 271770 404294 271834
rect 90831 271684 90897 271687
rect 116559 271684 116625 271687
rect 90831 271682 116625 271684
rect 90831 271626 90836 271682
rect 90892 271626 116564 271682
rect 116620 271626 116625 271682
rect 90831 271624 116625 271626
rect 90831 271621 90897 271624
rect 116559 271621 116625 271624
rect 121743 271684 121809 271687
rect 146895 271684 146961 271687
rect 121743 271682 146961 271684
rect 121743 271626 121748 271682
rect 121804 271626 146900 271682
rect 146956 271626 146961 271682
rect 121743 271624 146961 271626
rect 121743 271621 121809 271624
rect 146895 271621 146961 271624
rect 147087 271684 147153 271687
rect 157167 271684 157233 271687
rect 147087 271682 157233 271684
rect 147087 271626 147092 271682
rect 147148 271626 157172 271682
rect 157228 271626 157233 271682
rect 147087 271624 157233 271626
rect 147087 271621 147153 271624
rect 157167 271621 157233 271624
rect 166767 271684 166833 271687
rect 187215 271684 187281 271687
rect 166767 271682 187281 271684
rect 166767 271626 166772 271682
rect 166828 271626 187220 271682
rect 187276 271626 187281 271682
rect 166767 271624 187281 271626
rect 166767 271621 166833 271624
rect 187215 271621 187281 271624
rect 207279 271684 207345 271687
rect 227535 271684 227601 271687
rect 207279 271682 227601 271684
rect 207279 271626 207284 271682
rect 207340 271626 227540 271682
rect 227596 271626 227601 271682
rect 207279 271624 227601 271626
rect 207279 271621 207345 271624
rect 227535 271621 227601 271624
rect 247599 271684 247665 271687
rect 267855 271684 267921 271687
rect 247599 271682 267921 271684
rect 247599 271626 247604 271682
rect 247660 271626 267860 271682
rect 267916 271626 267921 271682
rect 247599 271624 267921 271626
rect 247599 271621 247665 271624
rect 267855 271621 267921 271624
rect 302415 271684 302481 271687
rect 324154 271684 324160 271686
rect 302415 271682 324160 271684
rect 302415 271626 302420 271682
rect 302476 271626 324160 271682
rect 302415 271624 324160 271626
rect 302415 271621 302481 271624
rect 324154 271622 324160 271624
rect 324224 271622 324230 271686
rect 324399 271684 324465 271687
rect 328815 271684 328881 271687
rect 324399 271682 328881 271684
rect 324399 271626 324404 271682
rect 324460 271626 328820 271682
rect 328876 271626 328881 271682
rect 324399 271624 328881 271626
rect 324399 271621 324465 271624
rect 328815 271621 328881 271624
rect 329007 271684 329073 271687
rect 379066 271684 379072 271686
rect 329007 271682 379072 271684
rect 329007 271626 329012 271682
rect 329068 271626 379072 271682
rect 329007 271624 379072 271626
rect 329007 271621 329073 271624
rect 379066 271622 379072 271624
rect 379136 271622 379142 271686
rect 379311 271684 379377 271687
rect 388047 271684 388113 271687
rect 379311 271682 388113 271684
rect 379311 271626 379316 271682
rect 379372 271626 388052 271682
rect 388108 271626 388113 271682
rect 379311 271624 388113 271626
rect 379311 271621 379377 271624
rect 388047 271621 388113 271624
rect 388623 271684 388689 271687
rect 388911 271684 388977 271687
rect 388623 271682 388977 271684
rect 388623 271626 388628 271682
rect 388684 271626 388916 271682
rect 388972 271626 388977 271682
rect 388623 271624 388977 271626
rect 388623 271621 388689 271624
rect 388911 271621 388977 271624
rect 390831 271684 390897 271687
rect 403834 271684 403840 271686
rect 390831 271682 403840 271684
rect 390831 271626 390836 271682
rect 390892 271626 403840 271682
rect 390831 271624 403840 271626
rect 390831 271621 390897 271624
rect 403834 271622 403840 271624
rect 403904 271622 403910 271686
rect 91983 271536 92049 271539
rect 270639 271536 270705 271539
rect 91983 271534 270705 271536
rect 91983 271478 91988 271534
rect 92044 271478 270644 271534
rect 270700 271478 270705 271534
rect 91983 271476 270705 271478
rect 91983 271473 92049 271476
rect 270639 271473 270705 271476
rect 315759 271536 315825 271539
rect 324975 271536 325041 271539
rect 315759 271534 325041 271536
rect 315759 271478 315764 271534
rect 315820 271478 324980 271534
rect 325036 271478 325041 271534
rect 315759 271476 325041 271478
rect 315759 271473 315825 271476
rect 324975 271473 325041 271476
rect 325359 271536 325425 271539
rect 356986 271536 356992 271538
rect 325359 271534 356992 271536
rect 325359 271478 325364 271534
rect 325420 271478 356992 271534
rect 325359 271476 356992 271478
rect 325359 271473 325425 271476
rect 356986 271474 356992 271476
rect 357056 271474 357062 271538
rect 370959 271536 371025 271539
rect 369282 271534 371025 271536
rect 369282 271478 370964 271534
rect 371020 271478 371025 271534
rect 369282 271476 371025 271478
rect 87183 271388 87249 271391
rect 211791 271388 211857 271391
rect 237519 271388 237585 271391
rect 87183 271386 211857 271388
rect 87183 271330 87188 271386
rect 87244 271330 211796 271386
rect 211852 271330 211857 271386
rect 87183 271328 211857 271330
rect 87183 271325 87249 271328
rect 211791 271325 211857 271328
rect 217218 271386 237585 271388
rect 217218 271330 237524 271386
rect 237580 271330 237585 271386
rect 217218 271328 237585 271330
rect 95631 271240 95697 271243
rect 211983 271240 212049 271243
rect 95631 271238 212049 271240
rect 95631 271182 95636 271238
rect 95692 271182 211988 271238
rect 212044 271182 212049 271238
rect 95631 271180 212049 271182
rect 95631 271177 95697 271180
rect 211983 271177 212049 271180
rect 156687 271092 156753 271095
rect 177231 271092 177297 271095
rect 156687 271090 177297 271092
rect 156687 271034 156692 271090
rect 156748 271034 177236 271090
rect 177292 271034 177297 271090
rect 156687 271032 177297 271034
rect 156687 271029 156753 271032
rect 177231 271029 177297 271032
rect 177423 271092 177489 271095
rect 197050 271092 197056 271094
rect 177423 271090 197056 271092
rect 177423 271034 177428 271090
rect 177484 271034 197056 271090
rect 177423 271032 197056 271034
rect 177423 271029 177489 271032
rect 197050 271030 197056 271032
rect 197120 271030 197126 271094
rect 197199 271092 197265 271095
rect 217218 271092 217278 271328
rect 237519 271325 237585 271328
rect 237711 271388 237777 271391
rect 250575 271388 250641 271391
rect 237711 271386 250641 271388
rect 237711 271330 237716 271386
rect 237772 271330 250580 271386
rect 250636 271330 250641 271386
rect 237711 271328 250641 271330
rect 237711 271325 237777 271328
rect 250575 271325 250641 271328
rect 267855 271388 267921 271391
rect 322479 271388 322545 271391
rect 267855 271386 322545 271388
rect 267855 271330 267860 271386
rect 267916 271330 322484 271386
rect 322540 271330 322545 271386
rect 267855 271328 322545 271330
rect 267855 271325 267921 271328
rect 322479 271325 322545 271328
rect 323247 271388 323313 271391
rect 336975 271388 337041 271391
rect 323247 271386 337041 271388
rect 323247 271330 323252 271386
rect 323308 271330 336980 271386
rect 337036 271330 337041 271386
rect 323247 271328 337041 271330
rect 323247 271325 323313 271328
rect 336975 271325 337041 271328
rect 363759 271388 363825 271391
rect 369282 271388 369342 271476
rect 370959 271473 371025 271476
rect 371439 271536 371505 271539
rect 559407 271536 559473 271539
rect 371439 271534 559473 271536
rect 371439 271478 371444 271534
rect 371500 271478 559412 271534
rect 559468 271478 559473 271534
rect 371439 271476 559473 271478
rect 371439 271473 371505 271476
rect 559407 271473 559473 271476
rect 363759 271386 369342 271388
rect 363759 271330 363764 271386
rect 363820 271330 369342 271386
rect 363759 271328 369342 271330
rect 370575 271388 370641 271391
rect 555855 271388 555921 271391
rect 370575 271386 555921 271388
rect 370575 271330 370580 271386
rect 370636 271330 555860 271386
rect 555916 271330 555921 271386
rect 370575 271328 555921 271330
rect 363759 271325 363825 271328
rect 370575 271325 370641 271328
rect 555855 271325 555921 271328
rect 237615 271240 237681 271243
rect 257679 271240 257745 271243
rect 237615 271238 257745 271240
rect 237615 271182 237620 271238
rect 237676 271182 257684 271238
rect 257740 271182 257745 271238
rect 237615 271180 257745 271182
rect 237615 271177 237681 271180
rect 257679 271177 257745 271180
rect 322575 271240 322641 271243
rect 327951 271240 328017 271243
rect 322575 271238 328017 271240
rect 322575 271182 322580 271238
rect 322636 271182 327956 271238
rect 328012 271182 328017 271238
rect 322575 271180 328017 271182
rect 322575 271177 322641 271180
rect 327951 271177 328017 271180
rect 328143 271240 328209 271243
rect 330831 271240 330897 271243
rect 328143 271238 330897 271240
rect 328143 271182 328148 271238
rect 328204 271182 330836 271238
rect 330892 271182 330897 271238
rect 328143 271180 330897 271182
rect 328143 271177 328209 271180
rect 330831 271177 330897 271180
rect 331066 271178 331072 271242
rect 331136 271240 331142 271242
rect 339759 271240 339825 271243
rect 552303 271240 552369 271243
rect 331136 271238 339825 271240
rect 331136 271182 339764 271238
rect 339820 271182 339825 271238
rect 331136 271180 339825 271182
rect 331136 271178 331142 271180
rect 339759 271177 339825 271180
rect 368754 271238 552369 271240
rect 368754 271182 552308 271238
rect 552364 271182 552369 271238
rect 368754 271180 552369 271182
rect 197199 271090 217278 271092
rect 197199 271034 197204 271090
rect 197260 271034 217278 271090
rect 197199 271032 217278 271034
rect 227535 271092 227601 271095
rect 247599 271092 247665 271095
rect 227535 271090 247665 271092
rect 227535 271034 227540 271090
rect 227596 271034 247604 271090
rect 247660 271034 247665 271090
rect 227535 271032 247665 271034
rect 197199 271029 197265 271032
rect 227535 271029 227601 271032
rect 247599 271029 247665 271032
rect 261135 271092 261201 271095
rect 325455 271092 325521 271095
rect 261135 271090 325521 271092
rect 261135 271034 261140 271090
rect 261196 271034 325460 271090
rect 325516 271034 325521 271090
rect 261135 271032 325521 271034
rect 261135 271029 261201 271032
rect 325455 271029 325521 271032
rect 325647 271092 325713 271095
rect 328623 271092 328689 271095
rect 325647 271090 328689 271092
rect 325647 271034 325652 271090
rect 325708 271034 328628 271090
rect 328684 271034 328689 271090
rect 325647 271032 328689 271034
rect 325647 271029 325713 271032
rect 328623 271029 328689 271032
rect 328815 271092 328881 271095
rect 342447 271092 342513 271095
rect 328815 271090 342513 271092
rect 328815 271034 328820 271090
rect 328876 271034 342452 271090
rect 342508 271034 342513 271090
rect 328815 271032 342513 271034
rect 328815 271029 328881 271032
rect 342447 271029 342513 271032
rect 368175 271092 368241 271095
rect 368754 271092 368814 271180
rect 552303 271177 552369 271180
rect 368175 271090 368814 271092
rect 368175 271034 368180 271090
rect 368236 271034 368814 271090
rect 368175 271032 368814 271034
rect 369807 271092 369873 271095
rect 548751 271092 548817 271095
rect 369807 271090 548817 271092
rect 369807 271034 369812 271090
rect 369868 271034 548756 271090
rect 548812 271034 548817 271090
rect 369807 271032 548817 271034
rect 368175 271029 368241 271032
rect 369807 271029 369873 271032
rect 548751 271029 548817 271032
rect 156975 270944 157041 270947
rect 177711 270944 177777 270947
rect 156975 270942 177777 270944
rect 156975 270886 156980 270942
rect 157036 270886 177716 270942
rect 177772 270886 177777 270942
rect 156975 270884 177777 270886
rect 156975 270881 157041 270884
rect 177711 270881 177777 270884
rect 197583 270944 197649 270947
rect 217359 270944 217425 270947
rect 197583 270942 217425 270944
rect 197583 270886 197588 270942
rect 197644 270886 217364 270942
rect 217420 270886 217425 270942
rect 197583 270884 217425 270886
rect 197583 270881 197649 270884
rect 217359 270881 217425 270884
rect 264879 270944 264945 270947
rect 351279 270944 351345 270947
rect 264879 270942 351345 270944
rect 264879 270886 264884 270942
rect 264940 270886 351284 270942
rect 351340 270886 351345 270942
rect 264879 270884 351345 270886
rect 264879 270881 264945 270884
rect 351279 270881 351345 270884
rect 356943 270944 357009 270947
rect 371439 270944 371505 270947
rect 356943 270942 371505 270944
rect 356943 270886 356948 270942
rect 357004 270886 371444 270942
rect 371500 270886 371505 270942
rect 356943 270884 371505 270886
rect 356943 270881 357009 270884
rect 371439 270881 371505 270884
rect 376623 270944 376689 270947
rect 386031 270944 386097 270947
rect 376623 270942 386097 270944
rect 376623 270886 376628 270942
rect 376684 270886 386036 270942
rect 386092 270886 386097 270942
rect 376623 270884 386097 270886
rect 376623 270881 376689 270884
rect 386031 270881 386097 270884
rect 387130 270882 387136 270946
rect 387200 270944 387206 270946
rect 401583 270944 401649 270947
rect 387200 270942 401649 270944
rect 387200 270886 401588 270942
rect 401644 270886 401649 270942
rect 387200 270884 401649 270886
rect 387200 270882 387206 270884
rect 401583 270881 401649 270884
rect 673978 270882 673984 270946
rect 674048 270944 674054 270946
rect 674754 270944 674814 271432
rect 674048 270884 674814 270944
rect 674048 270882 674054 270884
rect 146895 270796 146961 270799
rect 166767 270796 166833 270799
rect 146895 270794 166833 270796
rect 146895 270738 146900 270794
rect 146956 270738 166772 270794
rect 166828 270738 166833 270794
rect 146895 270736 166833 270738
rect 146895 270733 146961 270736
rect 166767 270733 166833 270736
rect 194511 270796 194577 270799
rect 212559 270796 212625 270799
rect 194511 270794 212625 270796
rect 194511 270738 194516 270794
rect 194572 270738 212564 270794
rect 212620 270738 212625 270794
rect 194511 270736 212625 270738
rect 194511 270733 194577 270736
rect 212559 270733 212625 270736
rect 212751 270796 212817 270799
rect 355215 270796 355281 270799
rect 212751 270794 355281 270796
rect 212751 270738 212756 270794
rect 212812 270738 355220 270794
rect 355276 270738 355281 270794
rect 212751 270736 355281 270738
rect 212751 270733 212817 270736
rect 355215 270733 355281 270736
rect 368367 270796 368433 270799
rect 368751 270796 368817 270799
rect 368367 270794 368817 270796
rect 368367 270738 368372 270794
rect 368428 270738 368756 270794
rect 368812 270738 368817 270794
rect 368367 270736 368817 270738
rect 368367 270733 368433 270736
rect 368751 270733 368817 270736
rect 368943 270796 369009 270799
rect 373167 270796 373233 270799
rect 368943 270794 373233 270796
rect 368943 270738 368948 270794
rect 369004 270738 373172 270794
rect 373228 270738 373233 270794
rect 368943 270736 373233 270738
rect 368943 270733 369009 270736
rect 373167 270733 373233 270736
rect 373551 270796 373617 270799
rect 383919 270796 383985 270799
rect 373551 270794 383985 270796
rect 373551 270738 373556 270794
rect 373612 270738 383924 270794
rect 383980 270738 383985 270794
rect 373551 270736 383985 270738
rect 373551 270733 373617 270736
rect 383919 270733 383985 270736
rect 384058 270734 384064 270798
rect 384128 270796 384134 270798
rect 387567 270796 387633 270799
rect 384128 270794 387633 270796
rect 384128 270738 387572 270794
rect 387628 270738 387633 270794
rect 384128 270736 387633 270738
rect 384128 270734 384134 270736
rect 387567 270733 387633 270736
rect 387759 270796 387825 270799
rect 394575 270796 394641 270799
rect 387759 270794 394641 270796
rect 387759 270738 387764 270794
rect 387820 270738 394580 270794
rect 394636 270738 394641 270794
rect 387759 270736 394641 270738
rect 387759 270733 387825 270736
rect 394575 270733 394641 270736
rect 395823 270796 395889 270799
rect 404026 270796 404032 270798
rect 395823 270794 404032 270796
rect 395823 270738 395828 270794
rect 395884 270738 404032 270794
rect 395823 270736 404032 270738
rect 395823 270733 395889 270736
rect 404026 270734 404032 270736
rect 404096 270734 404102 270798
rect 647535 270796 647601 270799
rect 639426 270794 647601 270796
rect 639426 270738 647540 270794
rect 647596 270738 647601 270794
rect 639426 270736 647601 270738
rect 40762 270586 40768 270650
rect 40832 270648 40838 270650
rect 41775 270648 41841 270651
rect 40832 270646 41841 270648
rect 40832 270590 41780 270646
rect 41836 270590 41841 270646
rect 40832 270588 41841 270590
rect 40832 270586 40838 270588
rect 41775 270585 41841 270588
rect 256431 270648 256497 270651
rect 276303 270648 276369 270651
rect 256431 270646 276369 270648
rect 256431 270590 256436 270646
rect 256492 270590 276308 270646
rect 276364 270590 276369 270646
rect 256431 270588 276369 270590
rect 256431 270585 256497 270588
rect 276303 270585 276369 270588
rect 312111 270648 312177 270651
rect 320559 270648 320625 270651
rect 312111 270646 320625 270648
rect 312111 270590 312116 270646
rect 312172 270590 320564 270646
rect 320620 270590 320625 270646
rect 312111 270588 320625 270590
rect 312111 270585 312177 270588
rect 320559 270585 320625 270588
rect 322479 270648 322545 270651
rect 328047 270648 328113 270651
rect 322479 270646 328113 270648
rect 322479 270590 322484 270646
rect 322540 270590 328052 270646
rect 328108 270590 328113 270646
rect 322479 270588 328113 270590
rect 322479 270585 322545 270588
rect 328047 270585 328113 270588
rect 328623 270648 328689 270651
rect 582063 270648 582129 270651
rect 328623 270646 582129 270648
rect 328623 270590 328628 270646
rect 328684 270590 582068 270646
rect 582124 270590 582129 270646
rect 328623 270588 582129 270590
rect 328623 270585 328689 270588
rect 582063 270585 582129 270588
rect 41722 270438 41728 270502
rect 41792 270500 41798 270502
rect 42543 270500 42609 270503
rect 41792 270498 42609 270500
rect 41792 270442 42548 270498
rect 42604 270442 42609 270498
rect 41792 270440 42609 270442
rect 41792 270438 41798 270440
rect 42543 270437 42609 270440
rect 257871 270500 257937 270503
rect 369807 270500 369873 270503
rect 257871 270498 369873 270500
rect 257871 270442 257876 270498
rect 257932 270442 369812 270498
rect 369868 270442 369873 270498
rect 257871 270440 369873 270442
rect 257871 270437 257937 270440
rect 369807 270437 369873 270440
rect 369999 270500 370065 270503
rect 388719 270500 388785 270503
rect 369999 270498 388785 270500
rect 369999 270442 370004 270498
rect 370060 270442 388724 270498
rect 388780 270442 388785 270498
rect 369999 270440 388785 270442
rect 369999 270437 370065 270440
rect 388719 270437 388785 270440
rect 388911 270500 388977 270503
rect 429135 270500 429201 270503
rect 388911 270498 429201 270500
rect 388911 270442 388916 270498
rect 388972 270442 429140 270498
rect 429196 270442 429201 270498
rect 388911 270440 429201 270442
rect 388911 270437 388977 270440
rect 429135 270437 429201 270440
rect 449199 270500 449265 270503
rect 469455 270500 469521 270503
rect 449199 270498 469521 270500
rect 449199 270442 449204 270498
rect 449260 270442 469460 270498
rect 469516 270442 469521 270498
rect 449199 270440 469521 270442
rect 449199 270437 449265 270440
rect 469455 270437 469521 270440
rect 489519 270500 489585 270503
rect 509775 270500 509841 270503
rect 489519 270498 509841 270500
rect 489519 270442 489524 270498
rect 489580 270442 509780 270498
rect 509836 270442 509841 270498
rect 489519 270440 509841 270442
rect 489519 270437 489585 270440
rect 509775 270437 509841 270440
rect 524367 270500 524433 270503
rect 552975 270500 553041 270503
rect 590415 270500 590481 270503
rect 524367 270498 553041 270500
rect 524367 270442 524372 270498
rect 524428 270442 552980 270498
rect 553036 270442 553041 270498
rect 524367 270440 553041 270442
rect 524367 270437 524433 270440
rect 552975 270437 553041 270440
rect 583170 270498 590481 270500
rect 583170 270442 590420 270498
rect 590476 270442 590481 270498
rect 583170 270440 590481 270442
rect 254607 270352 254673 270355
rect 523791 270352 523857 270355
rect 254607 270350 523857 270352
rect 254607 270294 254612 270350
rect 254668 270294 523796 270350
rect 523852 270294 523857 270350
rect 254607 270292 523857 270294
rect 254607 270289 254673 270292
rect 523791 270289 523857 270292
rect 573039 270352 573105 270355
rect 573186 270352 573630 270389
rect 583170 270352 583230 270440
rect 590415 270437 590481 270440
rect 600495 270500 600561 270503
rect 639426 270500 639486 270736
rect 647535 270733 647601 270736
rect 600495 270498 639486 270500
rect 600495 270442 600500 270498
rect 600556 270442 639486 270498
rect 600495 270440 639486 270442
rect 600495 270437 600561 270440
rect 573039 270350 583230 270352
rect 573039 270294 573044 270350
rect 573100 270329 583230 270350
rect 573100 270294 573246 270329
rect 573039 270292 573246 270294
rect 573570 270292 583230 270329
rect 573039 270289 573105 270292
rect 178575 270204 178641 270207
rect 195855 270204 195921 270207
rect 178575 270202 195921 270204
rect 178575 270146 178580 270202
rect 178636 270146 195860 270202
rect 195916 270146 195921 270202
rect 178575 270144 195921 270146
rect 178575 270141 178641 270144
rect 195855 270141 195921 270144
rect 276591 270204 276657 270207
rect 296559 270204 296625 270207
rect 276591 270202 296625 270204
rect 276591 270146 276596 270202
rect 276652 270146 296564 270202
rect 296620 270146 296625 270202
rect 276591 270144 296625 270146
rect 276591 270141 276657 270144
rect 296559 270141 296625 270144
rect 319119 270204 319185 270207
rect 336975 270204 337041 270207
rect 573135 270204 573201 270207
rect 319119 270202 330942 270204
rect 319119 270146 319124 270202
rect 319180 270146 330942 270202
rect 319119 270144 330942 270146
rect 319119 270141 319185 270144
rect 41338 269994 41344 270058
rect 41408 270056 41414 270058
rect 41775 270056 41841 270059
rect 41408 270054 41841 270056
rect 41408 269998 41780 270054
rect 41836 269998 41841 270054
rect 41408 269996 41841 269998
rect 41408 269994 41414 269996
rect 41775 269993 41841 269996
rect 195951 270056 196017 270059
rect 312879 270056 312945 270059
rect 317487 270056 317553 270059
rect 195951 270054 199038 270056
rect 195951 269998 195956 270054
rect 196012 269998 199038 270054
rect 195951 269996 199038 269998
rect 195951 269993 196017 269996
rect 118095 269908 118161 269911
rect 138106 269908 138112 269910
rect 118095 269906 138112 269908
rect 118095 269850 118100 269906
rect 118156 269850 138112 269906
rect 118095 269848 138112 269850
rect 118095 269845 118161 269848
rect 138106 269846 138112 269848
rect 138176 269846 138182 269910
rect 198978 269908 199038 269996
rect 312879 270054 317553 270056
rect 312879 269998 312884 270054
rect 312940 269998 317492 270054
rect 317548 269998 317553 270054
rect 312879 269996 317553 269998
rect 312879 269993 312945 269996
rect 317487 269993 317553 269996
rect 318735 270056 318801 270059
rect 323247 270056 323313 270059
rect 318735 270054 323313 270056
rect 318735 269998 318740 270054
rect 318796 269998 323252 270054
rect 323308 269998 323313 270054
rect 318735 269996 323313 269998
rect 318735 269993 318801 269996
rect 323247 269993 323313 269996
rect 323439 270056 323505 270059
rect 329007 270056 329073 270059
rect 323439 270054 329073 270056
rect 323439 269998 323444 270054
rect 323500 269998 329012 270054
rect 329068 269998 329073 270054
rect 323439 269996 329073 269998
rect 330882 270056 330942 270144
rect 336975 270202 573201 270204
rect 336975 270146 336980 270202
rect 337036 270146 573140 270202
rect 573196 270146 573201 270202
rect 336975 270144 573201 270146
rect 336975 270141 337041 270144
rect 573135 270141 573201 270144
rect 674170 270142 674176 270206
rect 674240 270204 674246 270206
rect 674754 270204 674814 270766
rect 674240 270144 674814 270204
rect 674240 270142 674246 270144
rect 596367 270056 596433 270059
rect 330882 270054 596433 270056
rect 330882 269998 596372 270054
rect 596428 269998 596433 270054
rect 330882 269996 596433 269998
rect 323439 269993 323505 269996
rect 329007 269993 329073 269996
rect 596367 269993 596433 269996
rect 216015 269908 216081 269911
rect 161154 269848 161406 269908
rect 198978 269906 216081 269908
rect 198978 269850 216020 269906
rect 216076 269850 216081 269906
rect 198978 269848 216081 269850
rect 141135 269760 141201 269763
rect 161154 269760 161214 269848
rect 141135 269758 161214 269760
rect 141135 269702 141140 269758
rect 141196 269702 161214 269758
rect 141135 269700 161214 269702
rect 161346 269760 161406 269848
rect 216015 269845 216081 269848
rect 243279 269908 243345 269911
rect 253359 269908 253425 269911
rect 243279 269906 253425 269908
rect 243279 269850 243284 269906
rect 243340 269850 253364 269906
rect 253420 269850 253425 269906
rect 243279 269848 253425 269850
rect 243279 269845 243345 269848
rect 253359 269845 253425 269848
rect 276303 269908 276369 269911
rect 276495 269908 276561 269911
rect 276303 269906 276561 269908
rect 276303 269850 276308 269906
rect 276364 269850 276500 269906
rect 276556 269850 276561 269906
rect 276303 269848 276561 269850
rect 276303 269845 276369 269848
rect 276495 269845 276561 269848
rect 296559 269908 296625 269911
rect 299487 269908 299553 269911
rect 296559 269906 299553 269908
rect 296559 269850 296564 269906
rect 296620 269850 299492 269906
rect 299548 269850 299553 269906
rect 296559 269848 299553 269850
rect 296559 269845 296625 269848
rect 299487 269845 299553 269848
rect 317487 269908 317553 269911
rect 324687 269908 324753 269911
rect 317487 269906 324753 269908
rect 317487 269850 317492 269906
rect 317548 269850 324692 269906
rect 324748 269850 324753 269906
rect 317487 269848 324753 269850
rect 317487 269845 317553 269848
rect 324687 269845 324753 269848
rect 327087 269908 327153 269911
rect 328431 269908 328497 269911
rect 327087 269906 328497 269908
rect 327087 269850 327092 269906
rect 327148 269850 328436 269906
rect 328492 269850 328497 269906
rect 327087 269848 328497 269850
rect 327087 269845 327153 269848
rect 328431 269845 328497 269848
rect 342543 269908 342609 269911
rect 383151 269908 383217 269911
rect 342543 269906 383217 269908
rect 342543 269850 342548 269906
rect 342604 269850 383156 269906
rect 383212 269850 383217 269906
rect 342543 269848 383217 269850
rect 342543 269845 342609 269848
rect 383151 269845 383217 269848
rect 403119 269908 403185 269911
rect 414735 269908 414801 269911
rect 403119 269906 414801 269908
rect 403119 269850 403124 269906
rect 403180 269850 414740 269906
rect 414796 269850 414801 269906
rect 403119 269848 414801 269850
rect 403119 269845 403185 269848
rect 414735 269845 414801 269848
rect 427599 269908 427665 269911
rect 437583 269908 437649 269911
rect 469359 269908 469425 269911
rect 427599 269906 437649 269908
rect 427599 269850 427604 269906
rect 427660 269850 437588 269906
rect 437644 269850 437649 269906
rect 427599 269848 437649 269850
rect 427599 269845 427665 269848
rect 437583 269845 437649 269848
rect 437826 269906 469425 269908
rect 437826 269850 469364 269906
rect 469420 269850 469425 269906
rect 437826 269848 469425 269850
rect 178575 269760 178641 269763
rect 161346 269758 178641 269760
rect 161346 269702 178580 269758
rect 178636 269702 178641 269758
rect 161346 269700 178641 269702
rect 141135 269697 141201 269700
rect 178575 269697 178641 269700
rect 253359 269758 253425 269763
rect 253359 269702 253364 269758
rect 253420 269702 253425 269758
rect 253359 269697 253425 269702
rect 299727 269760 299793 269763
rect 323002 269760 323008 269762
rect 299727 269758 323008 269760
rect 299727 269702 299732 269758
rect 299788 269702 323008 269758
rect 299727 269700 323008 269702
rect 299727 269697 299793 269700
rect 323002 269698 323008 269700
rect 323072 269698 323078 269762
rect 323151 269760 323217 269763
rect 336591 269760 336657 269763
rect 323151 269758 336657 269760
rect 323151 269702 323156 269758
rect 323212 269702 336596 269758
rect 336652 269702 336657 269758
rect 323151 269700 336657 269702
rect 323151 269697 323217 269700
rect 336591 269697 336657 269700
rect 342586 269698 342592 269762
rect 342656 269760 342662 269762
rect 368559 269760 368625 269763
rect 342656 269758 368625 269760
rect 342656 269702 368564 269758
rect 368620 269702 368625 269758
rect 342656 269700 368625 269702
rect 342656 269698 342662 269700
rect 368559 269697 368625 269700
rect 368751 269760 368817 269763
rect 380175 269760 380241 269763
rect 368751 269758 380241 269760
rect 368751 269702 368756 269758
rect 368812 269702 380180 269758
rect 380236 269702 380241 269758
rect 368751 269700 380241 269702
rect 368751 269697 368817 269700
rect 380175 269697 380241 269700
rect 380559 269760 380625 269763
rect 398895 269760 398961 269763
rect 380559 269758 398961 269760
rect 380559 269702 380564 269758
rect 380620 269702 398900 269758
rect 398956 269702 398961 269758
rect 380559 269700 398961 269702
rect 380559 269697 380625 269700
rect 398895 269697 398961 269700
rect 399034 269698 399040 269762
rect 399104 269760 399110 269762
rect 406095 269760 406161 269763
rect 399104 269758 406161 269760
rect 399104 269702 406100 269758
rect 406156 269702 406161 269758
rect 399104 269700 406161 269702
rect 399104 269698 399110 269700
rect 406095 269697 406161 269700
rect 434799 269760 434865 269763
rect 437826 269760 437886 269848
rect 469359 269845 469425 269848
rect 469551 269908 469617 269911
rect 489423 269908 489489 269911
rect 469551 269906 489489 269908
rect 469551 269850 469556 269906
rect 469612 269850 489428 269906
rect 489484 269850 489489 269906
rect 469551 269848 489489 269850
rect 469551 269845 469617 269848
rect 489423 269845 489489 269848
rect 529935 269908 530001 269911
rect 552975 269908 553041 269911
rect 529935 269906 553041 269908
rect 529935 269850 529940 269906
rect 529996 269850 552980 269906
rect 553036 269850 553041 269906
rect 529935 269848 553041 269850
rect 529935 269845 530001 269848
rect 552975 269845 553041 269848
rect 434799 269758 437886 269760
rect 434799 269702 434804 269758
rect 434860 269702 437886 269758
rect 434799 269700 437886 269702
rect 457935 269760 458001 269763
rect 458607 269760 458673 269763
rect 457935 269758 458673 269760
rect 457935 269702 457940 269758
rect 457996 269702 458612 269758
rect 458668 269702 458673 269758
rect 457935 269700 458673 269702
rect 434799 269697 434865 269700
rect 457935 269697 458001 269700
rect 458607 269697 458673 269700
rect 469455 269760 469521 269763
rect 483855 269760 483921 269763
rect 469455 269758 483921 269760
rect 469455 269702 469460 269758
rect 469516 269702 483860 269758
rect 483916 269702 483921 269758
rect 469455 269700 483921 269702
rect 469455 269697 469521 269700
rect 483855 269697 483921 269700
rect 518319 269760 518385 269763
rect 529839 269760 529905 269763
rect 518319 269758 529905 269760
rect 518319 269702 518324 269758
rect 518380 269702 529844 269758
rect 529900 269702 529905 269758
rect 518319 269700 529905 269702
rect 518319 269697 518385 269700
rect 529839 269697 529905 269700
rect 553071 269760 553137 269763
rect 593199 269760 593265 269763
rect 610575 269760 610641 269763
rect 675138 269762 675198 269878
rect 553071 269758 570366 269760
rect 553071 269702 553076 269758
rect 553132 269702 570366 269758
rect 553071 269700 570366 269702
rect 553071 269697 553137 269700
rect 77775 269612 77841 269615
rect 85263 269612 85329 269615
rect 77775 269610 85329 269612
rect 77775 269554 77780 269610
rect 77836 269554 85268 269610
rect 85324 269554 85329 269610
rect 77775 269552 85329 269554
rect 77775 269549 77841 269552
rect 85263 269549 85329 269552
rect 138106 269550 138112 269614
rect 138176 269612 138182 269614
rect 141135 269612 141201 269615
rect 138176 269610 141201 269612
rect 138176 269554 141140 269610
rect 141196 269554 141201 269610
rect 138176 269552 141201 269554
rect 253362 269612 253422 269697
rect 260559 269612 260625 269615
rect 483855 269612 483921 269615
rect 253362 269552 256398 269612
rect 138176 269550 138182 269552
rect 141135 269549 141201 269552
rect 256338 269467 256398 269552
rect 260559 269610 483921 269612
rect 260559 269554 260564 269610
rect 260620 269554 483860 269610
rect 483916 269554 483921 269610
rect 260559 269552 483921 269554
rect 260559 269549 260625 269552
rect 483855 269549 483921 269552
rect 484143 269612 484209 269615
rect 570159 269612 570225 269615
rect 484143 269610 570225 269612
rect 484143 269554 484148 269610
rect 484204 269554 570164 269610
rect 570220 269554 570225 269610
rect 484143 269552 570225 269554
rect 570306 269612 570366 269700
rect 593199 269758 610641 269760
rect 593199 269702 593204 269758
rect 593260 269702 610580 269758
rect 610636 269702 610641 269758
rect 593199 269700 610641 269702
rect 593199 269697 593265 269700
rect 610575 269697 610641 269700
rect 674554 269698 674560 269762
rect 674624 269760 674630 269762
rect 675130 269760 675136 269762
rect 674624 269700 675136 269760
rect 674624 269698 674630 269700
rect 675130 269698 675136 269700
rect 675200 269698 675206 269762
rect 573135 269612 573201 269615
rect 570306 269610 573201 269612
rect 570306 269554 573140 269610
rect 573196 269554 573201 269610
rect 570306 269552 573201 269554
rect 484143 269549 484209 269552
rect 570159 269549 570225 269552
rect 573135 269549 573201 269552
rect 86511 269464 86577 269467
rect 106426 269464 106432 269466
rect 86511 269462 106432 269464
rect 86511 269406 86516 269462
rect 86572 269406 106432 269462
rect 86511 269404 106432 269406
rect 86511 269401 86577 269404
rect 106426 269402 106432 269404
rect 106496 269402 106502 269466
rect 106618 269402 106624 269466
rect 106688 269464 106694 269466
rect 118095 269464 118161 269467
rect 106688 269462 118161 269464
rect 106688 269406 118100 269462
rect 118156 269406 118161 269462
rect 106688 269404 118161 269406
rect 106688 269402 106694 269404
rect 118095 269401 118161 269404
rect 256335 269462 256401 269467
rect 256335 269406 256340 269462
rect 256396 269406 256401 269462
rect 256335 269401 256401 269406
rect 268143 269464 268209 269467
rect 318159 269464 318225 269467
rect 268143 269462 318225 269464
rect 268143 269406 268148 269462
rect 268204 269406 318164 269462
rect 318220 269406 318225 269462
rect 268143 269404 318225 269406
rect 268143 269401 268209 269404
rect 318159 269401 318225 269404
rect 320847 269464 320913 269467
rect 324399 269464 324465 269467
rect 320847 269462 324465 269464
rect 320847 269406 320852 269462
rect 320908 269406 324404 269462
rect 324460 269406 324465 269462
rect 320847 269404 324465 269406
rect 320847 269401 320913 269404
rect 324399 269401 324465 269404
rect 325455 269464 325521 269467
rect 328815 269464 328881 269467
rect 325455 269462 328881 269464
rect 325455 269406 325460 269462
rect 325516 269406 328820 269462
rect 328876 269406 328881 269462
rect 325455 269404 328881 269406
rect 325455 269401 325521 269404
rect 328815 269401 328881 269404
rect 329007 269464 329073 269467
rect 632079 269464 632145 269467
rect 329007 269462 632145 269464
rect 329007 269406 329012 269462
rect 329068 269406 632084 269462
rect 632140 269406 632145 269462
rect 329007 269404 632145 269406
rect 329007 269401 329073 269404
rect 632079 269401 632145 269404
rect 261615 269316 261681 269319
rect 580911 269316 580977 269319
rect 261615 269314 580977 269316
rect 261615 269258 261620 269314
rect 261676 269258 580916 269314
rect 580972 269258 580977 269314
rect 261615 269256 580977 269258
rect 261615 269253 261681 269256
rect 580911 269253 580977 269256
rect 40954 269106 40960 269170
rect 41024 269168 41030 269170
rect 41775 269168 41841 269171
rect 41024 269166 41841 269168
rect 41024 269110 41780 269166
rect 41836 269110 41841 269166
rect 41024 269108 41841 269110
rect 41024 269106 41030 269108
rect 41775 269105 41841 269108
rect 253359 269168 253425 269171
rect 513039 269168 513105 269171
rect 253359 269166 513105 269168
rect 253359 269110 253364 269166
rect 253420 269110 513044 269166
rect 513100 269110 513105 269166
rect 253359 269108 513105 269110
rect 253359 269105 253425 269108
rect 513039 269105 513105 269108
rect 674127 269168 674193 269171
rect 674127 269166 674784 269168
rect 674127 269110 674132 269166
rect 674188 269110 674784 269166
rect 674127 269108 674784 269110
rect 674127 269105 674193 269108
rect 252879 269020 252945 269023
rect 509487 269020 509553 269023
rect 252879 269018 509553 269020
rect 252879 268962 252884 269018
rect 252940 268962 509492 269018
rect 509548 268962 509553 269018
rect 252879 268960 509553 268962
rect 252879 268957 252945 268960
rect 509487 268957 509553 268960
rect 509775 269020 509841 269023
rect 524367 269020 524433 269023
rect 509775 269018 524433 269020
rect 509775 268962 509780 269018
rect 509836 268962 524372 269018
rect 524428 268962 524433 269018
rect 509775 268960 524433 268962
rect 509775 268957 509841 268960
rect 524367 268957 524433 268960
rect 252015 268872 252081 268875
rect 502287 268872 502353 268875
rect 252015 268870 502353 268872
rect 252015 268814 252020 268870
rect 252076 268814 502292 268870
rect 502348 268814 502353 268870
rect 252015 268812 502353 268814
rect 252015 268809 252081 268812
rect 502287 268809 502353 268812
rect 269199 268724 269265 268727
rect 322767 268724 322833 268727
rect 269199 268722 322833 268724
rect 269199 268666 269204 268722
rect 269260 268666 322772 268722
rect 322828 268666 322833 268722
rect 269199 268664 322833 268666
rect 269199 268661 269265 268664
rect 322767 268661 322833 268664
rect 324591 268724 324657 268727
rect 328623 268724 328689 268727
rect 324591 268722 328689 268724
rect 324591 268666 324596 268722
rect 324652 268666 328628 268722
rect 328684 268666 328689 268722
rect 324591 268664 328689 268666
rect 324591 268661 324657 268664
rect 328623 268661 328689 268664
rect 328815 268724 328881 268727
rect 577263 268724 577329 268727
rect 328815 268722 577329 268724
rect 328815 268666 328820 268722
rect 328876 268666 577268 268722
rect 577324 268666 577329 268722
rect 328815 268664 577329 268666
rect 328815 268661 328881 268664
rect 577263 268661 577329 268664
rect 258543 268576 258609 268579
rect 370575 268576 370641 268579
rect 258543 268574 370641 268576
rect 258543 268518 258548 268574
rect 258604 268518 370580 268574
rect 370636 268518 370641 268574
rect 258543 268516 370641 268518
rect 258543 268513 258609 268516
rect 370575 268513 370641 268516
rect 370767 268576 370833 268579
rect 371002 268576 371008 268578
rect 370767 268574 371008 268576
rect 370767 268518 370772 268574
rect 370828 268518 371008 268574
rect 370767 268516 371008 268518
rect 370767 268513 370833 268516
rect 371002 268514 371008 268516
rect 371072 268514 371078 268578
rect 371439 268576 371505 268579
rect 393903 268576 393969 268579
rect 371439 268574 393969 268576
rect 371439 268518 371444 268574
rect 371500 268518 393908 268574
rect 393964 268518 393969 268574
rect 371439 268516 393969 268518
rect 371439 268513 371505 268516
rect 393903 268513 393969 268516
rect 394095 268576 394161 268579
rect 398650 268576 398656 268578
rect 394095 268574 398656 268576
rect 394095 268518 394100 268574
rect 394156 268518 398656 268574
rect 394095 268516 398656 268518
rect 394095 268513 394161 268516
rect 398650 268514 398656 268516
rect 398720 268514 398726 268578
rect 398895 268576 398961 268579
rect 620079 268576 620145 268579
rect 398895 268574 620145 268576
rect 398895 268518 398900 268574
rect 398956 268518 620084 268574
rect 620140 268518 620145 268574
rect 398895 268516 620145 268518
rect 398895 268513 398961 268516
rect 620079 268513 620145 268516
rect 265071 268428 265137 268431
rect 389242 268428 389248 268430
rect 265071 268426 389248 268428
rect 265071 268370 265076 268426
rect 265132 268370 389248 268426
rect 265071 268368 389248 268370
rect 265071 268365 265137 268368
rect 389242 268366 389248 268368
rect 389312 268366 389318 268430
rect 389391 268428 389457 268431
rect 400527 268428 400593 268431
rect 389391 268426 400593 268428
rect 389391 268370 389396 268426
rect 389452 268370 400532 268426
rect 400588 268370 400593 268426
rect 389391 268368 400593 268370
rect 389391 268365 389457 268368
rect 400527 268365 400593 268368
rect 401103 268430 401169 268431
rect 401103 268426 401152 268430
rect 401216 268428 401222 268430
rect 429135 268428 429201 268431
rect 449199 268428 449265 268431
rect 401103 268370 401108 268426
rect 401103 268366 401152 268370
rect 401216 268368 401260 268428
rect 429135 268426 449265 268428
rect 429135 268370 429140 268426
rect 429196 268370 449204 268426
rect 449260 268370 449265 268426
rect 429135 268368 449265 268370
rect 401216 268366 401222 268368
rect 401103 268365 401169 268366
rect 429135 268365 429201 268368
rect 449199 268365 449265 268368
rect 260655 268280 260721 268283
rect 368367 268280 368433 268283
rect 260655 268278 368433 268280
rect 260655 268222 260660 268278
rect 260716 268222 368372 268278
rect 368428 268222 368433 268278
rect 260655 268220 368433 268222
rect 260655 268217 260721 268220
rect 368367 268217 368433 268220
rect 369231 268280 369297 268283
rect 630831 268280 630897 268283
rect 369231 268278 630897 268280
rect 369231 268222 369236 268278
rect 369292 268222 630836 268278
rect 630892 268222 630897 268278
rect 369231 268220 630897 268222
rect 369231 268217 369297 268220
rect 630831 268217 630897 268220
rect 258927 268132 258993 268135
rect 356943 268132 357009 268135
rect 368175 268132 368241 268135
rect 258927 268130 357009 268132
rect 258927 268074 258932 268130
rect 258988 268074 356948 268130
rect 357004 268074 357009 268130
rect 258927 268072 357009 268074
rect 258927 268069 258993 268072
rect 356943 268069 357009 268072
rect 357186 268130 368241 268132
rect 357186 268074 368180 268130
rect 368236 268074 368241 268130
rect 357186 268072 368241 268074
rect 258351 267984 258417 267987
rect 357186 267984 357246 268072
rect 368175 268069 368241 268072
rect 368751 268132 368817 268135
rect 389007 268132 389073 268135
rect 368751 268130 389073 268132
rect 368751 268074 368756 268130
rect 368812 268074 389012 268130
rect 389068 268074 389073 268130
rect 368751 268072 389073 268074
rect 368751 268069 368817 268072
rect 389007 268069 389073 268072
rect 389242 268070 389248 268134
rect 389312 268132 389318 268134
rect 393711 268132 393777 268135
rect 389312 268130 393777 268132
rect 389312 268074 393716 268130
rect 393772 268074 393777 268130
rect 389312 268072 393777 268074
rect 389312 268070 389318 268072
rect 393711 268069 393777 268072
rect 393903 268132 393969 268135
rect 486735 268132 486801 268135
rect 393903 268130 486801 268132
rect 393903 268074 393908 268130
rect 393964 268074 486740 268130
rect 486796 268074 486801 268130
rect 393903 268072 486801 268074
rect 393903 268069 393969 268072
rect 486735 268069 486801 268072
rect 377103 267986 377169 267987
rect 372922 267984 372928 267986
rect 258351 267982 357246 267984
rect 258351 267926 258356 267982
rect 258412 267926 357246 267982
rect 258351 267924 357246 267926
rect 357330 267924 372928 267984
rect 258351 267921 258417 267924
rect 116943 267836 117009 267839
rect 328431 267836 328497 267839
rect 116943 267834 328497 267836
rect 116943 267778 116948 267834
rect 117004 267778 328436 267834
rect 328492 267778 328497 267834
rect 116943 267776 328497 267778
rect 116943 267773 117009 267776
rect 328431 267773 328497 267776
rect 328570 267774 328576 267838
rect 328640 267836 328646 267838
rect 348783 267836 348849 267839
rect 328640 267834 348849 267836
rect 328640 267778 348788 267834
rect 348844 267778 348849 267834
rect 328640 267776 348849 267778
rect 328640 267774 328646 267776
rect 348783 267773 348849 267776
rect 348975 267836 349041 267839
rect 357330 267836 357390 267924
rect 372922 267922 372928 267924
rect 372992 267922 372998 267986
rect 377103 267982 377152 267986
rect 377216 267984 377222 267986
rect 377391 267984 377457 267987
rect 396730 267984 396736 267986
rect 377103 267926 377108 267982
rect 377103 267922 377152 267926
rect 377216 267924 377260 267984
rect 377391 267982 396736 267984
rect 377391 267926 377396 267982
rect 377452 267926 396736 267982
rect 377391 267924 396736 267926
rect 377216 267922 377222 267924
rect 377103 267921 377169 267922
rect 377391 267921 377457 267924
rect 396730 267922 396736 267924
rect 396800 267922 396806 267986
rect 396879 267984 396945 267987
rect 400378 267984 400384 267986
rect 396879 267982 400384 267984
rect 396879 267926 396884 267982
rect 396940 267926 400384 267982
rect 396879 267924 400384 267926
rect 396879 267921 396945 267924
rect 400378 267922 400384 267924
rect 400448 267922 400454 267986
rect 400527 267984 400593 267987
rect 480975 267984 481041 267987
rect 674946 267986 675006 268250
rect 400527 267982 481041 267984
rect 400527 267926 400532 267982
rect 400588 267926 480980 267982
rect 481036 267926 481041 267982
rect 400527 267924 481041 267926
rect 400527 267921 400593 267924
rect 480975 267921 481041 267924
rect 674938 267922 674944 267986
rect 675008 267922 675014 267986
rect 348975 267834 357390 267836
rect 348975 267778 348980 267834
rect 349036 267778 357390 267834
rect 348975 267776 357390 267778
rect 357807 267836 357873 267839
rect 372687 267836 372753 267839
rect 357807 267834 372753 267836
rect 357807 267778 357812 267834
rect 357868 267778 372692 267834
rect 372748 267778 372753 267834
rect 357807 267776 372753 267778
rect 348975 267773 349041 267776
rect 357807 267773 357873 267776
rect 372687 267773 372753 267776
rect 376815 267836 376881 267839
rect 389242 267836 389248 267838
rect 376815 267834 389248 267836
rect 376815 267778 376820 267834
rect 376876 267778 389248 267834
rect 376815 267776 389248 267778
rect 376815 267773 376881 267776
rect 389242 267774 389248 267776
rect 389312 267774 389318 267838
rect 391023 267836 391089 267839
rect 408591 267836 408657 267839
rect 391023 267834 408657 267836
rect 391023 267778 391028 267834
rect 391084 267778 408596 267834
rect 408652 267778 408657 267834
rect 391023 267776 408657 267778
rect 391023 267773 391089 267776
rect 408591 267773 408657 267776
rect 408783 267836 408849 267839
rect 528495 267836 528561 267839
rect 408783 267834 528561 267836
rect 408783 267778 408788 267834
rect 408844 267778 528500 267834
rect 528556 267778 528561 267834
rect 408783 267776 528561 267778
rect 408783 267773 408849 267776
rect 528495 267773 528561 267776
rect 256143 267688 256209 267691
rect 267514 267688 267520 267690
rect 256143 267686 267520 267688
rect 256143 267630 256148 267686
rect 256204 267630 267520 267686
rect 256143 267628 267520 267630
rect 256143 267625 256209 267628
rect 267514 267626 267520 267628
rect 267584 267626 267590 267690
rect 267759 267688 267825 267691
rect 530895 267688 530961 267691
rect 267759 267686 530961 267688
rect 267759 267630 267764 267686
rect 267820 267630 530900 267686
rect 530956 267630 530961 267686
rect 267759 267628 530961 267630
rect 267759 267625 267825 267628
rect 530895 267625 530961 267628
rect 188367 267540 188433 267543
rect 267855 267540 267921 267543
rect 188367 267538 267921 267540
rect 188367 267482 188372 267538
rect 188428 267482 267860 267538
rect 267916 267482 267921 267538
rect 188367 267480 267921 267482
rect 188367 267477 188433 267480
rect 267855 267477 267921 267480
rect 268047 267540 268113 267543
rect 376815 267540 376881 267543
rect 378735 267542 378801 267543
rect 268047 267538 376881 267540
rect 268047 267482 268052 267538
rect 268108 267482 376820 267538
rect 376876 267482 376881 267538
rect 268047 267480 376881 267482
rect 268047 267477 268113 267480
rect 376815 267477 376881 267480
rect 378682 267478 378688 267542
rect 378752 267540 378801 267542
rect 378752 267538 378844 267540
rect 378796 267482 378844 267538
rect 378752 267480 378844 267482
rect 378752 267478 378801 267480
rect 379066 267478 379072 267542
rect 379136 267540 379142 267542
rect 388911 267540 388977 267543
rect 379136 267538 388977 267540
rect 379136 267482 388916 267538
rect 388972 267482 388977 267538
rect 379136 267480 388977 267482
rect 379136 267478 379142 267480
rect 378735 267477 378801 267478
rect 388911 267477 388977 267480
rect 389050 267478 389056 267542
rect 389120 267540 389126 267542
rect 408687 267540 408753 267543
rect 389120 267538 408753 267540
rect 389120 267482 408692 267538
rect 408748 267482 408753 267538
rect 389120 267480 408753 267482
rect 389120 267478 389126 267480
rect 408687 267477 408753 267480
rect 408879 267540 408945 267543
rect 537999 267540 538065 267543
rect 408879 267538 538065 267540
rect 408879 267482 408884 267538
rect 408940 267482 538004 267538
rect 538060 267482 538065 267538
rect 408879 267480 538065 267482
rect 408879 267477 408945 267480
rect 537999 267477 538065 267480
rect 256335 267392 256401 267395
rect 267567 267392 267633 267395
rect 256335 267390 267633 267392
rect 256335 267334 256340 267390
rect 256396 267334 267572 267390
rect 267628 267334 267633 267390
rect 256335 267332 267633 267334
rect 256335 267329 256401 267332
rect 267567 267329 267633 267332
rect 267706 267330 267712 267394
rect 267776 267392 267782 267394
rect 396591 267392 396657 267395
rect 396783 267394 396849 267395
rect 267776 267390 396657 267392
rect 267776 267334 396596 267390
rect 396652 267334 396657 267390
rect 267776 267332 396657 267334
rect 267776 267330 267782 267332
rect 396591 267329 396657 267332
rect 396730 267330 396736 267394
rect 396800 267392 396849 267394
rect 397167 267392 397233 267395
rect 534447 267392 534513 267395
rect 396800 267390 396892 267392
rect 396844 267334 396892 267390
rect 396800 267332 396892 267334
rect 397167 267390 534513 267392
rect 397167 267334 397172 267390
rect 397228 267334 534452 267390
rect 534508 267334 534513 267390
rect 397167 267332 534513 267334
rect 396800 267330 396849 267332
rect 396783 267329 396849 267330
rect 397167 267329 397233 267332
rect 534447 267329 534513 267332
rect 256815 267244 256881 267247
rect 374127 267244 374193 267247
rect 374415 267246 374481 267247
rect 374415 267244 374464 267246
rect 256815 267242 374193 267244
rect 256815 267186 256820 267242
rect 256876 267186 374132 267242
rect 374188 267186 374193 267242
rect 256815 267184 374193 267186
rect 374372 267242 374464 267244
rect 374372 267186 374420 267242
rect 374372 267184 374464 267186
rect 256815 267181 256881 267184
rect 374127 267181 374193 267184
rect 374415 267182 374464 267184
rect 374528 267182 374534 267246
rect 374607 267244 374673 267247
rect 541551 267244 541617 267247
rect 374607 267242 541617 267244
rect 374607 267186 374612 267242
rect 374668 267186 541556 267242
rect 541612 267186 541617 267242
rect 374607 267184 541617 267186
rect 374415 267181 374481 267182
rect 374607 267181 374673 267184
rect 541551 267181 541617 267184
rect 674511 267244 674577 267247
rect 674754 267244 674814 267510
rect 674511 267242 674814 267244
rect 674511 267186 674516 267242
rect 674572 267186 674814 267242
rect 674511 267184 674814 267186
rect 674511 267181 674577 267184
rect 257199 267096 257265 267099
rect 328047 267096 328113 267099
rect 328335 267098 328401 267099
rect 328335 267096 328384 267098
rect 257199 267094 328113 267096
rect 257199 267038 257204 267094
rect 257260 267038 328052 267094
rect 328108 267038 328113 267094
rect 257199 267036 328113 267038
rect 328292 267094 328384 267096
rect 328292 267038 328340 267094
rect 328292 267036 328384 267038
rect 257199 267033 257265 267036
rect 328047 267033 328113 267036
rect 328335 267034 328384 267036
rect 328448 267034 328454 267098
rect 328570 267034 328576 267098
rect 328640 267096 328646 267098
rect 349359 267096 349425 267099
rect 368506 267096 368512 267098
rect 328640 267036 348222 267096
rect 328640 267034 328646 267036
rect 328335 267033 328401 267034
rect 72975 266948 73041 266951
rect 328431 266948 328497 266951
rect 72975 266946 328497 266948
rect 72975 266890 72980 266946
rect 73036 266890 328436 266946
rect 328492 266890 328497 266946
rect 72975 266888 328497 266890
rect 72975 266885 73041 266888
rect 328431 266885 328497 266888
rect 328623 266948 328689 266951
rect 347823 266948 347889 266951
rect 328623 266946 347889 266948
rect 328623 266890 328628 266946
rect 328684 266890 347828 266946
rect 347884 266890 347889 266946
rect 328623 266888 347889 266890
rect 348162 266948 348222 267036
rect 349359 267094 368512 267096
rect 349359 267038 349364 267094
rect 349420 267038 368512 267094
rect 349359 267036 368512 267038
rect 349359 267033 349425 267036
rect 368506 267034 368512 267036
rect 368576 267034 368582 267098
rect 368751 267096 368817 267099
rect 388090 267096 388096 267098
rect 368751 267094 388096 267096
rect 368751 267038 368756 267094
rect 368812 267038 388096 267094
rect 368751 267036 388096 267038
rect 368751 267033 368817 267036
rect 388090 267034 388096 267036
rect 388160 267034 388166 267098
rect 388282 267034 388288 267098
rect 388352 267096 388358 267098
rect 545199 267096 545265 267099
rect 388352 267094 545265 267096
rect 388352 267038 545204 267094
rect 545260 267038 545265 267094
rect 388352 267036 545265 267038
rect 388352 267034 388358 267036
rect 545199 267033 545265 267036
rect 348495 266948 348561 266951
rect 348162 266946 348561 266948
rect 348162 266890 348500 266946
rect 348556 266890 348561 266946
rect 348162 266888 348561 266890
rect 328623 266885 328689 266888
rect 347823 266885 347889 266888
rect 348495 266885 348561 266888
rect 348783 266948 348849 266951
rect 368463 266948 368529 266951
rect 348783 266946 368529 266948
rect 348783 266890 348788 266946
rect 348844 266890 368468 266946
rect 368524 266890 368529 266946
rect 348783 266888 368529 266890
rect 348783 266885 348849 266888
rect 368463 266885 368529 266888
rect 368655 266948 368721 266951
rect 388815 266948 388881 266951
rect 368655 266946 388881 266948
rect 368655 266890 368660 266946
rect 368716 266890 388820 266946
rect 388876 266890 388881 266946
rect 368655 266888 388881 266890
rect 368655 266885 368721 266888
rect 388815 266885 388881 266888
rect 389434 266886 389440 266950
rect 389504 266948 389510 266950
rect 408495 266948 408561 266951
rect 389504 266946 408561 266948
rect 389504 266890 408500 266946
rect 408556 266890 408561 266946
rect 389504 266888 408561 266890
rect 389504 266886 389510 266888
rect 408495 266885 408561 266888
rect 408783 266948 408849 266951
rect 419151 266948 419217 266951
rect 408783 266946 419217 266948
rect 408783 266890 408788 266946
rect 408844 266890 419156 266946
rect 419212 266890 419217 266946
rect 408783 266888 419217 266890
rect 408783 266885 408849 266888
rect 419151 266885 419217 266888
rect 419343 266948 419409 266951
rect 542799 266948 542865 266951
rect 419343 266946 542865 266948
rect 419343 266890 419348 266946
rect 419404 266890 542804 266946
rect 542860 266890 542865 266946
rect 419343 266888 542865 266890
rect 419343 266885 419409 266888
rect 542799 266885 542865 266888
rect 132495 266800 132561 266803
rect 287631 266800 287697 266803
rect 132495 266798 287697 266800
rect 132495 266742 132500 266798
rect 132556 266742 287636 266798
rect 287692 266742 287697 266798
rect 132495 266740 287697 266742
rect 132495 266737 132561 266740
rect 287631 266737 287697 266740
rect 287919 266800 287985 266803
rect 328378 266800 328384 266802
rect 287919 266798 328384 266800
rect 287919 266742 287924 266798
rect 287980 266742 328384 266798
rect 287919 266740 328384 266742
rect 287919 266737 287985 266740
rect 328378 266738 328384 266740
rect 328448 266738 328454 266802
rect 328762 266738 328768 266802
rect 328832 266800 328838 266802
rect 348687 266800 348753 266803
rect 389050 266800 389056 266802
rect 328832 266740 348030 266800
rect 328832 266738 328838 266740
rect 206991 266652 207057 266655
rect 287631 266652 287697 266655
rect 206991 266650 287697 266652
rect 206991 266594 206996 266650
rect 207052 266594 287636 266650
rect 287692 266594 287697 266650
rect 206991 266592 287697 266594
rect 206991 266589 207057 266592
rect 287631 266589 287697 266592
rect 287919 266652 287985 266655
rect 328527 266652 328593 266655
rect 287919 266650 328593 266652
rect 287919 266594 287924 266650
rect 287980 266594 328532 266650
rect 328588 266594 328593 266650
rect 287919 266592 328593 266594
rect 287919 266589 287985 266592
rect 328527 266589 328593 266592
rect 329295 266652 329361 266655
rect 347727 266652 347793 266655
rect 329295 266650 347793 266652
rect 329295 266594 329300 266650
rect 329356 266594 347732 266650
rect 347788 266594 347793 266650
rect 329295 266592 347793 266594
rect 347970 266652 348030 266740
rect 348687 266798 389056 266800
rect 348687 266742 348692 266798
rect 348748 266742 389056 266798
rect 348687 266740 389056 266742
rect 348687 266737 348753 266740
rect 389050 266738 389056 266740
rect 389120 266738 389126 266802
rect 389626 266738 389632 266802
rect 389696 266800 389702 266802
rect 439119 266800 439185 266803
rect 389696 266798 439185 266800
rect 389696 266742 439124 266798
rect 439180 266742 439185 266798
rect 389696 266740 439185 266742
rect 389696 266738 389702 266740
rect 439119 266737 439185 266740
rect 459279 266800 459345 266803
rect 479343 266800 479409 266803
rect 459279 266798 479409 266800
rect 459279 266742 459284 266798
rect 459340 266742 479348 266798
rect 479404 266742 479409 266798
rect 459279 266740 479409 266742
rect 459279 266737 459345 266740
rect 479343 266737 479409 266740
rect 479535 266800 479601 266803
rect 642735 266800 642801 266803
rect 479535 266798 642801 266800
rect 479535 266742 479540 266798
rect 479596 266742 642740 266798
rect 642796 266742 642801 266798
rect 479535 266740 642801 266742
rect 479535 266737 479601 266740
rect 642735 266737 642801 266740
rect 349071 266652 349137 266655
rect 347970 266650 349137 266652
rect 347970 266594 349076 266650
rect 349132 266594 349137 266650
rect 347970 266592 349137 266594
rect 329295 266589 329361 266592
rect 347727 266589 347793 266592
rect 349071 266589 349137 266592
rect 349839 266652 349905 266655
rect 368367 266652 368433 266655
rect 349839 266650 368433 266652
rect 349839 266594 349844 266650
rect 349900 266594 368372 266650
rect 368428 266594 368433 266650
rect 349839 266592 368433 266594
rect 349839 266589 349905 266592
rect 368367 266589 368433 266592
rect 368506 266590 368512 266654
rect 368576 266652 368582 266654
rect 388623 266652 388689 266655
rect 368576 266650 388689 266652
rect 368576 266594 388628 266650
rect 388684 266594 388689 266650
rect 368576 266592 388689 266594
rect 368576 266590 368582 266592
rect 388623 266589 388689 266592
rect 389434 266590 389440 266654
rect 389504 266652 389510 266654
rect 399279 266652 399345 266655
rect 389504 266650 399345 266652
rect 389504 266594 399284 266650
rect 399340 266594 399345 266650
rect 389504 266592 399345 266594
rect 389504 266590 389510 266592
rect 399279 266589 399345 266592
rect 399471 266652 399537 266655
rect 400143 266654 400209 266655
rect 399994 266652 400000 266654
rect 399471 266650 400000 266652
rect 399471 266594 399476 266650
rect 399532 266594 400000 266650
rect 399471 266592 400000 266594
rect 399471 266589 399537 266592
rect 399994 266590 400000 266592
rect 400064 266590 400070 266654
rect 400143 266650 400192 266654
rect 400256 266652 400262 266654
rect 400431 266652 400497 266655
rect 400570 266652 400576 266654
rect 400143 266594 400148 266650
rect 400143 266590 400192 266594
rect 400256 266592 400300 266652
rect 400431 266650 400576 266652
rect 400431 266594 400436 266650
rect 400492 266594 400576 266650
rect 400431 266592 400576 266594
rect 400256 266590 400262 266592
rect 400143 266589 400209 266590
rect 400431 266589 400497 266592
rect 400570 266590 400576 266592
rect 400640 266590 400646 266654
rect 401199 266652 401265 266655
rect 401338 266652 401344 266654
rect 401199 266650 401344 266652
rect 401199 266594 401204 266650
rect 401260 266594 401344 266650
rect 401199 266592 401344 266594
rect 401199 266589 401265 266592
rect 401338 266590 401344 266592
rect 401408 266590 401414 266654
rect 401530 266590 401536 266654
rect 401600 266652 401606 266654
rect 402447 266652 402513 266655
rect 401600 266650 402513 266652
rect 401600 266594 402452 266650
rect 402508 266594 402513 266650
rect 401600 266592 402513 266594
rect 401600 266590 401606 266592
rect 402447 266589 402513 266592
rect 403215 266654 403281 266655
rect 403215 266650 403264 266654
rect 403328 266652 403334 266654
rect 403887 266652 403953 266655
rect 404751 266654 404817 266655
rect 405231 266654 405297 266655
rect 406191 266654 406257 266655
rect 406575 266654 406641 266655
rect 404602 266652 404608 266654
rect 403215 266594 403220 266650
rect 403215 266590 403264 266594
rect 403328 266592 403372 266652
rect 403887 266650 404608 266652
rect 403887 266594 403892 266650
rect 403948 266594 404608 266650
rect 403887 266592 404608 266594
rect 403328 266590 403334 266592
rect 403215 266589 403281 266590
rect 403887 266589 403953 266592
rect 404602 266590 404608 266592
rect 404672 266590 404678 266654
rect 404751 266650 404800 266654
rect 404864 266652 404870 266654
rect 405178 266652 405184 266654
rect 404751 266594 404756 266650
rect 404751 266590 404800 266594
rect 404864 266592 404908 266652
rect 405140 266592 405184 266652
rect 405248 266650 405297 266654
rect 406138 266652 406144 266654
rect 405292 266594 405297 266650
rect 404864 266590 404870 266592
rect 405178 266590 405184 266592
rect 405248 266590 405297 266594
rect 406100 266592 406144 266652
rect 406208 266650 406257 266654
rect 406522 266652 406528 266654
rect 406252 266594 406257 266650
rect 406138 266590 406144 266592
rect 406208 266590 406257 266594
rect 406484 266592 406528 266652
rect 406592 266650 406641 266654
rect 406863 266654 406929 266655
rect 407151 266654 407217 266655
rect 406863 266652 406912 266654
rect 406636 266594 406641 266650
rect 406522 266590 406528 266592
rect 406592 266590 406641 266594
rect 406820 266650 406912 266652
rect 406820 266594 406868 266650
rect 406820 266592 406912 266594
rect 404751 266589 404817 266590
rect 405231 266589 405297 266590
rect 406191 266589 406257 266590
rect 406575 266589 406641 266590
rect 406863 266590 406912 266592
rect 406976 266590 406982 266654
rect 407098 266652 407104 266654
rect 407060 266592 407104 266652
rect 407168 266650 407217 266654
rect 407212 266594 407217 266650
rect 407098 266590 407104 266592
rect 407168 266590 407217 266594
rect 406863 266589 406929 266590
rect 407151 266589 407217 266590
rect 407343 266652 407409 266655
rect 408783 266652 408849 266655
rect 409071 266654 409137 266655
rect 409455 266654 409521 266655
rect 409018 266652 409024 266654
rect 407343 266650 408849 266652
rect 407343 266594 407348 266650
rect 407404 266594 408788 266650
rect 408844 266594 408849 266650
rect 407343 266592 408849 266594
rect 408980 266592 409024 266652
rect 409088 266650 409137 266654
rect 409402 266652 409408 266654
rect 409132 266594 409137 266650
rect 407343 266589 407409 266592
rect 408783 266589 408849 266592
rect 409018 266590 409024 266592
rect 409088 266590 409137 266594
rect 409364 266592 409408 266652
rect 409472 266650 409521 266654
rect 409516 266594 409521 266650
rect 409402 266590 409408 266592
rect 409472 266590 409521 266594
rect 409071 266589 409137 266590
rect 409455 266589 409521 266590
rect 409647 266652 409713 266655
rect 419151 266652 419217 266655
rect 439215 266652 439281 266655
rect 409647 266650 419070 266652
rect 409647 266594 409652 266650
rect 409708 266594 419070 266650
rect 409647 266592 419070 266594
rect 409647 266589 409713 266592
rect 419010 266504 419070 266592
rect 419151 266650 439281 266652
rect 419151 266594 419156 266650
rect 419212 266594 439220 266650
rect 439276 266594 439281 266650
rect 419151 266592 439281 266594
rect 419151 266589 419217 266592
rect 439215 266589 439281 266592
rect 459375 266652 459441 266655
rect 479439 266652 479505 266655
rect 459375 266650 479505 266652
rect 459375 266594 459380 266650
rect 459436 266594 479444 266650
rect 479500 266594 479505 266650
rect 459375 266592 479505 266594
rect 459375 266589 459441 266592
rect 479439 266589 479505 266592
rect 479631 266652 479697 266655
rect 646287 266652 646353 266655
rect 479631 266650 646353 266652
rect 479631 266594 479636 266650
rect 479692 266594 646292 266650
rect 646348 266594 646353 266650
rect 479631 266592 646353 266594
rect 479631 266589 479697 266592
rect 646287 266589 646353 266592
rect 673935 266652 674001 266655
rect 673935 266650 674784 266652
rect 673935 266594 673940 266650
rect 673996 266594 674784 266650
rect 673935 266592 674784 266594
rect 673935 266589 674001 266592
rect 505263 266504 505329 266507
rect 419010 266502 505329 266504
rect 419010 266446 505268 266502
rect 505324 266446 505329 266502
rect 419010 266444 505329 266446
rect 505263 266441 505329 266444
rect 413775 266356 413841 266359
rect 419343 266356 419409 266359
rect 439023 266356 439089 266359
rect 413775 266354 419409 266356
rect 413775 266298 413780 266354
rect 413836 266298 419348 266354
rect 419404 266298 419409 266354
rect 413775 266296 419409 266298
rect 413775 266293 413841 266296
rect 419343 266293 419409 266296
rect 419586 266354 439089 266356
rect 419586 266298 439028 266354
rect 439084 266298 439089 266354
rect 419586 266296 439089 266298
rect 413679 266208 413745 266211
rect 419586 266208 419646 266296
rect 439023 266293 439089 266296
rect 458127 266356 458193 266359
rect 479535 266356 479601 266359
rect 458127 266354 479601 266356
rect 458127 266298 458132 266354
rect 458188 266298 479540 266354
rect 479596 266298 479601 266354
rect 458127 266296 479601 266298
rect 458127 266293 458193 266296
rect 479535 266293 479601 266296
rect 439311 266208 439377 266211
rect 413679 266206 419646 266208
rect 413679 266150 413684 266206
rect 413740 266150 419646 266206
rect 413679 266148 419646 266150
rect 419778 266206 439377 266208
rect 419778 266150 439316 266206
rect 439372 266150 439377 266206
rect 419778 266148 439377 266150
rect 413679 266145 413745 266148
rect 413391 265912 413457 265915
rect 419778 265912 419838 266148
rect 439311 266145 439377 266148
rect 479439 266208 479505 266211
rect 501231 266208 501297 266211
rect 479439 266206 501297 266208
rect 479439 266150 479444 266206
rect 479500 266150 501236 266206
rect 501292 266150 501297 266206
rect 479439 266148 501297 266150
rect 479439 266145 479505 266148
rect 501231 266145 501297 266148
rect 439119 266060 439185 266063
rect 459279 266060 459345 266063
rect 439119 266058 459345 266060
rect 439119 266002 439124 266058
rect 439180 266002 459284 266058
rect 459340 266002 459345 266058
rect 439119 266000 459345 266002
rect 439119 265997 439185 266000
rect 459279 265997 459345 266000
rect 479343 266060 479409 266063
rect 479343 266058 479934 266060
rect 479343 266002 479348 266058
rect 479404 266002 479934 266058
rect 479343 266000 479934 266002
rect 479343 265997 479409 266000
rect 413391 265910 419838 265912
rect 413391 265854 413396 265910
rect 413452 265854 419838 265910
rect 413391 265852 419838 265854
rect 439215 265912 439281 265915
rect 459375 265912 459441 265915
rect 439215 265910 459441 265912
rect 439215 265854 439220 265910
rect 439276 265854 459380 265910
rect 459436 265854 459441 265910
rect 439215 265852 459441 265854
rect 413391 265849 413457 265852
rect 439215 265849 439281 265852
rect 459375 265849 459441 265852
rect 459567 265912 459633 265915
rect 479631 265912 479697 265915
rect 459567 265910 479697 265912
rect 459567 265854 459572 265910
rect 459628 265854 479636 265910
rect 479692 265854 479697 265910
rect 459567 265852 479697 265854
rect 479874 265912 479934 266000
rect 497679 265912 497745 265915
rect 479874 265910 497745 265912
rect 479874 265854 497684 265910
rect 497740 265854 497745 265910
rect 479874 265852 497745 265854
rect 459567 265849 459633 265852
rect 479631 265849 479697 265852
rect 497679 265849 497745 265852
rect 413199 265764 413265 265767
rect 635535 265764 635601 265767
rect 413199 265762 635601 265764
rect 413199 265706 413204 265762
rect 413260 265706 635540 265762
rect 635596 265706 635601 265762
rect 413199 265704 635601 265706
rect 413199 265701 413265 265704
rect 635535 265701 635601 265704
rect 439023 265616 439089 265619
rect 458127 265616 458193 265619
rect 439023 265614 458193 265616
rect 439023 265558 439028 265614
rect 439084 265558 458132 265614
rect 458188 265558 458193 265614
rect 439023 265556 458193 265558
rect 439023 265553 439089 265556
rect 458127 265553 458193 265556
rect 439311 265468 439377 265471
rect 459567 265468 459633 265471
rect 439311 265466 459633 265468
rect 439311 265410 439316 265466
rect 439372 265410 459572 265466
rect 459628 265410 459633 265466
rect 439311 265408 459633 265410
rect 439311 265405 439377 265408
rect 459567 265405 459633 265408
rect 674554 265406 674560 265470
rect 674624 265468 674630 265470
rect 674754 265468 674814 266030
rect 674624 265408 674814 265468
rect 674624 265406 674630 265408
rect 413199 265320 413265 265323
rect 455055 265320 455121 265323
rect 413199 265318 455121 265320
rect 413199 265262 413204 265318
rect 413260 265262 455060 265318
rect 455116 265262 455121 265318
rect 413199 265260 455121 265262
rect 413199 265257 413265 265260
rect 455055 265257 455121 265260
rect 475119 265172 475185 265175
rect 483855 265172 483921 265175
rect 475119 265170 483921 265172
rect 475119 265114 475124 265170
rect 475180 265114 483860 265170
rect 483916 265114 483921 265170
rect 475119 265112 483921 265114
rect 475119 265109 475185 265112
rect 483855 265109 483921 265112
rect 511119 265172 511185 265175
rect 607023 265172 607089 265175
rect 511119 265170 523518 265172
rect 511119 265114 511124 265170
rect 511180 265114 523518 265170
rect 511119 265112 523518 265114
rect 511119 265109 511185 265112
rect 412527 265024 412593 265027
rect 521391 265024 521457 265027
rect 412527 265022 521457 265024
rect 325455 264989 325521 264990
rect 365007 264989 365073 264990
rect 325455 264987 325504 264989
rect 325412 264985 325504 264987
rect 325412 264929 325460 264985
rect 325412 264927 325504 264929
rect 325455 264925 325504 264927
rect 325568 264925 325574 264989
rect 365007 264987 365056 264989
rect 364964 264985 365056 264987
rect 364964 264929 365012 264985
rect 364964 264927 365056 264929
rect 365007 264925 365056 264927
rect 365120 264925 365126 264989
rect 400762 264925 400768 264989
rect 400832 264987 400838 264989
rect 401583 264987 401649 264990
rect 400832 264985 401649 264987
rect 400832 264929 401588 264985
rect 401644 264929 401649 264985
rect 412527 264966 412532 265022
rect 412588 264966 521396 265022
rect 521452 264966 521457 265022
rect 412527 264964 521457 264966
rect 523458 265024 523518 265112
rect 537474 265112 563262 265172
rect 537474 265024 537534 265112
rect 523458 264964 537534 265024
rect 563202 265024 563262 265112
rect 594690 265170 607089 265172
rect 594690 265114 607028 265170
rect 607084 265114 607089 265170
rect 594690 265112 607089 265114
rect 594690 265024 594750 265112
rect 607023 265109 607089 265112
rect 678210 265027 678270 265142
rect 563202 264964 594750 265024
rect 678159 265022 678270 265027
rect 678159 264966 678164 265022
rect 678220 264966 678270 265022
rect 678159 264964 678270 264966
rect 412527 264961 412593 264964
rect 521391 264961 521457 264964
rect 678159 264961 678225 264964
rect 400832 264927 401649 264929
rect 400832 264925 400838 264927
rect 325455 264924 325521 264925
rect 365007 264924 365073 264925
rect 401583 264924 401649 264927
rect 42255 264284 42321 264287
rect 42255 264282 42366 264284
rect 42255 264226 42260 264282
rect 42316 264226 42366 264282
rect 42255 264221 42366 264226
rect 42306 264106 42366 264221
rect 674607 264136 674673 264139
rect 674754 264136 674814 264402
rect 674607 264134 674814 264136
rect 674607 264078 674612 264134
rect 674668 264078 674814 264134
rect 674607 264076 674814 264078
rect 674607 264073 674673 264076
rect 674031 263544 674097 263547
rect 674031 263542 674784 263544
rect 674031 263486 674036 263542
rect 674092 263486 674784 263542
rect 674031 263484 674784 263486
rect 674031 263481 674097 263484
rect 42639 263248 42705 263251
rect 42336 263246 42705 263248
rect 42336 263190 42644 263246
rect 42700 263190 42705 263246
rect 42336 263188 42705 263190
rect 42639 263185 42705 263188
rect 674319 262804 674385 262807
rect 674319 262802 674784 262804
rect 674319 262746 674324 262802
rect 674380 262746 674784 262802
rect 674319 262744 674784 262746
rect 674319 262741 674385 262744
rect 42639 262508 42705 262511
rect 42336 262506 42705 262508
rect 42336 262450 42644 262506
rect 42700 262450 42705 262506
rect 42336 262448 42705 262450
rect 42639 262445 42705 262448
rect 211503 261906 211569 261909
rect 211503 261904 211872 261906
rect 211503 261848 211508 261904
rect 211564 261848 211872 261904
rect 211503 261846 211872 261848
rect 211503 261843 211569 261846
rect 676866 261771 676926 261886
rect 676866 261766 676977 261771
rect 676866 261710 676916 261766
rect 676972 261710 676977 261766
rect 676866 261708 676977 261710
rect 676911 261705 676977 261708
rect 43503 261620 43569 261623
rect 42336 261618 43569 261620
rect 42336 261562 43508 261618
rect 43564 261562 43569 261618
rect 42336 261560 43569 261562
rect 43503 261557 43569 261560
rect 676866 261031 676926 261220
rect 676815 261026 676926 261031
rect 676815 260970 676820 261026
rect 676876 260970 676926 261026
rect 676815 260968 676926 260970
rect 676815 260965 676881 260968
rect 43215 260880 43281 260883
rect 42336 260878 43281 260880
rect 42336 260822 43220 260878
rect 43276 260822 43281 260878
rect 42336 260820 43281 260822
rect 43215 260817 43281 260820
rect 42490 260436 42496 260438
rect 42306 260376 42496 260436
rect 42306 260140 42366 260376
rect 42490 260374 42496 260376
rect 42560 260374 42566 260438
rect 675330 260143 675390 260406
rect 41376 260110 42366 260140
rect 675279 260138 675390 260143
rect 41346 260080 42336 260110
rect 675279 260082 675284 260138
rect 675340 260082 675390 260138
rect 675279 260080 675390 260082
rect 41346 259551 41406 260080
rect 675279 260077 675345 260080
rect 41295 259546 41406 259551
rect 41295 259490 41300 259546
rect 41356 259490 41406 259546
rect 41295 259488 41406 259490
rect 41295 259485 41361 259488
rect 42106 259486 42112 259550
rect 42176 259486 42182 259550
rect 42114 259400 42174 259486
rect 675138 259403 675198 259592
rect 43407 259400 43473 259403
rect 42114 259398 43473 259400
rect 42114 259370 43412 259398
rect 42144 259342 43412 259370
rect 43468 259342 43473 259398
rect 42144 259340 43473 259342
rect 675138 259398 675249 259403
rect 675138 259342 675188 259398
rect 675244 259342 675249 259398
rect 675138 259340 675249 259342
rect 43407 259337 43473 259340
rect 675183 259337 675249 259340
rect 674223 258808 674289 258811
rect 674223 258806 674784 258808
rect 674223 258750 674228 258806
rect 674284 258750 674784 258806
rect 674223 258748 674784 258750
rect 674223 258745 674289 258748
rect 41538 257922 41598 258482
rect 41530 257858 41536 257922
rect 41600 257858 41606 257922
rect 42114 257183 42174 257742
rect 679746 257479 679806 257964
rect 679746 257474 679857 257479
rect 679746 257418 679796 257474
rect 679852 257418 679857 257474
rect 679746 257416 679857 257418
rect 679791 257413 679857 257416
rect 42063 257178 42174 257183
rect 42063 257122 42068 257178
rect 42124 257122 42174 257178
rect 42063 257120 42174 257122
rect 42063 257117 42129 257120
rect 679791 256884 679857 256887
rect 679746 256882 679857 256884
rect 40386 256294 40446 256854
rect 679746 256826 679796 256882
rect 679852 256826 679857 256882
rect 679746 256821 679857 256826
rect 679746 256410 679806 256821
rect 40378 256230 40384 256294
rect 40448 256230 40454 256294
rect 40962 255702 41022 256114
rect 40954 255638 40960 255702
rect 41024 255638 41030 255702
rect 207279 255404 207345 255407
rect 211842 255404 211902 255864
rect 207279 255402 211902 255404
rect 41154 254814 41214 255374
rect 207279 255346 207284 255402
rect 207340 255346 211902 255402
rect 207279 255344 211902 255346
rect 207279 255341 207345 255344
rect 41146 254750 41152 254814
rect 41216 254750 41222 254814
rect 41730 254371 41790 254560
rect 41730 254366 41841 254371
rect 41730 254310 41780 254366
rect 41836 254310 41841 254366
rect 41730 254308 41841 254310
rect 41775 254305 41841 254308
rect 40770 253482 40830 253746
rect 40762 253418 40768 253482
rect 40832 253418 40838 253482
rect 675706 253418 675712 253482
rect 675776 253480 675782 253482
rect 678159 253480 678225 253483
rect 675776 253478 678225 253480
rect 675776 253422 678164 253478
rect 678220 253422 678225 253478
rect 675776 253420 678225 253422
rect 675776 253418 675782 253420
rect 678159 253417 678225 253420
rect 41346 252742 41406 252932
rect 41338 252678 41344 252742
rect 41408 252678 41414 252742
rect 40194 251559 40254 252118
rect 40194 251554 40305 251559
rect 40194 251498 40244 251554
rect 40300 251498 40305 251554
rect 40194 251496 40305 251498
rect 40239 251493 40305 251496
rect 37314 250819 37374 251304
rect 37314 250814 37425 250819
rect 40047 250816 40113 250819
rect 37314 250758 37364 250814
rect 37420 250758 37425 250814
rect 37314 250756 37425 250758
rect 37359 250753 37425 250756
rect 40002 250814 40113 250816
rect 40002 250758 40052 250814
rect 40108 250758 40113 250814
rect 40002 250753 40113 250758
rect 40002 250638 40062 250753
rect 206895 249928 206961 249931
rect 206895 249926 211872 249928
rect 206895 249870 206900 249926
rect 206956 249870 211872 249926
rect 206895 249868 211872 249870
rect 206895 249865 206961 249868
rect 42306 249188 42366 249750
rect 42543 249188 42609 249191
rect 42306 249186 42609 249188
rect 42306 249130 42548 249186
rect 42604 249130 42609 249186
rect 42306 249128 42609 249130
rect 42543 249125 42609 249128
rect 40194 248451 40254 249010
rect 40143 248446 40254 248451
rect 40143 248390 40148 248446
rect 40204 248390 40254 248446
rect 40143 248388 40254 248390
rect 40143 248385 40209 248388
rect 42306 247560 42366 248122
rect 143919 247708 143985 247711
rect 156879 247708 156945 247711
rect 143919 247706 156945 247708
rect 143919 247650 143924 247706
rect 143980 247650 156884 247706
rect 156940 247650 156945 247706
rect 143919 247648 156945 247650
rect 143919 247645 143985 247648
rect 156879 247645 156945 247648
rect 161103 247708 161169 247711
rect 161103 247706 197310 247708
rect 161103 247650 161108 247706
rect 161164 247650 197310 247706
rect 161103 247648 197310 247650
rect 161103 247645 161169 247648
rect 43023 247560 43089 247563
rect 42306 247558 43089 247560
rect 42306 247502 43028 247558
rect 43084 247502 43089 247558
rect 42306 247500 43089 247502
rect 43023 247497 43089 247500
rect 140943 247560 141009 247563
rect 197250 247560 197310 247648
rect 404794 247560 404800 247562
rect 140943 247558 187902 247560
rect 140943 247502 140948 247558
rect 141004 247502 187902 247558
rect 140943 247500 187902 247502
rect 197250 247500 404800 247560
rect 140943 247497 141009 247500
rect 146703 247412 146769 247415
rect 187842 247412 187902 247500
rect 404794 247498 404800 247500
rect 404864 247498 404870 247562
rect 406330 247412 406336 247414
rect 146703 247410 187710 247412
rect 42159 247118 42225 247119
rect 42106 247116 42112 247118
rect 42068 247056 42112 247116
rect 42176 247114 42225 247118
rect 42220 247058 42225 247114
rect 42106 247054 42112 247056
rect 42176 247054 42225 247058
rect 42159 247053 42225 247054
rect 42306 246823 42366 247382
rect 146703 247354 146708 247410
rect 146764 247354 187710 247410
rect 146703 247352 187710 247354
rect 187842 247352 369150 247412
rect 146703 247349 146769 247352
rect 156879 247264 156945 247267
rect 171663 247264 171729 247267
rect 156879 247262 171729 247264
rect 156879 247206 156884 247262
rect 156940 247206 171668 247262
rect 171724 247206 171729 247262
rect 156879 247204 171729 247206
rect 187650 247264 187710 247352
rect 188175 247264 188241 247267
rect 187650 247204 188094 247264
rect 156879 247201 156945 247204
rect 171663 247201 171729 247204
rect 149583 247116 149649 247119
rect 187887 247116 187953 247119
rect 149583 247114 187953 247116
rect 149583 247058 149588 247114
rect 149644 247058 187892 247114
rect 187948 247058 187953 247114
rect 149583 247056 187953 247058
rect 188034 247116 188094 247204
rect 188175 247262 368574 247264
rect 188175 247206 188180 247262
rect 188236 247206 368574 247262
rect 188175 247204 368574 247206
rect 188175 247201 188241 247204
rect 188034 247056 368190 247116
rect 149583 247053 149649 247056
rect 187887 247053 187953 247056
rect 155343 246968 155409 246971
rect 187695 246968 187761 246971
rect 155343 246966 187761 246968
rect 155343 246910 155348 246966
rect 155404 246910 187700 246966
rect 187756 246910 187761 246966
rect 155343 246908 187761 246910
rect 155343 246905 155409 246908
rect 187695 246905 187761 246908
rect 201519 246968 201585 246971
rect 201519 246966 367806 246968
rect 201519 246910 201524 246966
rect 201580 246910 367806 246966
rect 201519 246908 367806 246910
rect 201519 246905 201585 246908
rect 42306 246818 42417 246823
rect 42306 246762 42356 246818
rect 42412 246762 42417 246818
rect 42306 246760 42417 246762
rect 42351 246757 42417 246760
rect 42874 246758 42880 246822
rect 42944 246820 42950 246822
rect 187599 246820 187665 246823
rect 216879 246820 216945 246823
rect 42944 246818 187665 246820
rect 42944 246762 187604 246818
rect 187660 246762 187665 246818
rect 42944 246760 187665 246762
rect 42944 246758 42950 246760
rect 187599 246757 187665 246760
rect 187842 246818 216945 246820
rect 187842 246762 216884 246818
rect 216940 246762 216945 246818
rect 187842 246760 216945 246762
rect 90639 246672 90705 246675
rect 100527 246672 100593 246675
rect 90639 246670 100593 246672
rect 90639 246614 90644 246670
rect 90700 246614 100532 246670
rect 100588 246614 100593 246670
rect 90639 246612 100593 246614
rect 90639 246609 90705 246612
rect 100527 246609 100593 246612
rect 177039 246672 177105 246675
rect 187842 246672 187902 246760
rect 216879 246757 216945 246760
rect 227919 246820 227985 246823
rect 246447 246820 246513 246823
rect 227919 246818 246513 246820
rect 227919 246762 227924 246818
rect 227980 246762 246452 246818
rect 246508 246762 246513 246818
rect 227919 246760 246513 246762
rect 227919 246757 227985 246760
rect 246447 246757 246513 246760
rect 247546 246758 247552 246822
rect 247616 246820 247622 246822
rect 247791 246820 247857 246823
rect 247616 246818 247857 246820
rect 247616 246762 247796 246818
rect 247852 246762 247857 246818
rect 247616 246760 247857 246762
rect 247616 246758 247622 246760
rect 247791 246757 247857 246760
rect 248367 246820 248433 246823
rect 259215 246820 259281 246823
rect 248367 246818 259281 246820
rect 248367 246762 248372 246818
rect 248428 246762 259220 246818
rect 259276 246762 259281 246818
rect 248367 246760 259281 246762
rect 248367 246757 248433 246760
rect 259215 246757 259281 246760
rect 267951 246820 268017 246823
rect 291951 246820 292017 246823
rect 267951 246818 292017 246820
rect 267951 246762 267956 246818
rect 268012 246762 291956 246818
rect 292012 246762 292017 246818
rect 267951 246760 292017 246762
rect 267951 246757 268017 246760
rect 291951 246757 292017 246760
rect 292143 246820 292209 246823
rect 307983 246820 308049 246823
rect 292143 246818 308049 246820
rect 292143 246762 292148 246818
rect 292204 246762 307988 246818
rect 308044 246762 308049 246818
rect 292143 246760 308049 246762
rect 292143 246757 292209 246760
rect 307983 246757 308049 246760
rect 311151 246820 311217 246823
rect 327087 246820 327153 246823
rect 311151 246818 327153 246820
rect 311151 246762 311156 246818
rect 311212 246762 327092 246818
rect 327148 246762 327153 246818
rect 311151 246760 327153 246762
rect 311151 246757 311217 246760
rect 327087 246757 327153 246760
rect 327951 246820 328017 246823
rect 328335 246820 328401 246823
rect 327951 246818 328401 246820
rect 327951 246762 327956 246818
rect 328012 246762 328340 246818
rect 328396 246762 328401 246818
rect 327951 246760 328401 246762
rect 327951 246757 328017 246760
rect 328335 246757 328401 246760
rect 328527 246820 328593 246823
rect 348111 246820 348177 246823
rect 328527 246818 348177 246820
rect 328527 246762 328532 246818
rect 328588 246762 348116 246818
rect 348172 246762 348177 246818
rect 328527 246760 348177 246762
rect 328527 246757 328593 246760
rect 348111 246757 348177 246760
rect 348591 246820 348657 246823
rect 360058 246820 360064 246822
rect 348591 246818 360064 246820
rect 348591 246762 348596 246818
rect 348652 246762 360064 246818
rect 348591 246760 360064 246762
rect 348591 246757 348657 246760
rect 360058 246758 360064 246760
rect 360128 246758 360134 246822
rect 360442 246758 360448 246822
rect 360512 246820 360518 246822
rect 367599 246820 367665 246823
rect 367746 246822 367806 246908
rect 360512 246818 367665 246820
rect 360512 246762 367604 246818
rect 367660 246762 367665 246818
rect 360512 246760 367665 246762
rect 360512 246758 360518 246760
rect 367599 246757 367665 246760
rect 367738 246758 367744 246822
rect 367808 246758 367814 246822
rect 367983 246820 368049 246823
rect 368130 246820 368190 247056
rect 368514 246822 368574 247204
rect 369090 247116 369150 247352
rect 369666 247352 406336 247412
rect 369090 247056 369342 247116
rect 369282 246822 369342 247056
rect 369666 246968 369726 247352
rect 406330 247350 406336 247352
rect 406400 247350 406406 247414
rect 407098 247264 407104 247266
rect 370242 247204 407104 247264
rect 370242 247116 370302 247204
rect 407098 247202 407104 247204
rect 407168 247202 407174 247266
rect 401338 247116 401344 247118
rect 369426 246908 369726 246968
rect 369906 247056 370302 247116
rect 370434 247056 401344 247116
rect 369426 246823 369486 246908
rect 369906 246823 369966 247056
rect 367983 246818 368190 246820
rect 367983 246762 367988 246818
rect 368044 246762 368190 246818
rect 367983 246760 368190 246762
rect 367983 246757 368049 246760
rect 368506 246758 368512 246822
rect 368576 246758 368582 246822
rect 369274 246758 369280 246822
rect 369344 246758 369350 246822
rect 369423 246818 369489 246823
rect 369423 246762 369428 246818
rect 369484 246762 369489 246818
rect 369423 246757 369489 246762
rect 369903 246818 369969 246823
rect 369903 246762 369908 246818
rect 369964 246762 369969 246818
rect 369903 246757 369969 246762
rect 370191 246820 370257 246823
rect 370434 246820 370494 247056
rect 401338 247054 401344 247056
rect 401408 247054 401414 247118
rect 401530 247054 401536 247118
rect 401600 247116 401606 247118
rect 406138 247116 406144 247118
rect 401600 247056 406144 247116
rect 401600 247054 401606 247056
rect 406138 247054 406144 247056
rect 406208 247054 406214 247118
rect 404410 246968 404416 246970
rect 370818 246908 392574 246968
rect 370191 246818 370494 246820
rect 370191 246762 370196 246818
rect 370252 246762 370494 246818
rect 370191 246760 370494 246762
rect 370671 246820 370737 246823
rect 370818 246820 370878 246908
rect 392514 246823 392574 246908
rect 393090 246908 404416 246968
rect 370671 246818 370878 246820
rect 370671 246762 370676 246818
rect 370732 246762 370878 246818
rect 370671 246760 370878 246762
rect 377199 246820 377265 246823
rect 388239 246820 388305 246823
rect 377199 246818 388305 246820
rect 377199 246762 377204 246818
rect 377260 246762 388244 246818
rect 388300 246762 388305 246818
rect 377199 246760 388305 246762
rect 392514 246818 392625 246823
rect 392514 246762 392564 246818
rect 392620 246762 392625 246818
rect 392514 246760 392625 246762
rect 370191 246757 370257 246760
rect 370671 246757 370737 246760
rect 377199 246757 377265 246760
rect 388239 246757 388305 246760
rect 392559 246757 392625 246760
rect 392943 246820 393009 246823
rect 393090 246820 393150 246908
rect 404410 246906 404416 246908
rect 404480 246906 404486 246970
rect 392943 246818 393150 246820
rect 392943 246762 392948 246818
rect 393004 246762 393150 246818
rect 392943 246760 393150 246762
rect 393423 246820 393489 246823
rect 674746 246820 674752 246822
rect 393423 246818 674752 246820
rect 393423 246762 393428 246818
rect 393484 246762 674752 246818
rect 393423 246760 674752 246762
rect 392943 246757 393009 246760
rect 393423 246757 393489 246760
rect 674746 246758 674752 246760
rect 674816 246758 674822 246822
rect 177039 246670 187902 246672
rect 177039 246614 177044 246670
rect 177100 246614 187902 246670
rect 177039 246612 187902 246614
rect 187983 246672 188049 246675
rect 211599 246672 211665 246675
rect 187983 246670 211665 246672
rect 187983 246614 187988 246670
rect 188044 246614 211604 246670
rect 211660 246614 211665 246670
rect 187983 246612 211665 246614
rect 177039 246609 177105 246612
rect 187983 246609 188049 246612
rect 211599 246609 211665 246612
rect 65103 246524 65169 246527
rect 202095 246524 202161 246527
rect 65103 246522 202161 246524
rect 65103 246466 65108 246522
rect 65164 246466 202100 246522
rect 202156 246466 202161 246522
rect 65103 246464 202161 246466
rect 65103 246461 65169 246464
rect 202095 246461 202161 246464
rect 211407 246376 211473 246379
rect 87618 246316 106686 246376
rect 65199 245932 65265 245935
rect 87618 245932 87678 246316
rect 106626 246228 106686 246316
rect 187650 246374 211473 246376
rect 187650 246318 211412 246374
rect 211468 246318 211473 246374
rect 187650 246316 211473 246318
rect 171759 246228 171825 246231
rect 187650 246228 187710 246316
rect 211407 246313 211473 246316
rect 211311 246228 211377 246231
rect 106626 246226 171825 246228
rect 106626 246170 171764 246226
rect 171820 246170 171825 246226
rect 106626 246168 171825 246170
rect 171759 246165 171825 246168
rect 177090 246168 187710 246228
rect 187842 246226 211377 246228
rect 187842 246170 211316 246226
rect 211372 246170 211377 246226
rect 187842 246168 211377 246170
rect 166863 246080 166929 246083
rect 177090 246080 177150 246168
rect 187842 246080 187902 246168
rect 211311 246165 211377 246168
rect 211119 246080 211185 246083
rect 166863 246078 177150 246080
rect 166863 246022 166868 246078
rect 166924 246022 177150 246078
rect 166863 246020 177150 246022
rect 177282 246020 187902 246080
rect 210738 246078 211185 246080
rect 210738 246022 211124 246078
rect 211180 246022 211185 246078
rect 210738 246020 211185 246022
rect 166863 246017 166929 246020
rect 65199 245930 87678 245932
rect 42306 245639 42366 245902
rect 65199 245874 65204 245930
rect 65260 245874 87678 245930
rect 65199 245872 87678 245874
rect 163983 245932 164049 245935
rect 177039 245932 177105 245935
rect 163983 245930 177105 245932
rect 163983 245874 163988 245930
rect 164044 245874 177044 245930
rect 177100 245874 177105 245930
rect 163983 245872 177105 245874
rect 65199 245869 65265 245872
rect 163983 245869 164049 245872
rect 177039 245869 177105 245872
rect 172719 245784 172785 245787
rect 177282 245784 177342 246020
rect 210738 245932 210798 246020
rect 211119 246017 211185 246020
rect 211023 245932 211089 245935
rect 674799 245934 674865 245935
rect 674746 245932 674752 245934
rect 172719 245782 177342 245784
rect 172719 245726 172724 245782
rect 172780 245726 177342 245782
rect 172719 245724 177342 245726
rect 177474 245872 210798 245932
rect 210882 245930 211089 245932
rect 210882 245874 211028 245930
rect 211084 245874 211089 245930
rect 210882 245872 211089 245874
rect 674708 245872 674752 245932
rect 674816 245930 674865 245934
rect 674860 245874 674865 245930
rect 172719 245721 172785 245724
rect 42306 245634 42417 245639
rect 42306 245578 42356 245634
rect 42412 245578 42417 245634
rect 42306 245576 42417 245578
rect 42351 245573 42417 245576
rect 175503 245636 175569 245639
rect 177474 245636 177534 245872
rect 178383 245784 178449 245787
rect 210882 245784 210942 245872
rect 211023 245869 211089 245872
rect 674746 245870 674752 245872
rect 674816 245870 674865 245874
rect 674799 245869 674865 245870
rect 178383 245782 210942 245784
rect 178383 245726 178388 245782
rect 178444 245726 210942 245782
rect 178383 245724 210942 245726
rect 178383 245721 178449 245724
rect 175503 245634 177534 245636
rect 175503 245578 175508 245634
rect 175564 245578 177534 245634
rect 175503 245576 177534 245578
rect 181359 245636 181425 245639
rect 210735 245636 210801 245639
rect 181359 245634 210801 245636
rect 181359 245578 181364 245634
rect 181420 245578 210740 245634
rect 210796 245578 210801 245634
rect 181359 245576 210801 245578
rect 175503 245573 175569 245576
rect 181359 245573 181425 245576
rect 210735 245573 210801 245576
rect 181263 245488 181329 245491
rect 186831 245488 186897 245491
rect 181263 245486 186897 245488
rect 181263 245430 181268 245486
rect 181324 245430 186836 245486
rect 186892 245430 186897 245486
rect 181263 245428 186897 245430
rect 181263 245425 181329 245428
rect 186831 245425 186897 245428
rect 187023 245488 187089 245491
rect 210543 245488 210609 245491
rect 187023 245486 210609 245488
rect 187023 245430 187028 245486
rect 187084 245430 210548 245486
rect 210604 245430 210609 245486
rect 187023 245428 210609 245430
rect 187023 245425 187089 245428
rect 210543 245425 210609 245428
rect 158319 245340 158385 245343
rect 168591 245340 168657 245343
rect 158319 245338 168657 245340
rect 158319 245282 158324 245338
rect 158380 245282 168596 245338
rect 168652 245282 168657 245338
rect 158319 245280 168657 245282
rect 158319 245277 158385 245280
rect 168591 245277 168657 245280
rect 171759 245340 171825 245343
rect 187983 245340 188049 245343
rect 202191 245340 202257 245343
rect 171759 245338 187902 245340
rect 171759 245282 171764 245338
rect 171820 245282 187902 245338
rect 171759 245280 187902 245282
rect 171759 245277 171825 245280
rect 171663 245192 171729 245195
rect 187695 245192 187761 245195
rect 171663 245190 187761 245192
rect 171663 245134 171668 245190
rect 171724 245134 187700 245190
rect 187756 245134 187761 245190
rect 171663 245132 187761 245134
rect 187842 245192 187902 245280
rect 187983 245338 202257 245340
rect 187983 245282 187988 245338
rect 188044 245282 202196 245338
rect 202252 245282 202257 245338
rect 187983 245280 202257 245282
rect 187983 245277 188049 245280
rect 202191 245277 202257 245280
rect 210298 245192 210304 245194
rect 187842 245132 210304 245192
rect 171663 245129 171729 245132
rect 187695 245129 187761 245132
rect 210298 245130 210304 245132
rect 210368 245130 210374 245194
rect 674895 245192 674961 245195
rect 675471 245194 675537 245195
rect 675471 245192 675520 245194
rect 674895 245190 675520 245192
rect 674895 245134 674900 245190
rect 674956 245134 675476 245190
rect 674895 245132 675520 245134
rect 674895 245129 674961 245132
rect 675471 245130 675520 245132
rect 675584 245130 675590 245194
rect 675471 245129 675537 245130
rect 187023 245044 187089 245047
rect 227055 245044 227121 245047
rect 187023 245042 227121 245044
rect 187023 244986 187028 245042
rect 187084 244986 227060 245042
rect 227116 244986 227121 245042
rect 187023 244984 227121 244986
rect 187023 244981 187089 244984
rect 227055 244981 227121 244984
rect 228111 245044 228177 245047
rect 247503 245044 247569 245047
rect 228111 245042 247569 245044
rect 228111 244986 228116 245042
rect 228172 244986 247508 245042
rect 247564 244986 247569 245042
rect 228111 244984 247569 244986
rect 228111 244981 228177 244984
rect 247503 244981 247569 244984
rect 247695 245044 247761 245047
rect 287919 245044 287985 245047
rect 247695 245042 287985 245044
rect 247695 244986 247700 245042
rect 247756 244986 287924 245042
rect 287980 244986 287985 245042
rect 247695 244984 287985 244986
rect 247695 244981 247761 244984
rect 287919 244981 287985 244984
rect 288111 245044 288177 245047
rect 290031 245044 290097 245047
rect 288111 245042 290097 245044
rect 288111 244986 288116 245042
rect 288172 244986 290036 245042
rect 290092 244986 290097 245042
rect 288111 244984 290097 244986
rect 288111 244981 288177 244984
rect 290031 244981 290097 244984
rect 292335 245044 292401 245047
rect 307791 245044 307857 245047
rect 292335 245042 307857 245044
rect 292335 244986 292340 245042
rect 292396 244986 307796 245042
rect 307852 244986 307857 245042
rect 292335 244984 307857 244986
rect 292335 244981 292401 244984
rect 307791 244981 307857 244984
rect 307983 245044 308049 245047
rect 308175 245044 308241 245047
rect 307983 245042 308241 245044
rect 307983 244986 307988 245042
rect 308044 244986 308180 245042
rect 308236 244986 308241 245042
rect 307983 244984 308241 244986
rect 307983 244981 308049 244984
rect 308175 244981 308241 244984
rect 309423 245044 309489 245047
rect 326799 245044 326865 245047
rect 309423 245042 326865 245044
rect 309423 244986 309428 245042
rect 309484 244986 326804 245042
rect 326860 244986 326865 245042
rect 309423 244984 326865 244986
rect 309423 244981 309489 244984
rect 326799 244981 326865 244984
rect 328239 245044 328305 245047
rect 328431 245044 328497 245047
rect 328239 245042 328497 245044
rect 328239 244986 328244 245042
rect 328300 244986 328436 245042
rect 328492 244986 328497 245042
rect 328239 244984 328497 244986
rect 328239 244981 328305 244984
rect 328431 244981 328497 244984
rect 328623 245044 328689 245047
rect 348207 245044 348273 245047
rect 328623 245042 348273 245044
rect 328623 244986 328628 245042
rect 328684 244986 348212 245042
rect 348268 244986 348273 245042
rect 328623 244984 348273 244986
rect 328623 244981 328689 244984
rect 348207 244981 348273 244984
rect 348879 245044 348945 245047
rect 368367 245044 368433 245047
rect 348879 245042 368433 245044
rect 348879 244986 348884 245042
rect 348940 244986 368372 245042
rect 368428 244986 368433 245042
rect 348879 244984 368433 244986
rect 348879 244981 348945 244984
rect 368367 244981 368433 244984
rect 369039 245044 369105 245047
rect 388527 245044 388593 245047
rect 369039 245042 388593 245044
rect 369039 244986 369044 245042
rect 369100 244986 388532 245042
rect 388588 244986 388593 245042
rect 369039 244984 388593 244986
rect 369039 244981 369105 244984
rect 388527 244981 388593 244984
rect 388719 245044 388785 245047
rect 388858 245044 388864 245046
rect 388719 245042 388864 245044
rect 388719 244986 388724 245042
rect 388780 244986 388864 245042
rect 388719 244984 388864 244986
rect 388719 244981 388785 244984
rect 388858 244982 388864 244984
rect 388928 244982 388934 245046
rect 389007 245044 389073 245047
rect 401338 245044 401344 245046
rect 389007 245042 401344 245044
rect 389007 244986 389012 245042
rect 389068 244986 401344 245042
rect 389007 244984 401344 244986
rect 389007 244981 389073 244984
rect 401338 244982 401344 244984
rect 401408 244982 401414 245046
rect 401487 245044 401553 245047
rect 401914 245044 401920 245046
rect 401487 245042 401920 245044
rect 401487 244986 401492 245042
rect 401548 244986 401920 245042
rect 401487 244984 401920 244986
rect 401487 244981 401553 244984
rect 401914 244982 401920 244984
rect 401984 244982 401990 245046
rect 403311 245044 403377 245047
rect 404218 245044 404224 245046
rect 403311 245042 404224 245044
rect 403311 244986 403316 245042
rect 403372 244986 404224 245042
rect 403311 244984 404224 244986
rect 403311 244981 403377 244984
rect 404218 244982 404224 244984
rect 404288 244982 404294 245046
rect 404367 245044 404433 245047
rect 404986 245044 404992 245046
rect 404367 245042 404992 245044
rect 404367 244986 404372 245042
rect 404428 244986 404992 245042
rect 404367 244984 404992 244986
rect 404367 244981 404433 244984
rect 404986 244982 404992 244984
rect 405056 244982 405062 245046
rect 405135 245044 405201 245047
rect 406906 245044 406912 245046
rect 405135 245042 406912 245044
rect 405135 244986 405140 245042
rect 405196 244986 406912 245042
rect 405135 244984 406912 244986
rect 405135 244981 405201 244984
rect 406906 244982 406912 244984
rect 406976 244982 406982 245046
rect 407055 245044 407121 245047
rect 409018 245044 409024 245046
rect 407055 245042 409024 245044
rect 407055 244986 407060 245042
rect 407116 244986 409024 245042
rect 407055 244984 409024 244986
rect 407055 244981 407121 244984
rect 409018 244982 409024 244984
rect 409088 244982 409094 245046
rect 409167 245044 409233 245047
rect 409402 245044 409408 245046
rect 409167 245042 409408 245044
rect 409167 244986 409172 245042
rect 409228 244986 409408 245042
rect 409167 244984 409408 244986
rect 409167 244981 409233 244984
rect 409402 244982 409408 244984
rect 409472 244982 409478 245046
rect 42106 244834 42112 244898
rect 42176 244896 42182 244898
rect 674895 244896 674961 244899
rect 42176 244894 674961 244896
rect 42176 244838 674900 244894
rect 674956 244838 674961 244894
rect 42176 244836 674961 244838
rect 42176 244834 42182 244836
rect 674895 244833 674961 244836
rect 202095 244748 202161 244751
rect 211215 244748 211281 244751
rect 202095 244746 211281 244748
rect 202095 244690 202100 244746
rect 202156 244690 211220 244746
rect 211276 244690 211281 244746
rect 202095 244688 211281 244690
rect 202095 244685 202161 244688
rect 211215 244685 211281 244688
rect 211407 244748 211473 244751
rect 226383 244748 226449 244751
rect 211407 244746 226449 244748
rect 211407 244690 211412 244746
rect 211468 244690 226388 244746
rect 226444 244690 226449 244746
rect 211407 244688 226449 244690
rect 211407 244685 211473 244688
rect 226383 244685 226449 244688
rect 227439 244748 227505 244751
rect 227631 244748 227697 244751
rect 227439 244746 227697 244748
rect 227439 244690 227444 244746
rect 227500 244690 227636 244746
rect 227692 244690 227697 244746
rect 227439 244688 227697 244690
rect 227439 244685 227505 244688
rect 227631 244685 227697 244688
rect 228207 244748 228273 244751
rect 247354 244748 247360 244750
rect 228207 244746 247360 244748
rect 228207 244690 228212 244746
rect 228268 244690 247360 244746
rect 228207 244688 247360 244690
rect 228207 244685 228273 244688
rect 247354 244686 247360 244688
rect 247424 244686 247430 244750
rect 247503 244748 247569 244751
rect 247695 244748 247761 244751
rect 247503 244746 247761 244748
rect 247503 244690 247508 244746
rect 247564 244690 247700 244746
rect 247756 244690 247761 244746
rect 247503 244688 247761 244690
rect 247503 244685 247569 244688
rect 247695 244685 247761 244688
rect 257679 244748 257745 244751
rect 344463 244748 344529 244751
rect 257679 244746 344529 244748
rect 257679 244690 257684 244746
rect 257740 244690 344468 244746
rect 344524 244690 344529 244746
rect 257679 244688 344529 244690
rect 257679 244685 257745 244688
rect 344463 244685 344529 244688
rect 348591 244748 348657 244751
rect 369135 244748 369201 244751
rect 348591 244746 369201 244748
rect 348591 244690 348596 244746
rect 348652 244690 369140 244746
rect 369196 244690 369201 244746
rect 348591 244688 369201 244690
rect 348591 244685 348657 244688
rect 369135 244685 369201 244688
rect 388527 244748 388593 244751
rect 400762 244748 400768 244750
rect 388527 244746 400768 244748
rect 388527 244690 388532 244746
rect 388588 244690 400768 244746
rect 388527 244688 400768 244690
rect 388527 244685 388593 244688
rect 400762 244686 400768 244688
rect 400832 244686 400838 244750
rect 400911 244748 400977 244751
rect 401146 244748 401152 244750
rect 400911 244746 401152 244748
rect 400911 244690 400916 244746
rect 400972 244690 401152 244746
rect 400911 244688 401152 244690
rect 400911 244685 400977 244688
rect 401146 244686 401152 244688
rect 401216 244686 401222 244750
rect 403887 244748 403953 244751
rect 404026 244748 404032 244750
rect 403887 244746 404032 244748
rect 403887 244690 403892 244746
rect 403948 244690 404032 244746
rect 403887 244688 404032 244690
rect 403887 244685 403953 244688
rect 404026 244686 404032 244688
rect 404096 244686 404102 244750
rect 404367 244748 404433 244751
rect 404602 244748 404608 244750
rect 404367 244746 404608 244748
rect 404367 244690 404372 244746
rect 404428 244690 404608 244746
rect 404367 244688 404608 244690
rect 404367 244685 404433 244688
rect 404602 244686 404608 244688
rect 404672 244686 404678 244750
rect 673359 244748 673425 244751
rect 674170 244748 674176 244750
rect 673359 244746 674176 244748
rect 673359 244690 673364 244746
rect 673420 244690 674176 244746
rect 673359 244688 674176 244690
rect 673359 244685 673425 244688
rect 674170 244686 674176 244688
rect 674240 244686 674246 244750
rect 212079 244600 212145 244603
rect 227535 244600 227601 244603
rect 212079 244598 227601 244600
rect 212079 244542 212084 244598
rect 212140 244542 227540 244598
rect 227596 244542 227601 244598
rect 212079 244540 227601 244542
rect 212079 244537 212145 244540
rect 227535 244537 227601 244540
rect 229551 244600 229617 244603
rect 328378 244600 328384 244602
rect 229551 244598 328384 244600
rect 229551 244542 229556 244598
rect 229612 244542 328384 244598
rect 229551 244540 328384 244542
rect 229551 244537 229617 244540
rect 328378 244538 328384 244540
rect 328448 244538 328454 244602
rect 348399 244600 348465 244603
rect 328578 244598 348465 244600
rect 328578 244542 348404 244598
rect 348460 244542 348465 244598
rect 328578 244540 348465 244542
rect 221007 244452 221073 244455
rect 308079 244452 308145 244455
rect 221007 244450 308145 244452
rect 221007 244394 221012 244450
rect 221068 244394 308084 244450
rect 308140 244394 308145 244450
rect 221007 244392 308145 244394
rect 221007 244389 221073 244392
rect 308079 244389 308145 244392
rect 308271 244452 308337 244455
rect 328578 244452 328638 244540
rect 348399 244537 348465 244540
rect 368463 244600 368529 244603
rect 368847 244600 368913 244603
rect 403791 244602 403857 244603
rect 368463 244598 368913 244600
rect 368463 244542 368468 244598
rect 368524 244542 368852 244598
rect 368908 244542 368913 244598
rect 368463 244540 368913 244542
rect 368463 244537 368529 244540
rect 368847 244537 368913 244540
rect 369274 244538 369280 244602
rect 369344 244600 369350 244602
rect 399994 244600 400000 244602
rect 369344 244540 400000 244600
rect 369344 244538 369350 244540
rect 399994 244538 400000 244540
rect 400064 244538 400070 244602
rect 403791 244600 403840 244602
rect 403748 244598 403840 244600
rect 403748 244542 403796 244598
rect 403748 244540 403840 244542
rect 403791 244538 403840 244540
rect 403904 244538 403910 244602
rect 673839 244600 673905 244603
rect 675130 244600 675136 244602
rect 673839 244598 675136 244600
rect 673839 244542 673844 244598
rect 673900 244542 675136 244598
rect 673839 244540 675136 244542
rect 403791 244537 403857 244538
rect 673839 244537 673905 244540
rect 675130 244538 675136 244540
rect 675200 244538 675206 244602
rect 308271 244450 328638 244452
rect 308271 244394 308276 244450
rect 308332 244394 328638 244450
rect 308271 244392 328638 244394
rect 328719 244452 328785 244455
rect 368559 244452 368625 244455
rect 328719 244450 368625 244452
rect 328719 244394 328724 244450
rect 328780 244394 368564 244450
rect 368620 244394 368625 244450
rect 328719 244392 368625 244394
rect 308271 244389 308337 244392
rect 328719 244389 328785 244392
rect 368559 244389 368625 244392
rect 368698 244390 368704 244454
rect 368768 244452 368774 244454
rect 400186 244452 400192 244454
rect 368768 244392 400192 244452
rect 368768 244390 368774 244392
rect 400186 244390 400192 244392
rect 400256 244390 400262 244454
rect 257583 244304 257649 244307
rect 343791 244304 343857 244307
rect 257583 244302 343857 244304
rect 257583 244246 257588 244302
rect 257644 244246 343796 244302
rect 343852 244246 343857 244302
rect 257583 244244 343857 244246
rect 257583 244241 257649 244244
rect 343791 244241 343857 244244
rect 367738 244242 367744 244306
rect 367808 244304 367814 244306
rect 400570 244304 400576 244306
rect 367808 244244 400576 244304
rect 367808 244242 367814 244244
rect 400570 244242 400576 244244
rect 400640 244242 400646 244306
rect 225807 244156 225873 244159
rect 257679 244156 257745 244159
rect 225807 244154 257745 244156
rect 225807 244098 225812 244154
rect 225868 244098 257684 244154
rect 257740 244098 257745 244154
rect 225807 244096 257745 244098
rect 225807 244093 225873 244096
rect 257679 244093 257745 244096
rect 257871 244156 257937 244159
rect 343311 244156 343377 244159
rect 257871 244154 343377 244156
rect 257871 244098 257876 244154
rect 257932 244098 343316 244154
rect 343372 244098 343377 244154
rect 257871 244096 343377 244098
rect 257871 244093 257937 244096
rect 343311 244093 343377 244096
rect 369135 244156 369201 244159
rect 400378 244156 400384 244158
rect 369135 244154 400384 244156
rect 369135 244098 369140 244154
rect 369196 244098 400384 244154
rect 369135 244096 400384 244098
rect 369135 244093 369201 244096
rect 400378 244094 400384 244096
rect 400448 244094 400454 244158
rect 219759 244008 219825 244011
rect 341583 244008 341649 244011
rect 219759 244006 341649 244008
rect 219759 243950 219764 244006
rect 219820 243950 341588 244006
rect 341644 243950 341649 244006
rect 219759 243948 341649 243950
rect 219759 243945 219825 243948
rect 341583 243945 341649 243948
rect 388858 243946 388864 244010
rect 388928 244008 388934 244010
rect 403258 244008 403264 244010
rect 388928 243948 403264 244008
rect 388928 243946 388934 243948
rect 403258 243946 403264 243948
rect 403328 243946 403334 244010
rect 218223 243860 218289 243863
rect 341103 243860 341169 243863
rect 218223 243858 341169 243860
rect 218223 243802 218228 243858
rect 218284 243802 341108 243858
rect 341164 243802 341169 243858
rect 218223 243800 341169 243802
rect 218223 243797 218289 243800
rect 341103 243797 341169 243800
rect 212367 243712 212433 243715
rect 335151 243712 335217 243715
rect 212367 243710 335217 243712
rect 212367 243654 212372 243710
rect 212428 243654 335156 243710
rect 335212 243654 335217 243710
rect 212367 243652 335217 243654
rect 212367 243649 212433 243652
rect 335151 243649 335217 243652
rect 214287 243564 214353 243567
rect 328431 243564 328497 243567
rect 214287 243562 328497 243564
rect 214287 243506 214292 243562
rect 214348 243506 328436 243562
rect 328492 243506 328497 243562
rect 214287 243504 328497 243506
rect 214287 243501 214353 243504
rect 328431 243501 328497 243504
rect 328570 243502 328576 243566
rect 328640 243564 328646 243566
rect 345999 243564 346065 243567
rect 328640 243562 346065 243564
rect 328640 243506 346004 243562
rect 346060 243506 346065 243562
rect 328640 243504 346065 243506
rect 328640 243502 328646 243504
rect 345999 243501 346065 243504
rect 674554 243502 674560 243566
rect 674624 243564 674630 243566
rect 675471 243564 675537 243567
rect 674624 243562 675537 243564
rect 674624 243506 675476 243562
rect 675532 243506 675537 243562
rect 674624 243504 675537 243506
rect 674624 243502 674630 243504
rect 675471 243501 675537 243504
rect 207279 243416 207345 243419
rect 385263 243416 385329 243419
rect 207279 243414 385329 243416
rect 207279 243358 207284 243414
rect 207340 243358 385268 243414
rect 385324 243358 385329 243414
rect 207279 243356 385329 243358
rect 207279 243353 207345 243356
rect 385263 243353 385329 243356
rect 232335 243268 232401 243271
rect 347727 243268 347793 243271
rect 232335 243266 347793 243268
rect 232335 243210 232340 243266
rect 232396 243210 347732 243266
rect 347788 243210 347793 243266
rect 232335 243208 347793 243210
rect 232335 243205 232401 243208
rect 347727 243205 347793 243208
rect 224559 243120 224625 243123
rect 257583 243120 257649 243123
rect 224559 243118 257649 243120
rect 224559 243062 224564 243118
rect 224620 243062 257588 243118
rect 257644 243062 257649 243118
rect 224559 243060 257649 243062
rect 224559 243057 224625 243060
rect 257583 243057 257649 243060
rect 296655 243120 296721 243123
rect 297231 243120 297297 243123
rect 296655 243118 297297 243120
rect 296655 243062 296660 243118
rect 296716 243062 297236 243118
rect 297292 243062 297297 243118
rect 296655 243060 297297 243062
rect 296655 243057 296721 243060
rect 297231 243057 297297 243060
rect 308175 243120 308241 243123
rect 342543 243120 342609 243123
rect 308175 243118 342609 243120
rect 308175 243062 308180 243118
rect 308236 243062 342548 243118
rect 342604 243062 342609 243118
rect 308175 243060 342609 243062
rect 308175 243057 308241 243060
rect 342543 243057 342609 243060
rect 223023 242972 223089 242975
rect 257871 242972 257937 242975
rect 223023 242970 257937 242972
rect 223023 242914 223028 242970
rect 223084 242914 257876 242970
rect 257932 242914 257937 242970
rect 223023 242912 257937 242914
rect 223023 242909 223089 242912
rect 257871 242909 257937 242912
rect 296751 242972 296817 242975
rect 305775 242972 305841 242975
rect 296751 242970 305841 242972
rect 296751 242914 296756 242970
rect 296812 242914 305780 242970
rect 305836 242914 305841 242970
rect 296751 242912 305841 242914
rect 296751 242909 296817 242912
rect 305775 242909 305841 242912
rect 328431 242972 328497 242975
rect 348399 242972 348465 242975
rect 328431 242970 348465 242972
rect 328431 242914 328436 242970
rect 328492 242914 348404 242970
rect 348460 242914 348465 242970
rect 328431 242912 348465 242914
rect 328431 242909 328497 242912
rect 348399 242909 348465 242912
rect 41914 242614 41920 242678
rect 41984 242676 41990 242678
rect 42874 242676 42880 242678
rect 41984 242616 42880 242676
rect 41984 242614 41990 242616
rect 42874 242614 42880 242616
rect 42944 242614 42950 242678
rect 285135 242676 285201 242679
rect 297903 242676 297969 242679
rect 285135 242674 297969 242676
rect 285135 242618 285140 242674
rect 285196 242618 297908 242674
rect 297964 242618 297969 242674
rect 285135 242616 297969 242618
rect 285135 242613 285201 242616
rect 297903 242613 297969 242616
rect 290703 242528 290769 242531
rect 298191 242528 298257 242531
rect 290703 242526 298257 242528
rect 290703 242470 290708 242526
rect 290764 242470 298196 242526
rect 298252 242470 298257 242526
rect 290703 242468 298257 242470
rect 290703 242465 290769 242468
rect 298191 242465 298257 242468
rect 157935 242380 158001 242383
rect 161199 242380 161265 242383
rect 140832 242378 158001 242380
rect 140832 242322 157940 242378
rect 157996 242322 158001 242378
rect 140832 242320 158001 242322
rect 157935 242317 158001 242320
rect 161154 242378 161265 242380
rect 161154 242322 161204 242378
rect 161260 242322 161265 242378
rect 161154 242317 161265 242322
rect 283215 242380 283281 242383
rect 290799 242380 290865 242383
rect 283215 242378 290865 242380
rect 283215 242322 283220 242378
rect 283276 242322 290804 242378
rect 290860 242322 290865 242378
rect 283215 242320 290865 242322
rect 283215 242317 283281 242320
rect 290799 242317 290865 242320
rect 297519 242380 297585 242383
rect 297999 242380 298065 242383
rect 297519 242378 298065 242380
rect 297519 242322 297524 242378
rect 297580 242322 298004 242378
rect 298060 242322 298065 242378
rect 297519 242320 298065 242322
rect 297519 242317 297585 242320
rect 297999 242317 298065 242320
rect 161154 242087 161214 242317
rect 282543 242232 282609 242235
rect 292431 242232 292497 242235
rect 282543 242230 292497 242232
rect 282543 242174 282548 242230
rect 282604 242174 292436 242230
rect 292492 242174 292497 242230
rect 282543 242172 292497 242174
rect 282543 242169 282609 242172
rect 292431 242169 292497 242172
rect 509775 242232 509841 242235
rect 673839 242232 673905 242235
rect 509775 242230 673905 242232
rect 509775 242174 509780 242230
rect 509836 242174 673844 242230
rect 673900 242174 673905 242230
rect 509775 242172 673905 242174
rect 509775 242169 509841 242172
rect 673839 242169 673905 242172
rect 40239 242084 40305 242087
rect 41722 242084 41728 242086
rect 40239 242082 41728 242084
rect 40239 242026 40244 242082
rect 40300 242026 41728 242082
rect 40239 242024 41728 242026
rect 40239 242021 40305 242024
rect 41722 242022 41728 242024
rect 41792 242022 41798 242086
rect 161154 242082 161265 242087
rect 161154 242026 161204 242082
rect 161260 242026 161265 242082
rect 161154 242024 161265 242026
rect 161199 242021 161265 242024
rect 235695 242084 235761 242087
rect 348879 242084 348945 242087
rect 235695 242082 348945 242084
rect 235695 242026 235700 242082
rect 235756 242026 348884 242082
rect 348940 242026 348945 242082
rect 235695 242024 348945 242026
rect 235695 242021 235761 242024
rect 348879 242021 348945 242024
rect 504015 242084 504081 242087
rect 673359 242084 673425 242087
rect 504015 242082 673425 242084
rect 504015 242026 504020 242082
rect 504076 242026 673364 242082
rect 673420 242026 673425 242082
rect 504015 242024 673425 242026
rect 504015 242021 504081 242024
rect 673359 242021 673425 242024
rect 40378 241874 40384 241938
rect 40448 241936 40454 241938
rect 42298 241936 42304 241938
rect 40448 241876 42304 241936
rect 40448 241874 40454 241876
rect 42298 241874 42304 241876
rect 42368 241874 42374 241938
rect 246159 241936 246225 241939
rect 355023 241936 355089 241939
rect 246159 241934 355089 241936
rect 246159 241878 246164 241934
rect 246220 241878 355028 241934
rect 355084 241878 355089 241934
rect 246159 241876 355089 241878
rect 246159 241873 246225 241876
rect 355023 241873 355089 241876
rect 674895 241936 674961 241939
rect 675322 241936 675328 241938
rect 674895 241934 675328 241936
rect 674895 241878 674900 241934
rect 674956 241878 675328 241934
rect 674895 241876 675328 241878
rect 674895 241873 674961 241876
rect 675322 241874 675328 241876
rect 675392 241874 675398 241938
rect 245391 241788 245457 241791
rect 356751 241788 356817 241791
rect 245391 241786 356817 241788
rect 245391 241730 245396 241786
rect 245452 241730 356756 241786
rect 356812 241730 356817 241786
rect 245391 241728 356817 241730
rect 245391 241725 245457 241728
rect 356751 241725 356817 241728
rect 383055 241790 383121 241791
rect 383055 241786 383104 241790
rect 383168 241788 383174 241790
rect 383055 241730 383060 241786
rect 383055 241726 383104 241730
rect 383168 241728 383212 241788
rect 383168 241726 383174 241728
rect 383055 241725 383121 241726
rect 259983 241640 260049 241643
rect 376143 241640 376209 241643
rect 259983 241638 376209 241640
rect 259983 241582 259988 241638
rect 260044 241582 376148 241638
rect 376204 241582 376209 241638
rect 259983 241580 376209 241582
rect 259983 241577 260049 241580
rect 376143 241577 376209 241580
rect 259599 241492 259665 241495
rect 376815 241492 376881 241495
rect 259599 241490 376881 241492
rect 259599 241434 259604 241490
rect 259660 241434 376820 241490
rect 376876 241434 376881 241490
rect 259599 241432 376881 241434
rect 259599 241429 259665 241432
rect 376815 241429 376881 241432
rect 243951 241344 244017 241347
rect 360015 241344 360081 241347
rect 243951 241342 360081 241344
rect 243951 241286 243956 241342
rect 244012 241286 360020 241342
rect 360076 241286 360081 241342
rect 243951 241284 360081 241286
rect 243951 241281 244017 241284
rect 360015 241281 360081 241284
rect 243183 241196 243249 241199
rect 361551 241196 361617 241199
rect 243183 241194 361617 241196
rect 243183 241138 243188 241194
rect 243244 241138 361556 241194
rect 361612 241138 361617 241194
rect 243183 241136 361617 241138
rect 243183 241133 243249 241136
rect 361551 241133 361617 241136
rect 140802 240604 140862 241092
rect 242703 241048 242769 241051
rect 363087 241048 363153 241051
rect 242703 241046 363153 241048
rect 242703 240990 242708 241046
rect 242764 240990 363092 241046
rect 363148 240990 363153 241046
rect 242703 240988 363153 240990
rect 242703 240985 242769 240988
rect 363087 240985 363153 240988
rect 258639 240900 258705 240903
rect 378831 240900 378897 240903
rect 258639 240898 378897 240900
rect 258639 240842 258644 240898
rect 258700 240842 378836 240898
rect 378892 240842 378897 240898
rect 258639 240840 378897 240842
rect 258639 240837 258705 240840
rect 378831 240837 378897 240840
rect 241743 240752 241809 240755
rect 364815 240752 364881 240755
rect 241743 240750 364881 240752
rect 241743 240694 241748 240750
rect 241804 240694 364820 240750
rect 364876 240694 364881 240750
rect 241743 240692 364881 240694
rect 241743 240689 241809 240692
rect 364815 240689 364881 240692
rect 146319 240604 146385 240607
rect 140802 240602 146385 240604
rect 140802 240546 146324 240602
rect 146380 240546 146385 240602
rect 140802 240544 146385 240546
rect 146319 240541 146385 240544
rect 240975 240604 241041 240607
rect 366543 240604 366609 240607
rect 240975 240602 366609 240604
rect 240975 240546 240980 240602
rect 241036 240546 366548 240602
rect 366604 240546 366609 240602
rect 240975 240544 366609 240546
rect 240975 240541 241041 240544
rect 366543 240541 366609 240544
rect 367599 240604 367665 240607
rect 409743 240604 409809 240607
rect 367599 240602 409809 240604
rect 367599 240546 367604 240602
rect 367660 240546 409748 240602
rect 409804 240546 409809 240602
rect 367599 240544 409809 240546
rect 367599 240541 367665 240544
rect 409743 240541 409809 240544
rect 282255 240456 282321 240459
rect 411471 240456 411537 240459
rect 282255 240454 411537 240456
rect 282255 240398 282260 240454
rect 282316 240398 411476 240454
rect 411532 240398 411537 240454
rect 282255 240396 411537 240398
rect 282255 240393 282321 240396
rect 411471 240393 411537 240396
rect 247119 240308 247185 240311
rect 353967 240308 354033 240311
rect 247119 240306 354033 240308
rect 247119 240250 247124 240306
rect 247180 240250 353972 240306
rect 354028 240250 354033 240306
rect 247119 240248 354033 240250
rect 247119 240245 247185 240248
rect 353967 240245 354033 240248
rect 247599 240160 247665 240163
rect 352239 240160 352305 240163
rect 247599 240158 352305 240160
rect 247599 240102 247604 240158
rect 247660 240102 352244 240158
rect 352300 240102 352305 240158
rect 247599 240100 352305 240102
rect 247599 240097 247665 240100
rect 352239 240097 352305 240100
rect 383055 240160 383121 240163
rect 389871 240160 389937 240163
rect 383055 240158 389937 240160
rect 383055 240102 383060 240158
rect 383116 240102 389876 240158
rect 389932 240102 389937 240158
rect 383055 240100 389937 240102
rect 383055 240097 383121 240100
rect 389871 240097 389937 240100
rect 198927 240012 198993 240015
rect 208719 240012 208785 240015
rect 198927 240010 208785 240012
rect 198927 239954 198932 240010
rect 198988 239954 208724 240010
rect 208780 239954 208785 240010
rect 198927 239952 208785 239954
rect 198927 239949 198993 239952
rect 208719 239949 208785 239952
rect 262575 240012 262641 240015
rect 370959 240012 371025 240015
rect 262575 240010 371025 240012
rect 262575 239954 262580 240010
rect 262636 239954 370964 240010
rect 371020 239954 371025 240010
rect 262575 239952 371025 239954
rect 262575 239949 262641 239952
rect 370959 239949 371025 239952
rect 383055 240012 383121 240015
rect 402351 240012 402417 240015
rect 383055 240010 402417 240012
rect 383055 239954 383060 240010
rect 383116 239954 402356 240010
rect 402412 239954 402417 240010
rect 383055 239952 402417 239954
rect 383055 239949 383121 239952
rect 402351 239949 402417 239952
rect 145402 239864 145408 239866
rect 140832 239804 145408 239864
rect 145402 239802 145408 239804
rect 145472 239802 145478 239866
rect 42351 239420 42417 239423
rect 42351 239418 42558 239420
rect 42351 239362 42356 239418
rect 42412 239362 42558 239418
rect 42351 239360 42558 239362
rect 42351 239357 42417 239360
rect 42498 238979 42558 239360
rect 208719 239124 208785 239127
rect 209871 239124 209937 239127
rect 351375 239124 351441 239127
rect 208719 239122 351441 239124
rect 208719 239066 208724 239122
rect 208780 239066 209876 239122
rect 209932 239066 351380 239122
rect 351436 239066 351441 239122
rect 208719 239064 351441 239066
rect 208719 239061 208785 239064
rect 209871 239061 209937 239064
rect 351375 239061 351441 239064
rect 383055 239126 383121 239127
rect 383055 239122 383104 239126
rect 383168 239124 383174 239126
rect 383055 239066 383060 239122
rect 383055 239062 383104 239066
rect 383168 239064 383212 239124
rect 383168 239062 383174 239064
rect 383055 239061 383121 239062
rect 42447 238974 42558 238979
rect 42447 238918 42452 238974
rect 42508 238918 42558 238974
rect 42447 238916 42558 238918
rect 244335 238976 244401 238979
rect 358959 238976 359025 238979
rect 244335 238974 359025 238976
rect 244335 238918 244340 238974
rect 244396 238918 358964 238974
rect 359020 238918 359025 238974
rect 244335 238916 359025 238918
rect 42447 238913 42513 238916
rect 244335 238913 244401 238916
rect 358959 238913 359025 238916
rect 674799 238976 674865 238979
rect 675514 238976 675520 238978
rect 674799 238974 675520 238976
rect 674799 238918 674804 238974
rect 674860 238918 675520 238974
rect 674799 238916 675520 238918
rect 674799 238913 674865 238916
rect 675514 238914 675520 238916
rect 675584 238914 675590 238978
rect 243567 238828 243633 238831
rect 360687 238828 360753 238831
rect 243567 238826 360753 238828
rect 243567 238770 243572 238826
rect 243628 238770 360692 238826
rect 360748 238770 360753 238826
rect 243567 238768 360753 238770
rect 243567 238765 243633 238768
rect 360687 238765 360753 238768
rect 146703 238680 146769 238683
rect 140832 238678 146769 238680
rect 140832 238622 146708 238678
rect 146764 238622 146769 238678
rect 140832 238620 146769 238622
rect 146703 238617 146769 238620
rect 242799 238680 242865 238683
rect 362703 238680 362769 238683
rect 242799 238678 362769 238680
rect 242799 238622 242804 238678
rect 242860 238622 362708 238678
rect 362764 238622 362769 238678
rect 242799 238620 362769 238622
rect 242799 238617 242865 238620
rect 362703 238617 362769 238620
rect 383055 238680 383121 238683
rect 395343 238680 395409 238683
rect 383055 238678 395409 238680
rect 383055 238622 383060 238678
rect 383116 238622 395348 238678
rect 395404 238622 395409 238678
rect 383055 238620 395409 238622
rect 383055 238617 383121 238620
rect 395343 238617 395409 238620
rect 674938 238618 674944 238682
rect 675008 238680 675014 238682
rect 675471 238680 675537 238683
rect 675008 238678 675537 238680
rect 675008 238622 675476 238678
rect 675532 238622 675537 238678
rect 675008 238620 675537 238622
rect 675008 238618 675014 238620
rect 675471 238617 675537 238620
rect 259023 238532 259089 238535
rect 377679 238532 377745 238535
rect 259023 238530 377745 238532
rect 259023 238474 259028 238530
rect 259084 238474 377684 238530
rect 377740 238474 377745 238530
rect 259023 238472 377745 238474
rect 259023 238469 259089 238472
rect 377679 238469 377745 238472
rect 242319 238384 242385 238387
rect 363855 238384 363921 238387
rect 242319 238382 363921 238384
rect 242319 238326 242324 238382
rect 242380 238326 363860 238382
rect 363916 238326 363921 238382
rect 242319 238324 363921 238326
rect 242319 238321 242385 238324
rect 363855 238321 363921 238324
rect 241359 238236 241425 238239
rect 365775 238236 365841 238239
rect 241359 238234 365841 238236
rect 241359 238178 241364 238234
rect 241420 238178 365780 238234
rect 365836 238178 365841 238234
rect 241359 238176 365841 238178
rect 241359 238173 241425 238176
rect 365775 238173 365841 238176
rect 215823 238088 215889 238091
rect 391407 238088 391473 238091
rect 215823 238086 391473 238088
rect 215823 238030 215828 238086
rect 215884 238030 391412 238086
rect 391468 238030 391473 238086
rect 215823 238028 391473 238030
rect 215823 238025 215889 238028
rect 391407 238025 391473 238028
rect 215247 237940 215313 237943
rect 393135 237940 393201 237943
rect 215247 237938 393201 237940
rect 215247 237882 215252 237938
rect 215308 237882 393140 237938
rect 393196 237882 393201 237938
rect 215247 237880 393201 237882
rect 215247 237877 215313 237880
rect 393135 237877 393201 237880
rect 214863 237792 214929 237795
rect 394671 237792 394737 237795
rect 214863 237790 394737 237792
rect 214863 237734 214868 237790
rect 214924 237734 394676 237790
rect 394732 237734 394737 237790
rect 214863 237732 394737 237734
rect 214863 237729 214929 237732
rect 394671 237729 394737 237732
rect 162735 237644 162801 237647
rect 212986 237644 212992 237646
rect 162735 237642 212992 237644
rect 162735 237586 162740 237642
rect 162796 237586 212992 237642
rect 162735 237584 212992 237586
rect 162735 237581 162801 237584
rect 212986 237582 212992 237584
rect 213056 237582 213062 237646
rect 215919 237644 215985 237647
rect 411951 237644 412017 237647
rect 215919 237642 412017 237644
rect 215919 237586 215924 237642
rect 215980 237586 411956 237642
rect 412012 237586 412017 237642
rect 215919 237584 412017 237586
rect 215919 237581 215985 237584
rect 411951 237581 412017 237584
rect 321903 237496 321969 237499
rect 335343 237496 335409 237499
rect 321903 237494 335409 237496
rect 321903 237438 321908 237494
rect 321964 237438 335348 237494
rect 335404 237438 335409 237494
rect 321903 237436 335409 237438
rect 321903 237433 321969 237436
rect 335343 237433 335409 237436
rect 140802 236904 140862 237392
rect 322287 237348 322353 237351
rect 322767 237348 322833 237351
rect 322287 237346 322833 237348
rect 322287 237290 322292 237346
rect 322348 237290 322772 237346
rect 322828 237290 322833 237346
rect 322287 237288 322833 237290
rect 322287 237285 322353 237288
rect 322767 237285 322833 237288
rect 145551 236904 145617 236907
rect 140802 236902 145617 236904
rect 140802 236846 145556 236902
rect 145612 236846 145617 236902
rect 140802 236844 145617 236846
rect 145551 236841 145617 236844
rect 286863 236904 286929 236907
rect 295887 236904 295953 236907
rect 675759 236906 675825 236907
rect 286863 236902 295953 236904
rect 286863 236846 286868 236902
rect 286924 236846 295892 236902
rect 295948 236846 295953 236902
rect 286863 236844 295953 236846
rect 286863 236841 286929 236844
rect 295887 236841 295953 236844
rect 675706 236842 675712 236906
rect 675776 236904 675825 236906
rect 675776 236902 675868 236904
rect 675820 236846 675868 236902
rect 675776 236844 675868 236846
rect 675776 236842 675825 236844
rect 675759 236841 675825 236842
rect 209775 236756 209841 236759
rect 497487 236756 497553 236759
rect 209775 236754 497553 236756
rect 209775 236698 209780 236754
rect 209836 236698 497492 236754
rect 497548 236698 497553 236754
rect 209775 236696 497553 236698
rect 209775 236693 209841 236696
rect 497487 236693 497553 236696
rect 209679 236608 209745 236611
rect 209679 236606 211710 236608
rect 209679 236550 209684 236606
rect 209740 236550 211710 236606
rect 209679 236548 211710 236550
rect 209679 236545 209745 236548
rect 211650 236460 211710 236548
rect 212986 236546 212992 236610
rect 213056 236608 213062 236610
rect 359247 236608 359313 236611
rect 213056 236606 359313 236608
rect 213056 236550 359252 236606
rect 359308 236550 359313 236606
rect 213056 236548 359313 236550
rect 213056 236546 213062 236548
rect 359247 236545 359313 236548
rect 420591 236460 420657 236463
rect 211650 236458 420657 236460
rect 211650 236402 420596 236458
rect 420652 236402 420657 236458
rect 211650 236400 420657 236402
rect 420591 236397 420657 236400
rect 146799 236312 146865 236315
rect 140802 236310 146865 236312
rect 140802 236254 146804 236310
rect 146860 236254 146865 236310
rect 140802 236252 146865 236254
rect 140802 236210 140862 236252
rect 146799 236249 146865 236252
rect 210298 236250 210304 236314
rect 210368 236312 210374 236314
rect 210927 236312 210993 236315
rect 210368 236310 210993 236312
rect 210368 236254 210932 236310
rect 210988 236254 210993 236310
rect 210368 236252 210993 236254
rect 210368 236250 210374 236252
rect 210927 236249 210993 236252
rect 289359 236312 289425 236315
rect 293775 236312 293841 236315
rect 289359 236310 293841 236312
rect 289359 236254 289364 236310
rect 289420 236254 293780 236310
rect 293836 236254 293841 236310
rect 289359 236252 293841 236254
rect 289359 236249 289425 236252
rect 293775 236249 293841 236252
rect 228591 236164 228657 236167
rect 345615 236164 345681 236167
rect 228591 236162 345681 236164
rect 228591 236106 228596 236162
rect 228652 236106 345620 236162
rect 345676 236106 345681 236162
rect 228591 236104 345681 236106
rect 228591 236101 228657 236104
rect 345615 236101 345681 236104
rect 229743 236016 229809 236019
rect 346575 236016 346641 236019
rect 229743 236014 346641 236016
rect 229743 235958 229748 236014
rect 229804 235958 346580 236014
rect 346636 235958 346641 236014
rect 229743 235956 346641 235958
rect 229743 235953 229809 235956
rect 346575 235953 346641 235956
rect 217167 235868 217233 235871
rect 338991 235868 339057 235871
rect 217167 235866 339057 235868
rect 217167 235810 217172 235866
rect 217228 235810 338996 235866
rect 339052 235810 339057 235866
rect 217167 235808 339057 235810
rect 217167 235805 217233 235808
rect 338991 235805 339057 235808
rect 223983 235720 224049 235723
rect 343407 235720 343473 235723
rect 223983 235718 343473 235720
rect 223983 235662 223988 235718
rect 224044 235662 343412 235718
rect 343468 235662 343473 235718
rect 223983 235660 343473 235662
rect 223983 235657 224049 235660
rect 343407 235657 343473 235660
rect 220815 235572 220881 235575
rect 342159 235572 342225 235575
rect 220815 235570 342225 235572
rect 220815 235514 220820 235570
rect 220876 235514 342164 235570
rect 342220 235514 342225 235570
rect 220815 235512 342225 235514
rect 220815 235509 220881 235512
rect 342159 235509 342225 235512
rect 222159 235424 222225 235427
rect 342927 235424 342993 235427
rect 222159 235422 342993 235424
rect 222159 235366 222164 235422
rect 222220 235366 342932 235422
rect 342988 235366 342993 235422
rect 222159 235364 342993 235366
rect 222159 235361 222225 235364
rect 342927 235361 342993 235364
rect 219183 235276 219249 235279
rect 341199 235276 341265 235279
rect 219183 235274 341265 235276
rect 219183 235218 219188 235274
rect 219244 235218 341204 235274
rect 341260 235218 341265 235274
rect 219183 235216 341265 235218
rect 219183 235213 219249 235216
rect 341199 235213 341265 235216
rect 146415 235128 146481 235131
rect 140832 235126 146481 235128
rect 140832 235070 146420 235126
rect 146476 235070 146481 235126
rect 140832 235068 146481 235070
rect 146415 235065 146481 235068
rect 213231 235128 213297 235131
rect 344367 235128 344433 235131
rect 213231 235126 344433 235128
rect 213231 235070 213236 235126
rect 213292 235070 344372 235126
rect 344428 235070 344433 235126
rect 213231 235068 344433 235070
rect 213231 235065 213297 235068
rect 344367 235065 344433 235068
rect 214959 234980 215025 234983
rect 352239 234980 352305 234983
rect 214959 234978 352305 234980
rect 214959 234922 214964 234978
rect 215020 234922 352244 234978
rect 352300 234922 352305 234978
rect 214959 234920 352305 234922
rect 214959 234917 215025 234920
rect 352239 234917 352305 234920
rect 210159 234832 210225 234835
rect 379407 234832 379473 234835
rect 210159 234830 379473 234832
rect 210159 234774 210164 234830
rect 210220 234774 379412 234830
rect 379468 234774 379473 234830
rect 210159 234772 379473 234774
rect 210159 234769 210225 234772
rect 379407 234769 379473 234772
rect 211450 234622 211456 234686
rect 211520 234684 211526 234686
rect 541455 234684 541521 234687
rect 211520 234682 541521 234684
rect 211520 234626 541460 234682
rect 541516 234626 541521 234682
rect 211520 234624 541521 234626
rect 211520 234622 211526 234624
rect 541455 234621 541521 234624
rect 272943 234536 273009 234539
rect 354447 234536 354513 234539
rect 272943 234534 354513 234536
rect 272943 234478 272948 234534
rect 273004 234478 354452 234534
rect 354508 234478 354513 234534
rect 272943 234476 354513 234478
rect 272943 234473 273009 234476
rect 354447 234473 354513 234476
rect 286767 234388 286833 234391
rect 297423 234388 297489 234391
rect 286767 234386 297489 234388
rect 286767 234330 286772 234386
rect 286828 234330 297428 234386
rect 297484 234330 297489 234386
rect 286767 234328 297489 234330
rect 286767 234325 286833 234328
rect 297423 234325 297489 234328
rect 140802 233648 140862 233840
rect 211887 233796 211953 233799
rect 212026 233796 212032 233798
rect 211887 233794 212032 233796
rect 211887 233738 211892 233794
rect 211948 233738 212032 233794
rect 211887 233736 212032 233738
rect 211887 233733 211953 233736
rect 212026 233734 212032 233736
rect 212096 233734 212102 233798
rect 637306 233734 637312 233798
rect 637376 233796 637382 233798
rect 638127 233796 638193 233799
rect 638703 233796 638769 233799
rect 637376 233794 638769 233796
rect 637376 233738 638132 233794
rect 638188 233738 638708 233794
rect 638764 233738 638769 233794
rect 637376 233736 638769 233738
rect 637376 233734 637382 233736
rect 638127 233733 638193 233736
rect 638703 233733 638769 233736
rect 146799 233648 146865 233651
rect 140802 233646 146865 233648
rect 140802 233590 146804 233646
rect 146860 233590 146865 233646
rect 140802 233588 146865 233590
rect 146799 233585 146865 233588
rect 211023 233650 211089 233651
rect 211023 233646 211072 233650
rect 211136 233648 211142 233650
rect 211311 233648 211377 233651
rect 211695 233650 211761 233651
rect 211642 233648 211648 233650
rect 211023 233590 211028 233646
rect 211023 233586 211072 233590
rect 211136 233588 211180 233648
rect 211311 233646 211648 233648
rect 211712 233648 211761 233650
rect 212175 233650 212241 233651
rect 212175 233648 212224 233650
rect 211712 233646 211804 233648
rect 211311 233590 211316 233646
rect 211372 233590 211648 233646
rect 211756 233590 211804 233646
rect 211311 233588 211648 233590
rect 211136 233586 211142 233588
rect 211023 233585 211089 233586
rect 211311 233585 211377 233588
rect 211642 233586 211648 233588
rect 211712 233588 211804 233590
rect 212132 233646 212224 233648
rect 212132 233590 212180 233646
rect 212132 233588 212224 233590
rect 211712 233586 211761 233588
rect 211695 233585 211761 233586
rect 212175 233586 212224 233588
rect 212288 233586 212294 233650
rect 212410 233586 212416 233650
rect 212480 233648 212486 233650
rect 212986 233648 212992 233650
rect 212480 233588 212992 233648
rect 212480 233586 212486 233588
rect 212986 233586 212992 233588
rect 213056 233586 213062 233650
rect 636922 233586 636928 233650
rect 636992 233648 636998 233650
rect 637071 233648 637137 233651
rect 636992 233646 637137 233648
rect 636992 233590 637076 233646
rect 637132 233590 637137 233646
rect 636992 233588 637137 233590
rect 636992 233586 636998 233588
rect 212175 233585 212241 233586
rect 637071 233585 637137 233588
rect 637498 233586 637504 233650
rect 637568 233648 637574 233650
rect 638511 233648 638577 233651
rect 637568 233646 638577 233648
rect 637568 233590 638516 233646
rect 638572 233590 638577 233646
rect 637568 233588 638577 233590
rect 637568 233586 637574 233588
rect 638511 233585 638577 233588
rect 211407 233500 211473 233503
rect 212986 233500 212992 233502
rect 211407 233498 212992 233500
rect 211407 233442 211412 233498
rect 211468 233442 212992 233498
rect 211407 233440 212992 233442
rect 211407 233437 211473 233440
rect 212986 233438 212992 233440
rect 213056 233438 213062 233502
rect 214287 233498 214353 233503
rect 214287 233442 214292 233498
rect 214348 233442 214353 233498
rect 214287 233437 214353 233442
rect 637114 233438 637120 233502
rect 637184 233500 637190 233502
rect 637551 233500 637617 233503
rect 637935 233502 638001 233503
rect 637184 233498 637617 233500
rect 637184 233442 637556 233498
rect 637612 233442 637617 233498
rect 637184 233440 637617 233442
rect 637184 233438 637190 233440
rect 637551 233437 637617 233440
rect 637882 233438 637888 233502
rect 637952 233500 638001 233502
rect 638991 233500 639057 233503
rect 637952 233498 638044 233500
rect 637996 233442 638044 233498
rect 637952 233440 638044 233442
rect 638658 233498 639057 233500
rect 638658 233442 638996 233498
rect 639052 233442 639057 233498
rect 638658 233440 639057 233442
rect 637952 233438 638001 233440
rect 637935 233437 638001 233438
rect 41146 233290 41152 233354
rect 41216 233352 41222 233354
rect 41775 233352 41841 233355
rect 41216 233350 41841 233352
rect 41216 233294 41780 233350
rect 41836 233294 41841 233350
rect 41216 233292 41841 233294
rect 41216 233290 41222 233292
rect 41775 233289 41841 233292
rect 210874 233290 210880 233354
rect 210944 233352 210950 233354
rect 214290 233352 214350 233437
rect 210944 233292 214350 233352
rect 210944 233290 210950 233292
rect 637690 233290 637696 233354
rect 637760 233352 637766 233354
rect 638658 233352 638718 233440
rect 638991 233437 639057 233440
rect 637760 233292 638718 233352
rect 637760 233290 637766 233292
rect 210298 232846 210304 232910
rect 210368 232908 210374 232910
rect 212410 232908 212416 232910
rect 210368 232848 212416 232908
rect 210368 232846 210374 232848
rect 212410 232846 212416 232848
rect 212480 232846 212486 232910
rect 140802 232168 140862 232656
rect 205551 232316 205617 232319
rect 210498 232316 210558 232656
rect 640386 232464 640446 232656
rect 645711 232464 645777 232467
rect 640386 232462 645777 232464
rect 640386 232406 645716 232462
rect 645772 232406 645777 232462
rect 640386 232404 645777 232406
rect 645711 232401 645777 232404
rect 645135 232316 645201 232319
rect 205551 232314 210558 232316
rect 205551 232258 205556 232314
rect 205612 232258 210558 232314
rect 205551 232256 210558 232258
rect 640194 232314 645201 232316
rect 640194 232258 645140 232314
rect 645196 232258 645201 232314
rect 640194 232256 645201 232258
rect 205551 232253 205617 232256
rect 144399 232168 144465 232171
rect 140802 232166 144465 232168
rect 140802 232110 144404 232166
rect 144460 232110 144465 232166
rect 140802 232108 144465 232110
rect 144399 232105 144465 232108
rect 204879 232168 204945 232171
rect 207375 232168 207441 232171
rect 204879 232166 210528 232168
rect 204879 232110 204884 232166
rect 204940 232110 207380 232166
rect 207436 232110 210528 232166
rect 640194 232138 640254 232256
rect 645135 232253 645201 232256
rect 204879 232108 210528 232110
rect 204879 232105 204945 232108
rect 207375 232105 207441 232108
rect 41967 231726 42033 231727
rect 41914 231662 41920 231726
rect 41984 231724 42033 231726
rect 41984 231722 42076 231724
rect 42028 231666 42076 231722
rect 41984 231664 42076 231666
rect 41984 231662 42033 231664
rect 41967 231661 42033 231662
rect 204783 231576 204849 231579
rect 209583 231576 209649 231579
rect 645135 231576 645201 231579
rect 204783 231574 210528 231576
rect 204783 231518 204788 231574
rect 204844 231518 209588 231574
rect 209644 231518 210528 231574
rect 204783 231516 210528 231518
rect 640416 231574 645201 231576
rect 640416 231518 645140 231574
rect 645196 231518 645201 231574
rect 640416 231516 645201 231518
rect 204783 231513 204849 231516
rect 209583 231513 209649 231516
rect 645135 231513 645201 231516
rect 146799 231428 146865 231431
rect 140832 231426 146865 231428
rect 140832 231370 146804 231426
rect 146860 231370 146865 231426
rect 140832 231368 146865 231370
rect 146799 231365 146865 231368
rect 645135 231132 645201 231135
rect 640386 231130 645201 231132
rect 640386 231074 645140 231130
rect 645196 231074 645201 231130
rect 640386 231072 645201 231074
rect 41967 230984 42033 230987
rect 42106 230984 42112 230986
rect 41922 230982 42112 230984
rect 41922 230926 41972 230982
rect 42028 230926 42112 230982
rect 41922 230924 42112 230926
rect 41922 230921 42033 230924
rect 42106 230922 42112 230924
rect 42176 230922 42182 230986
rect 204687 230984 204753 230987
rect 207951 230984 208017 230987
rect 204687 230982 210528 230984
rect 204687 230926 204692 230982
rect 204748 230926 207956 230982
rect 208012 230926 210528 230982
rect 640386 230954 640446 231072
rect 645135 231069 645201 231072
rect 204687 230924 210528 230926
rect 204687 230921 204753 230924
rect 207951 230921 208017 230924
rect 41775 230394 41841 230395
rect 41722 230392 41728 230394
rect 41684 230332 41728 230392
rect 41792 230390 41841 230394
rect 41836 230334 41841 230390
rect 41722 230330 41728 230332
rect 41792 230330 41841 230334
rect 41775 230329 41841 230330
rect 41722 230182 41728 230246
rect 41792 230244 41798 230246
rect 41922 230244 41982 230921
rect 645135 230688 645201 230691
rect 640194 230686 645201 230688
rect 640194 230630 645140 230686
rect 645196 230630 645201 230686
rect 640194 230628 645201 230630
rect 205935 230540 206001 230543
rect 209391 230540 209457 230543
rect 205935 230538 210528 230540
rect 205935 230482 205940 230538
rect 205996 230482 209396 230538
rect 209452 230482 210528 230538
rect 640194 230510 640254 230628
rect 645135 230625 645201 230628
rect 205935 230480 210528 230482
rect 205935 230477 206001 230480
rect 209391 230477 209457 230480
rect 146703 230244 146769 230247
rect 41792 230184 41982 230244
rect 140832 230242 146769 230244
rect 140832 230186 146708 230242
rect 146764 230186 146769 230242
rect 140832 230184 146769 230186
rect 41792 230182 41798 230184
rect 146703 230181 146769 230184
rect 206799 229948 206865 229951
rect 207087 229948 207153 229951
rect 206799 229946 210528 229948
rect 206799 229890 206804 229946
rect 206860 229890 207092 229946
rect 207148 229890 210528 229946
rect 206799 229888 210528 229890
rect 206799 229885 206865 229888
rect 207087 229885 207153 229888
rect 41338 229738 41344 229802
rect 41408 229800 41414 229802
rect 41775 229800 41841 229803
rect 41408 229798 41841 229800
rect 41408 229742 41780 229798
rect 41836 229742 41841 229798
rect 41408 229740 41841 229742
rect 41408 229738 41414 229740
rect 41775 229737 41841 229740
rect 674415 229504 674481 229507
rect 674415 229502 674784 229504
rect 674415 229446 674420 229502
rect 674476 229446 674784 229502
rect 674415 229444 674784 229446
rect 674415 229441 674481 229444
rect 206127 229356 206193 229359
rect 206127 229354 210528 229356
rect 206127 229298 206132 229354
rect 206188 229298 210528 229354
rect 206127 229296 210528 229298
rect 206127 229293 206193 229296
rect 40954 228998 40960 229062
rect 41024 229060 41030 229062
rect 41775 229060 41841 229063
rect 146799 229060 146865 229063
rect 41024 229058 41841 229060
rect 41024 229002 41780 229058
rect 41836 229002 41841 229058
rect 41024 229000 41841 229002
rect 140832 229058 146865 229060
rect 140832 229002 146804 229058
rect 146860 229002 146865 229058
rect 140832 229000 146865 229002
rect 41024 228998 41030 229000
rect 41775 228997 41841 229000
rect 146799 228997 146865 229000
rect 210159 228912 210225 228915
rect 674703 228912 674769 228915
rect 210159 228910 210528 228912
rect 210159 228854 210164 228910
rect 210220 228854 210528 228910
rect 210159 228852 210528 228854
rect 674703 228910 674814 228912
rect 674703 228854 674708 228910
rect 674764 228854 674814 228910
rect 210159 228849 210225 228852
rect 674703 228849 674814 228854
rect 674754 228660 674814 228849
rect 205167 228320 205233 228323
rect 205167 228318 210528 228320
rect 205167 228262 205172 228318
rect 205228 228262 210528 228318
rect 205167 228260 210528 228262
rect 205167 228257 205233 228260
rect 140802 227728 140862 227914
rect 674415 227876 674481 227879
rect 674415 227874 674784 227876
rect 674415 227818 674420 227874
rect 674476 227818 674784 227874
rect 674415 227816 674784 227818
rect 674415 227813 674481 227816
rect 146799 227728 146865 227731
rect 140802 227726 146865 227728
rect 140802 227670 146804 227726
rect 146860 227670 146865 227726
rect 140802 227668 146865 227670
rect 146799 227665 146865 227668
rect 204495 227728 204561 227731
rect 204495 227726 210528 227728
rect 204495 227670 204500 227726
rect 204556 227670 210528 227726
rect 204495 227668 210528 227670
rect 204495 227665 204561 227668
rect 673978 227370 673984 227434
rect 674048 227432 674054 227434
rect 674048 227372 674814 227432
rect 674048 227370 674054 227372
rect 41530 227222 41536 227286
rect 41600 227284 41606 227286
rect 41775 227284 41841 227287
rect 41600 227282 41841 227284
rect 41600 227226 41780 227282
rect 41836 227226 41841 227282
rect 41600 227224 41841 227226
rect 41600 227222 41606 227224
rect 41775 227221 41841 227224
rect 205647 227284 205713 227287
rect 205647 227282 210528 227284
rect 205647 227226 205652 227282
rect 205708 227226 210528 227282
rect 205647 227224 210528 227226
rect 205647 227221 205713 227224
rect 674754 227032 674814 227372
rect 40762 226630 40768 226694
rect 40832 226692 40838 226694
rect 41775 226692 41841 226695
rect 144015 226692 144081 226695
rect 40832 226690 41841 226692
rect 40832 226634 41780 226690
rect 41836 226634 41841 226690
rect 40832 226632 41841 226634
rect 140832 226690 144081 226692
rect 140832 226634 144020 226690
rect 144076 226634 144081 226690
rect 140832 226632 144081 226634
rect 40832 226630 40838 226632
rect 41775 226629 41841 226632
rect 144015 226629 144081 226632
rect 204879 226692 204945 226695
rect 204879 226690 210528 226692
rect 204879 226634 204884 226690
rect 204940 226634 210528 226690
rect 204879 226632 210528 226634
rect 204879 226629 204945 226632
rect 42063 226248 42129 226251
rect 42298 226248 42304 226250
rect 42063 226246 42304 226248
rect 42063 226190 42068 226246
rect 42124 226190 42304 226246
rect 42063 226188 42304 226190
rect 42063 226185 42129 226188
rect 42298 226186 42304 226188
rect 42368 226186 42374 226250
rect 673978 226186 673984 226250
rect 674048 226248 674054 226250
rect 674048 226188 674784 226248
rect 674048 226186 674054 226188
rect 205263 226100 205329 226103
rect 205263 226098 210528 226100
rect 205263 226042 205268 226098
rect 205324 226042 210528 226098
rect 205263 226040 210528 226042
rect 205263 226037 205329 226040
rect 674703 225804 674769 225807
rect 674703 225802 674814 225804
rect 674703 225746 674708 225802
rect 674764 225746 674814 225802
rect 674703 225741 674814 225746
rect 205455 225656 205521 225659
rect 205455 225654 210528 225656
rect 205455 225598 205460 225654
rect 205516 225598 210528 225654
rect 205455 225596 210528 225598
rect 205455 225593 205521 225596
rect 674754 225552 674814 225741
rect 140802 225064 140862 225466
rect 144015 225064 144081 225067
rect 140802 225062 144081 225064
rect 140802 225006 144020 225062
rect 144076 225006 144081 225062
rect 140802 225004 144081 225006
rect 144015 225001 144081 225004
rect 206991 225064 207057 225067
rect 206991 225062 210528 225064
rect 206991 225006 206996 225062
rect 207052 225006 210528 225062
rect 206991 225004 210528 225006
rect 206991 225001 207057 225004
rect 673839 224768 673905 224771
rect 673839 224766 674784 224768
rect 673839 224710 673844 224766
rect 673900 224710 674784 224766
rect 673839 224708 674784 224710
rect 673839 224705 673905 224708
rect 205743 224472 205809 224475
rect 205743 224470 210528 224472
rect 205743 224414 205748 224470
rect 205804 224414 210528 224470
rect 205743 224412 210528 224414
rect 205743 224409 205809 224412
rect 140802 223732 140862 224220
rect 204495 224028 204561 224031
rect 204495 224026 210528 224028
rect 204495 223970 204500 224026
rect 204556 223970 210528 224026
rect 204495 223968 210528 223970
rect 204495 223965 204561 223968
rect 673935 223880 674001 223883
rect 673935 223878 674784 223880
rect 673935 223822 673940 223878
rect 673996 223822 674784 223878
rect 673935 223820 674784 223822
rect 673935 223817 674001 223820
rect 144111 223732 144177 223735
rect 140802 223730 144177 223732
rect 140802 223674 144116 223730
rect 144172 223674 144177 223730
rect 140802 223672 144177 223674
rect 144111 223669 144177 223672
rect 205455 223436 205521 223439
rect 205455 223434 210528 223436
rect 205455 223378 205460 223434
rect 205516 223378 210528 223434
rect 205455 223376 210528 223378
rect 205455 223373 205521 223376
rect 210490 223078 210496 223142
rect 210560 223140 210566 223142
rect 211066 223140 211072 223142
rect 210560 223080 211072 223140
rect 210560 223078 210566 223080
rect 211066 223078 211072 223080
rect 211136 223078 211142 223142
rect 674362 223078 674368 223142
rect 674432 223140 674438 223142
rect 674432 223080 674784 223140
rect 674432 223078 674438 223080
rect 144015 222992 144081 222995
rect 140832 222990 144081 222992
rect 140832 222934 144020 222990
rect 144076 222934 144081 222990
rect 140832 222932 144081 222934
rect 144015 222929 144081 222932
rect 204591 222844 204657 222847
rect 204591 222842 210528 222844
rect 204591 222786 204596 222842
rect 204652 222786 210528 222842
rect 204591 222784 210528 222786
rect 204591 222781 204657 222784
rect 206895 222400 206961 222403
rect 206895 222398 210528 222400
rect 206895 222342 206900 222398
rect 206956 222342 210528 222398
rect 206895 222340 210528 222342
rect 206895 222337 206961 222340
rect 674415 222252 674481 222255
rect 674415 222250 674784 222252
rect 674415 222194 674420 222250
rect 674476 222194 674784 222250
rect 674415 222192 674784 222194
rect 674415 222189 674481 222192
rect 145594 221808 145600 221810
rect 140832 221748 145600 221808
rect 145594 221746 145600 221748
rect 145664 221746 145670 221810
rect 206415 221808 206481 221811
rect 206415 221806 210528 221808
rect 206415 221750 206420 221806
rect 206476 221750 210528 221806
rect 206415 221748 210528 221750
rect 206415 221745 206481 221748
rect 674946 221219 675006 221482
rect 204495 221216 204561 221219
rect 204495 221214 210528 221216
rect 204495 221158 204500 221214
rect 204556 221158 210528 221214
rect 204495 221156 210528 221158
rect 674946 221214 675057 221219
rect 674946 221158 674996 221214
rect 675052 221158 675057 221214
rect 674946 221156 675057 221158
rect 204495 221153 204561 221156
rect 674991 221153 675057 221156
rect 42351 221068 42417 221071
rect 42306 221066 42417 221068
rect 42306 221010 42356 221066
rect 42412 221010 42417 221066
rect 42306 221005 42417 221010
rect 204975 221068 205041 221071
rect 204975 221066 210558 221068
rect 204975 221010 204980 221066
rect 205036 221010 210558 221066
rect 204975 221008 210558 221010
rect 204975 221005 205041 221008
rect 42306 220890 42366 221005
rect 210498 220668 210558 221008
rect 42351 220328 42417 220331
rect 42306 220326 42417 220328
rect 42306 220270 42356 220326
rect 42412 220270 42417 220326
rect 42306 220265 42417 220270
rect 42306 220076 42366 220265
rect 140802 220180 140862 220668
rect 677058 220627 677118 220742
rect 677007 220622 677118 220627
rect 677007 220566 677012 220622
rect 677068 220566 677118 220622
rect 677007 220564 677118 220566
rect 677007 220561 677073 220564
rect 144015 220180 144081 220183
rect 140802 220178 144081 220180
rect 140802 220122 144020 220178
rect 144076 220122 144081 220178
rect 140802 220120 144081 220122
rect 144015 220117 144081 220120
rect 205359 220180 205425 220183
rect 205359 220178 210528 220180
rect 205359 220122 205364 220178
rect 205420 220122 210528 220178
rect 205359 220120 210528 220122
rect 205359 220117 205425 220120
rect 677058 219739 677118 220002
rect 677058 219734 677169 219739
rect 677058 219678 677108 219734
rect 677164 219678 677169 219734
rect 677058 219676 677169 219678
rect 677103 219673 677169 219676
rect 206895 219588 206961 219591
rect 206895 219586 210528 219588
rect 206895 219530 206900 219586
rect 206956 219530 210528 219586
rect 206895 219528 210528 219530
rect 206895 219525 206961 219528
rect 42351 219440 42417 219443
rect 42306 219438 42417 219440
rect 42306 219382 42356 219438
rect 42412 219382 42417 219438
rect 42306 219377 42417 219382
rect 42306 219262 42366 219377
rect 140802 218996 140862 219482
rect 204591 219440 204657 219443
rect 204591 219438 210558 219440
rect 204591 219382 204596 219438
rect 204652 219382 210558 219438
rect 204591 219380 210558 219382
rect 204591 219377 204657 219380
rect 210498 219040 210558 219380
rect 675138 218999 675198 219114
rect 145359 218996 145425 218999
rect 140802 218994 145425 218996
rect 140802 218938 145364 218994
rect 145420 218938 145425 218994
rect 140802 218936 145425 218938
rect 675138 218994 675249 218999
rect 675138 218938 675188 218994
rect 675244 218938 675249 218994
rect 675138 218936 675249 218938
rect 145359 218933 145425 218936
rect 675183 218933 675249 218936
rect 204495 218552 204561 218555
rect 204495 218550 210528 218552
rect 204495 218494 204500 218550
rect 204556 218494 210528 218550
rect 204495 218492 210528 218494
rect 204495 218489 204561 218492
rect 144015 218256 144081 218259
rect 140832 218254 144081 218256
rect 140832 218198 144020 218254
rect 144076 218198 144081 218254
rect 140832 218196 144081 218198
rect 144015 218193 144081 218196
rect 204591 217960 204657 217963
rect 204591 217958 210528 217960
rect 204591 217902 204596 217958
rect 204652 217902 210528 217958
rect 204591 217900 210528 217902
rect 204591 217897 204657 217900
rect 675138 217815 675198 218374
rect 204687 217812 204753 217815
rect 204687 217810 210558 217812
rect 204687 217754 204692 217810
rect 204748 217754 210558 217810
rect 204687 217752 210558 217754
rect 204687 217749 204753 217752
rect 43215 217664 43281 217667
rect 42336 217662 43281 217664
rect 42336 217606 43220 217662
rect 43276 217606 43281 217662
rect 42336 217604 43281 217606
rect 43215 217601 43281 217604
rect 210498 217412 210558 217752
rect 675087 217810 675198 217815
rect 675087 217754 675092 217810
rect 675148 217754 675198 217810
rect 675087 217752 675198 217754
rect 675087 217749 675153 217752
rect 674031 217516 674097 217519
rect 674031 217514 674784 217516
rect 674031 217458 674036 217514
rect 674092 217458 674784 217514
rect 674031 217456 674784 217458
rect 674031 217453 674097 217456
rect 43311 216924 43377 216927
rect 42336 216922 43377 216924
rect 42336 216866 43316 216922
rect 43372 216866 43377 216922
rect 42336 216864 43377 216866
rect 43311 216861 43377 216864
rect 140802 216480 140862 217034
rect 205359 216924 205425 216927
rect 205359 216922 210528 216924
rect 205359 216866 205364 216922
rect 205420 216866 210528 216922
rect 205359 216864 210528 216866
rect 205359 216861 205425 216864
rect 676866 216483 676926 216746
rect 145455 216480 145521 216483
rect 140802 216478 145521 216480
rect 140802 216422 145460 216478
rect 145516 216422 145521 216478
rect 140802 216420 145521 216422
rect 676866 216478 676977 216483
rect 676866 216422 676916 216478
rect 676972 216422 676977 216478
rect 676866 216420 676977 216422
rect 145455 216417 145521 216420
rect 676911 216417 676977 216420
rect 206703 216332 206769 216335
rect 206703 216330 210528 216332
rect 206703 216274 206708 216330
rect 206764 216274 210528 216330
rect 206703 216272 210528 216274
rect 206703 216269 206769 216272
rect 43407 216184 43473 216187
rect 42336 216182 43473 216184
rect 42336 216126 43412 216182
rect 43468 216126 43473 216182
rect 42336 216124 43473 216126
rect 43407 216121 43473 216124
rect 676866 215891 676926 216006
rect 204783 215888 204849 215891
rect 204783 215886 210558 215888
rect 204783 215830 204788 215886
rect 204844 215830 210558 215886
rect 204783 215828 210558 215830
rect 204783 215825 204849 215828
rect 210498 215784 210558 215828
rect 676815 215886 676926 215891
rect 676815 215830 676820 215886
rect 676876 215830 676926 215886
rect 676815 215828 676926 215830
rect 676815 215825 676881 215828
rect 140802 215296 140862 215784
rect 144111 215296 144177 215299
rect 140802 215294 144177 215296
rect 40386 214706 40446 215266
rect 140802 215238 144116 215294
rect 144172 215238 144177 215294
rect 140802 215236 144177 215238
rect 144111 215233 144177 215236
rect 204495 215296 204561 215299
rect 204495 215294 210528 215296
rect 204495 215238 204500 215294
rect 204556 215238 210528 215294
rect 204495 215236 210528 215238
rect 204495 215233 204561 215236
rect 674946 214707 675006 215192
rect 40378 214642 40384 214706
rect 40448 214642 40454 214706
rect 206127 214704 206193 214707
rect 206127 214702 210528 214704
rect 206127 214646 206132 214702
rect 206188 214646 210528 214702
rect 206127 214644 210528 214646
rect 674895 214702 675006 214707
rect 674895 214646 674900 214702
rect 674956 214646 675006 214702
rect 674895 214644 675006 214646
rect 206127 214641 206193 214644
rect 674895 214641 674961 214644
rect 144015 214556 144081 214559
rect 140832 214554 144081 214556
rect 41922 213967 41982 214526
rect 140832 214498 144020 214554
rect 144076 214498 144081 214554
rect 140832 214496 144081 214498
rect 144015 214493 144081 214496
rect 206319 214556 206385 214559
rect 206319 214554 210558 214556
rect 206319 214498 206324 214554
rect 206380 214498 210558 214554
rect 206319 214496 210558 214498
rect 206319 214493 206385 214496
rect 210498 214156 210558 214496
rect 674754 214263 674814 214378
rect 674754 214258 674865 214263
rect 674754 214202 674804 214258
rect 674860 214202 674865 214258
rect 674754 214200 674865 214202
rect 674799 214197 674865 214200
rect 41922 213962 42033 213967
rect 41922 213906 41972 213962
rect 42028 213906 42033 213962
rect 41922 213904 42033 213906
rect 41967 213901 42033 213904
rect 206511 213668 206577 213671
rect 206511 213666 210528 213668
rect 40578 213226 40638 213638
rect 206511 213610 206516 213666
rect 206572 213610 210528 213666
rect 206511 213608 210528 213610
rect 206511 213605 206577 213608
rect 674754 213375 674814 213564
rect 146415 213372 146481 213375
rect 140832 213370 146481 213372
rect 140832 213314 146420 213370
rect 146476 213314 146481 213370
rect 140832 213312 146481 213314
rect 146415 213309 146481 213312
rect 674703 213370 674814 213375
rect 674703 213314 674708 213370
rect 674764 213314 674814 213370
rect 674703 213312 674814 213314
rect 674703 213309 674769 213312
rect 40570 213162 40576 213226
rect 40640 213162 40646 213226
rect 206607 213076 206673 213079
rect 206607 213074 210528 213076
rect 206607 213018 206612 213074
rect 206668 213018 210528 213074
rect 206607 213016 210528 213018
rect 206607 213013 206673 213016
rect 204879 212928 204945 212931
rect 204879 212926 210558 212928
rect 40962 212486 41022 212898
rect 204879 212870 204884 212926
rect 204940 212870 210558 212926
rect 204879 212868 210558 212870
rect 204879 212865 204945 212868
rect 210498 212528 210558 212868
rect 40954 212422 40960 212486
rect 41024 212422 41030 212486
rect 41154 211598 41214 212158
rect 140802 211744 140862 212232
rect 679746 212191 679806 212750
rect 679746 212186 679857 212191
rect 679746 212130 679796 212186
rect 679852 212130 679857 212186
rect 679746 212128 679857 212130
rect 679791 212125 679857 212128
rect 206223 212040 206289 212043
rect 206223 212038 210528 212040
rect 206223 211982 206228 212038
rect 206284 211982 210528 212038
rect 206223 211980 210528 211982
rect 206223 211977 206289 211980
rect 145551 211744 145617 211747
rect 140802 211742 145617 211744
rect 140802 211686 145556 211742
rect 145612 211686 145617 211742
rect 140802 211684 145617 211686
rect 145551 211681 145617 211684
rect 41146 211534 41152 211598
rect 41216 211534 41222 211598
rect 206799 211448 206865 211451
rect 679791 211448 679857 211451
rect 206799 211446 210528 211448
rect 40194 210859 40254 211418
rect 206799 211390 206804 211446
rect 206860 211390 210528 211446
rect 206799 211388 210528 211390
rect 679746 211446 679857 211448
rect 679746 211390 679796 211446
rect 679852 211390 679857 211446
rect 206799 211385 206865 211388
rect 679746 211385 679857 211390
rect 679746 211270 679806 211385
rect 40194 210854 40305 210859
rect 40194 210798 40244 210854
rect 40300 210798 40305 210854
rect 40194 210796 40305 210798
rect 40239 210793 40305 210796
rect 140802 210560 140862 211048
rect 145743 210560 145809 210563
rect 140802 210558 145809 210560
rect 40770 210414 40830 210530
rect 140802 210502 145748 210558
rect 145804 210502 145809 210558
rect 140802 210500 145809 210502
rect 145743 210497 145809 210500
rect 40762 210350 40768 210414
rect 40832 210350 40838 210414
rect 640194 210412 640254 210826
rect 645615 210412 645681 210415
rect 647919 210412 647985 210415
rect 640194 210410 647985 210412
rect 640194 210354 645620 210410
rect 645676 210354 647924 210410
rect 647980 210354 647985 210410
rect 640194 210352 647985 210354
rect 645615 210349 645681 210352
rect 647919 210349 647985 210352
rect 204879 210264 204945 210267
rect 205071 210264 205137 210267
rect 207183 210266 207249 210267
rect 207183 210264 207232 210266
rect 204879 210262 205137 210264
rect 204879 210206 204884 210262
rect 204940 210206 205076 210262
rect 205132 210206 205137 210262
rect 204879 210204 205137 210206
rect 207140 210262 207232 210264
rect 207140 210206 207188 210262
rect 207140 210204 207232 210206
rect 204879 210201 204945 210204
rect 205071 210201 205137 210204
rect 207183 210202 207232 210204
rect 207296 210202 207302 210266
rect 676474 210202 676480 210266
rect 676544 210264 676550 210266
rect 680079 210264 680145 210267
rect 676544 210262 680145 210264
rect 676544 210206 680084 210262
rect 680140 210206 680145 210262
rect 676544 210204 680145 210206
rect 676544 210202 676550 210204
rect 207183 210201 207249 210202
rect 680079 210201 680145 210204
rect 676666 210054 676672 210118
rect 676736 210116 676742 210118
rect 679983 210116 680049 210119
rect 676736 210114 680049 210116
rect 676736 210058 679988 210114
rect 680044 210058 680049 210114
rect 676736 210056 680049 210058
rect 676736 210054 676742 210056
rect 679983 210053 680049 210056
rect 144111 209820 144177 209823
rect 140832 209818 144177 209820
rect 42114 209231 42174 209790
rect 140832 209762 144116 209818
rect 144172 209762 144177 209818
rect 140832 209760 144177 209762
rect 144111 209757 144177 209760
rect 42063 209226 42174 209231
rect 42063 209170 42068 209226
rect 42124 209170 42174 209226
rect 42063 209168 42174 209170
rect 42063 209165 42129 209168
rect 42831 208932 42897 208935
rect 42336 208930 42897 208932
rect 42336 208874 42836 208930
rect 42892 208874 42897 208930
rect 42336 208872 42897 208874
rect 42831 208869 42897 208872
rect 42306 207899 42366 208088
rect 140802 208044 140862 208602
rect 145647 208044 145713 208047
rect 140802 208042 145713 208044
rect 140802 207986 145652 208042
rect 145708 207986 145713 208042
rect 140802 207984 145713 207986
rect 145647 207981 145713 207984
rect 42306 207894 42417 207899
rect 42306 207838 42356 207894
rect 42412 207838 42417 207894
rect 42306 207836 42417 207838
rect 42351 207833 42417 207836
rect 675898 207686 675904 207750
rect 675968 207748 675974 207750
rect 677007 207748 677073 207751
rect 675968 207746 677073 207748
rect 675968 207690 677012 207746
rect 677068 207690 677073 207746
rect 675968 207688 677073 207690
rect 675968 207686 675974 207688
rect 677007 207685 677073 207688
rect 676282 207538 676288 207602
rect 676352 207600 676358 207602
rect 677103 207600 677169 207603
rect 676352 207598 677169 207600
rect 676352 207542 677108 207598
rect 677164 207542 677169 207598
rect 676352 207540 677169 207542
rect 676352 207538 676358 207540
rect 677103 207537 677169 207540
rect 144015 207452 144081 207455
rect 140832 207450 144081 207452
rect 40002 207159 40062 207422
rect 140832 207394 144020 207450
rect 144076 207394 144081 207450
rect 140832 207392 144081 207394
rect 144015 207389 144081 207392
rect 676090 207390 676096 207454
rect 676160 207452 676166 207454
rect 676911 207452 676977 207455
rect 676160 207450 676977 207452
rect 676160 207394 676916 207450
rect 676972 207394 676977 207450
rect 676160 207392 676977 207394
rect 676160 207390 676166 207392
rect 676911 207389 676977 207392
rect 40002 207154 40113 207159
rect 40002 207098 40052 207154
rect 40108 207098 40113 207154
rect 40002 207096 40113 207098
rect 40047 207093 40113 207096
rect 37314 206123 37374 206608
rect 37314 206118 37425 206123
rect 37314 206062 37364 206118
rect 37420 206062 37425 206118
rect 37314 206060 37425 206062
rect 37359 206057 37425 206060
rect 40194 205235 40254 205794
rect 140802 205676 140862 206154
rect 144015 205676 144081 205679
rect 140802 205674 144081 205676
rect 140802 205618 144020 205674
rect 144076 205618 144081 205674
rect 140802 205616 144081 205618
rect 144015 205613 144081 205616
rect 40143 205230 40254 205235
rect 40143 205174 40148 205230
rect 40204 205174 40254 205230
rect 40143 205172 40254 205174
rect 40143 205169 40209 205172
rect 145839 205084 145905 205087
rect 140832 205082 145905 205084
rect 140832 205026 145844 205082
rect 145900 205026 145905 205082
rect 140832 205024 145905 205026
rect 145839 205021 145905 205024
rect 42306 204936 42366 204980
rect 43119 204936 43185 204939
rect 42306 204934 43185 204936
rect 42306 204878 43124 204934
rect 43180 204878 43185 204934
rect 42306 204876 43185 204878
rect 43119 204873 43185 204876
rect 42351 204344 42417 204347
rect 42306 204342 42417 204344
rect 42306 204286 42356 204342
rect 42412 204286 42417 204342
rect 42306 204281 42417 204286
rect 42306 204166 42366 204281
rect 140802 203456 140862 203796
rect 144015 203456 144081 203459
rect 140802 203454 144081 203456
rect 140802 203398 144020 203454
rect 144076 203398 144081 203454
rect 140802 203396 144081 203398
rect 144015 203393 144081 203396
rect 42351 202864 42417 202867
rect 42306 202862 42417 202864
rect 42306 202806 42356 202862
rect 42412 202806 42417 202862
rect 42306 202801 42417 202806
rect 42306 202686 42366 202801
rect 205647 202716 205713 202719
rect 209295 202716 209361 202719
rect 205647 202714 210528 202716
rect 205647 202658 205652 202714
rect 205708 202658 209300 202714
rect 209356 202658 210528 202714
rect 205647 202656 210528 202658
rect 205647 202653 205713 202656
rect 209295 202653 209361 202656
rect 140802 202124 140862 202612
rect 144591 202124 144657 202127
rect 140802 202122 144657 202124
rect 140802 202066 144596 202122
rect 144652 202066 144657 202122
rect 140802 202064 144657 202066
rect 144591 202061 144657 202064
rect 144111 201384 144177 201387
rect 140832 201382 144177 201384
rect 140832 201326 144116 201382
rect 144172 201326 144177 201382
rect 140832 201324 144177 201326
rect 144111 201321 144177 201324
rect 210298 200582 210304 200646
rect 210368 200644 210374 200646
rect 211066 200644 211072 200646
rect 210368 200584 211072 200644
rect 210368 200582 210374 200584
rect 211066 200582 211072 200584
rect 211136 200582 211142 200646
rect 140802 199608 140862 200142
rect 146223 199608 146289 199611
rect 140802 199606 146289 199608
rect 140802 199550 146228 199606
rect 146284 199550 146289 199606
rect 140802 199548 146289 199550
rect 146223 199545 146289 199548
rect 675375 199314 675441 199315
rect 675322 199250 675328 199314
rect 675392 199312 675441 199314
rect 675392 199310 675484 199312
rect 675436 199254 675484 199310
rect 675392 199252 675484 199254
rect 675392 199250 675441 199252
rect 675375 199249 675441 199250
rect 144015 199016 144081 199019
rect 140832 199014 144081 199016
rect 140832 198958 144020 199014
rect 144076 198958 144081 199014
rect 140832 198956 144081 198958
rect 144015 198953 144081 198956
rect 210490 198954 210496 199018
rect 210560 198954 210566 199018
rect 210498 198868 210558 198954
rect 211066 198868 211072 198870
rect 210498 198808 211072 198868
rect 211066 198806 211072 198808
rect 211136 198806 211142 198870
rect 40911 198720 40977 198723
rect 675471 198722 675537 198723
rect 41338 198720 41344 198722
rect 40911 198718 41344 198720
rect 40911 198662 40916 198718
rect 40972 198662 41344 198718
rect 40911 198660 41344 198662
rect 40911 198657 40977 198660
rect 41338 198658 41344 198660
rect 41408 198658 41414 198722
rect 675471 198720 675520 198722
rect 675428 198718 675520 198720
rect 675428 198662 675476 198718
rect 675428 198660 675520 198662
rect 675471 198658 675520 198660
rect 675584 198658 675590 198722
rect 675471 198657 675537 198658
rect 675759 198424 675825 198427
rect 675898 198424 675904 198426
rect 675759 198422 675904 198424
rect 675759 198366 675764 198422
rect 675820 198366 675904 198422
rect 675759 198364 675904 198366
rect 675759 198361 675825 198364
rect 675898 198362 675904 198364
rect 675968 198362 675974 198426
rect 144015 197832 144081 197835
rect 140832 197830 144081 197832
rect 140832 197774 144020 197830
rect 144076 197774 144081 197830
rect 140832 197772 144081 197774
rect 144015 197769 144081 197772
rect 42159 197536 42225 197539
rect 42298 197536 42304 197538
rect 42159 197534 42304 197536
rect 42159 197478 42164 197534
rect 42220 197478 42304 197534
rect 42159 197476 42304 197478
rect 42159 197473 42225 197476
rect 42298 197474 42304 197476
rect 42368 197474 42374 197538
rect 144399 196648 144465 196651
rect 140832 196646 144465 196648
rect 140832 196590 144404 196646
rect 144460 196590 144465 196646
rect 140832 196588 144465 196590
rect 144399 196585 144465 196588
rect 42351 195170 42417 195171
rect 42298 195168 42304 195170
rect 42260 195108 42304 195168
rect 42368 195166 42417 195170
rect 42412 195110 42417 195166
rect 42298 195106 42304 195108
rect 42368 195106 42417 195110
rect 42351 195105 42417 195106
rect 140802 194872 140862 195360
rect 675759 195316 675825 195319
rect 676090 195316 676096 195318
rect 675759 195314 676096 195316
rect 675759 195258 675764 195314
rect 675820 195258 676096 195314
rect 675759 195256 676096 195258
rect 675759 195253 675825 195256
rect 676090 195254 676096 195256
rect 676160 195254 676166 195318
rect 144303 194872 144369 194875
rect 140802 194870 144369 194872
rect 140802 194814 144308 194870
rect 144364 194814 144369 194870
rect 140802 194812 144369 194814
rect 144303 194809 144369 194812
rect 140802 193688 140862 194176
rect 145935 193688 146001 193691
rect 140802 193686 146001 193688
rect 140802 193630 145940 193686
rect 145996 193630 146001 193686
rect 140802 193628 146001 193630
rect 145935 193625 146001 193628
rect 674362 193478 674368 193542
rect 674432 193540 674438 193542
rect 675375 193540 675441 193543
rect 674432 193538 675441 193540
rect 674432 193482 675380 193538
rect 675436 193482 675441 193538
rect 674432 193480 675441 193482
rect 674432 193478 674438 193480
rect 675375 193477 675441 193480
rect 144015 192948 144081 192951
rect 140832 192946 144081 192948
rect 140832 192890 144020 192946
rect 144076 192890 144081 192946
rect 140832 192888 144081 192890
rect 144015 192885 144081 192888
rect 146031 191764 146097 191767
rect 140832 191762 146097 191764
rect 140832 191706 146036 191762
rect 146092 191706 146097 191762
rect 140832 191704 146097 191706
rect 146031 191701 146097 191704
rect 675759 191616 675825 191619
rect 676282 191616 676288 191618
rect 675759 191614 676288 191616
rect 675759 191558 675764 191614
rect 675820 191558 676288 191614
rect 675759 191556 676288 191558
rect 675759 191553 675825 191556
rect 676282 191554 676288 191556
rect 676352 191554 676358 191618
rect 41338 190962 41344 191026
rect 41408 191024 41414 191026
rect 41775 191024 41841 191027
rect 41408 191022 41841 191024
rect 41408 190966 41780 191022
rect 41836 190966 41841 191022
rect 41408 190964 41841 190966
rect 41408 190962 41414 190964
rect 41775 190961 41841 190964
rect 41146 190074 41152 190138
rect 41216 190136 41222 190138
rect 41775 190136 41841 190139
rect 41216 190134 41841 190136
rect 41216 190078 41780 190134
rect 41836 190078 41841 190134
rect 41216 190076 41841 190078
rect 140802 190136 140862 190476
rect 146223 190136 146289 190139
rect 207279 190138 207345 190139
rect 207226 190136 207232 190138
rect 140802 190134 146289 190136
rect 140802 190078 146228 190134
rect 146284 190078 146289 190134
rect 140802 190076 146289 190078
rect 207188 190076 207232 190136
rect 207296 190134 207345 190138
rect 207340 190078 207345 190134
rect 41216 190074 41222 190076
rect 41775 190073 41841 190076
rect 146223 190073 146289 190076
rect 207226 190074 207232 190076
rect 207296 190074 207345 190078
rect 207279 190073 207345 190074
rect 146127 189396 146193 189399
rect 140832 189394 146193 189396
rect 140832 189338 146132 189394
rect 146188 189338 146193 189394
rect 140832 189336 146193 189338
rect 146127 189333 146193 189336
rect 41967 189102 42033 189103
rect 41914 189100 41920 189102
rect 41876 189040 41920 189100
rect 41984 189098 42033 189102
rect 42028 189042 42033 189098
rect 41914 189038 41920 189040
rect 41984 189038 42033 189042
rect 41967 189037 42033 189038
rect 41775 188362 41841 188363
rect 41722 188298 41728 188362
rect 41792 188360 41841 188362
rect 41792 188358 41884 188360
rect 41836 188302 41884 188358
rect 41792 188300 41884 188302
rect 41792 188298 41841 188300
rect 41775 188297 41841 188298
rect 146415 188212 146481 188215
rect 140832 188210 146481 188212
rect 140832 188154 146420 188210
rect 146476 188154 146481 188210
rect 140832 188152 146481 188154
rect 146415 188149 146481 188152
rect 140802 186436 140862 186924
rect 146415 186436 146481 186439
rect 140802 186434 146481 186436
rect 140802 186378 146420 186434
rect 146476 186378 146481 186434
rect 140802 186376 146481 186378
rect 146415 186373 146481 186376
rect 40954 185930 40960 185994
rect 41024 185992 41030 185994
rect 41775 185992 41841 185995
rect 41024 185990 41841 185992
rect 41024 185934 41780 185990
rect 41836 185934 41841 185990
rect 41024 185932 41841 185934
rect 41024 185930 41030 185932
rect 41775 185929 41841 185932
rect 140802 185252 140862 185740
rect 144495 185252 144561 185255
rect 140802 185250 144561 185252
rect 140802 185194 144500 185250
rect 144556 185194 144561 185250
rect 140802 185192 144561 185194
rect 144495 185189 144561 185192
rect 146799 184512 146865 184515
rect 140832 184510 146865 184512
rect 140832 184454 146804 184510
rect 146860 184454 146865 184510
rect 140832 184452 146865 184454
rect 146799 184449 146865 184452
rect 674415 184512 674481 184515
rect 674415 184510 674784 184512
rect 674415 184454 674420 184510
rect 674476 184454 674784 184510
rect 674415 184452 674784 184454
rect 674415 184449 674481 184452
rect 40378 184154 40384 184218
rect 40448 184216 40454 184218
rect 41775 184216 41841 184219
rect 40448 184214 41841 184216
rect 40448 184158 41780 184214
rect 41836 184158 41841 184214
rect 40448 184156 41841 184158
rect 40448 184154 40454 184156
rect 41775 184153 41841 184156
rect 674703 183920 674769 183923
rect 674703 183918 674814 183920
rect 674703 183862 674708 183918
rect 674764 183862 674814 183918
rect 674703 183857 674814 183862
rect 674754 183668 674814 183857
rect 40762 183562 40768 183626
rect 40832 183624 40838 183626
rect 41775 183624 41841 183627
rect 40832 183622 41841 183624
rect 40832 183566 41780 183622
rect 41836 183566 41841 183622
rect 40832 183564 41841 183566
rect 40832 183562 40838 183564
rect 41775 183561 41841 183564
rect 146607 183328 146673 183331
rect 140832 183326 146673 183328
rect 140832 183270 146612 183326
rect 146668 183270 146673 183326
rect 140832 183268 146673 183270
rect 146607 183265 146673 183268
rect 40570 182822 40576 182886
rect 40640 182884 40646 182886
rect 41775 182884 41841 182887
rect 40640 182882 41841 182884
rect 40640 182826 41780 182882
rect 41836 182826 41841 182882
rect 40640 182824 41841 182826
rect 40640 182822 40646 182824
rect 41775 182821 41841 182824
rect 674415 182884 674481 182887
rect 674415 182882 674784 182884
rect 674415 182826 674420 182882
rect 674476 182826 674784 182882
rect 674415 182824 674784 182826
rect 674415 182821 674481 182824
rect 673978 182526 673984 182590
rect 674048 182588 674054 182590
rect 674048 182528 674814 182588
rect 674048 182526 674054 182528
rect 140802 181848 140862 182188
rect 674754 182040 674814 182528
rect 146799 181848 146865 181851
rect 140802 181846 146865 181848
rect 140802 181790 146804 181846
rect 146860 181790 146865 181846
rect 140802 181788 146865 181790
rect 146799 181785 146865 181788
rect 673978 181194 673984 181258
rect 674048 181256 674054 181258
rect 674048 181196 674784 181256
rect 674048 181194 674054 181196
rect 140802 180516 140862 180994
rect 676474 180898 676480 180962
rect 676544 180898 676550 180962
rect 144687 180516 144753 180519
rect 140802 180514 144753 180516
rect 140802 180458 144692 180514
rect 144748 180458 144753 180514
rect 140802 180456 144753 180458
rect 144687 180453 144753 180456
rect 676482 179924 676542 180898
rect 679695 179924 679761 179927
rect 676482 179922 679761 179924
rect 676482 179866 679700 179922
rect 679756 179866 679761 179922
rect 676482 179864 679761 179866
rect 679695 179861 679761 179864
rect 145263 179776 145329 179779
rect 140832 179774 145329 179776
rect 140832 179718 145268 179774
rect 145324 179718 145329 179774
rect 140832 179716 145329 179718
rect 145263 179713 145329 179716
rect 676674 179482 676734 179746
rect 676666 179418 676672 179482
rect 676736 179480 676742 179482
rect 679791 179480 679857 179483
rect 676736 179478 679857 179480
rect 676736 179422 679796 179478
rect 679852 179422 679857 179478
rect 676736 179420 679857 179422
rect 676736 179418 676742 179420
rect 679791 179417 679857 179420
rect 146799 178592 146865 178595
rect 674754 178594 674814 178858
rect 140832 178590 146865 178592
rect 140832 178534 146804 178590
rect 146860 178534 146865 178590
rect 140832 178532 146865 178534
rect 146799 178529 146865 178532
rect 674746 178530 674752 178594
rect 674816 178530 674822 178594
rect 674170 178086 674176 178150
rect 674240 178148 674246 178150
rect 674240 178088 674784 178148
rect 674240 178086 674246 178088
rect 140802 176816 140862 177304
rect 674946 177115 675006 177230
rect 674895 177110 675006 177115
rect 674895 177054 674900 177110
rect 674956 177054 675006 177110
rect 674895 177052 675006 177054
rect 674895 177049 674961 177052
rect 146799 176816 146865 176819
rect 140802 176814 146865 176816
rect 140802 176758 146804 176814
rect 146860 176758 146865 176814
rect 140802 176756 146865 176758
rect 146799 176753 146865 176756
rect 677058 176227 677118 176490
rect 677007 176222 677118 176227
rect 677007 176166 677012 176222
rect 677068 176166 677118 176222
rect 677007 176164 677118 176166
rect 677007 176161 677073 176164
rect 145263 176076 145329 176079
rect 140832 176074 145329 176076
rect 140832 176018 145268 176074
rect 145324 176018 145329 176074
rect 140832 176016 145329 176018
rect 145263 176013 145329 176016
rect 676911 175632 676977 175635
rect 677058 175632 677118 175750
rect 676911 175630 677118 175632
rect 676911 175574 676916 175630
rect 676972 175574 677118 175630
rect 676911 175572 677118 175574
rect 676911 175569 676977 175572
rect 140802 174448 140862 174982
rect 677250 174747 677310 175010
rect 677199 174742 677310 174747
rect 677199 174686 677204 174742
rect 677260 174686 677310 174742
rect 677199 174684 677310 174686
rect 677199 174681 677265 174684
rect 145167 174448 145233 174451
rect 140802 174446 145233 174448
rect 140802 174390 145172 174446
rect 145228 174390 145233 174446
rect 140802 174388 145233 174390
rect 145167 174385 145233 174388
rect 674946 174007 675006 174122
rect 674946 174002 675057 174007
rect 674946 173946 674996 174002
rect 675052 173946 675057 174002
rect 674946 173944 675057 173946
rect 674991 173941 675057 173944
rect 140802 173412 140862 173752
rect 146799 173412 146865 173415
rect 140802 173410 146865 173412
rect 140802 173354 146804 173410
rect 146860 173354 146865 173410
rect 140802 173352 146865 173354
rect 146799 173349 146865 173352
rect 674754 173119 674814 173382
rect 674754 173114 674865 173119
rect 674754 173058 674804 173114
rect 674860 173058 674865 173114
rect 674754 173056 674865 173058
rect 674799 173053 674865 173056
rect 211066 172758 211072 172822
rect 211136 172758 211142 172822
rect 210159 172672 210225 172675
rect 210874 172672 210880 172674
rect 210159 172670 210880 172672
rect 210159 172614 210164 172670
rect 210220 172614 210880 172670
rect 210159 172612 210880 172614
rect 210159 172609 210225 172612
rect 210874 172610 210880 172612
rect 210944 172610 210950 172674
rect 140802 172080 140862 172562
rect 210298 172462 210304 172526
rect 210368 172524 210374 172526
rect 211074 172524 211134 172758
rect 210368 172464 211134 172524
rect 210368 172462 210374 172464
rect 674511 172376 674577 172379
rect 674754 172376 674814 172494
rect 674511 172374 674814 172376
rect 674511 172318 674516 172374
rect 674572 172318 674814 172374
rect 674511 172316 674814 172318
rect 674511 172313 674577 172316
rect 144879 172080 144945 172083
rect 140802 172078 144945 172080
rect 140802 172022 144884 172078
rect 144940 172022 144945 172078
rect 140802 172020 144945 172022
rect 144879 172017 144945 172020
rect 677058 171491 677118 171754
rect 677058 171486 677169 171491
rect 677058 171430 677108 171486
rect 677164 171430 677169 171486
rect 677058 171428 677169 171430
rect 677103 171425 677169 171428
rect 146799 171340 146865 171343
rect 140832 171338 146865 171340
rect 140832 171282 146804 171338
rect 146860 171282 146865 171338
rect 140832 171280 146865 171282
rect 146799 171277 146865 171280
rect 676866 170899 676926 171014
rect 676815 170894 676926 170899
rect 676815 170838 676820 170894
rect 676876 170838 676926 170894
rect 676815 170836 676926 170838
rect 676815 170833 676881 170836
rect 145071 170156 145137 170159
rect 140832 170154 145137 170156
rect 140832 170098 145076 170154
rect 145132 170098 145137 170154
rect 140832 170096 145137 170098
rect 145071 170093 145137 170096
rect 675138 170011 675198 170200
rect 675087 170006 675198 170011
rect 675087 169950 675092 170006
rect 675148 169950 675198 170006
rect 675087 169948 675198 169950
rect 675087 169945 675153 169948
rect 674223 169416 674289 169419
rect 674223 169414 674784 169416
rect 674223 169358 674228 169414
rect 674284 169358 674784 169414
rect 674223 169356 674784 169358
rect 674223 169353 674289 169356
rect 140802 168380 140862 168868
rect 674127 168528 674193 168531
rect 674754 168528 674814 168572
rect 674127 168526 674814 168528
rect 674127 168470 674132 168526
rect 674188 168470 674814 168526
rect 674127 168468 674814 168470
rect 674127 168465 674193 168468
rect 144975 168380 145041 168383
rect 140802 168378 145041 168380
rect 140802 168322 144980 168378
rect 145036 168322 145041 168378
rect 140802 168320 145041 168322
rect 144975 168317 145041 168320
rect 146799 167640 146865 167643
rect 140832 167638 146865 167640
rect 140832 167582 146804 167638
rect 146860 167582 146865 167638
rect 140832 167580 146865 167582
rect 146799 167577 146865 167580
rect 674754 167347 674814 167758
rect 674703 167342 674814 167347
rect 674703 167286 674708 167342
rect 674764 167286 674814 167342
rect 674703 167284 674814 167286
rect 674703 167281 674769 167284
rect 144015 166604 144081 166607
rect 140832 166602 144081 166604
rect 140832 166546 144020 166602
rect 144076 166546 144081 166602
rect 140832 166544 144081 166546
rect 640386 166604 640446 166870
rect 646287 166604 646353 166607
rect 640386 166602 646353 166604
rect 640386 166546 646292 166602
rect 646348 166546 646353 166602
rect 640386 166544 646353 166546
rect 144015 166541 144081 166544
rect 646287 166541 646353 166544
rect 674607 166604 674673 166607
rect 674754 166604 674814 166944
rect 679695 166604 679761 166607
rect 674607 166602 674814 166604
rect 674607 166546 674612 166602
rect 674668 166546 674814 166602
rect 674607 166544 674814 166546
rect 674946 166602 679761 166604
rect 674946 166546 679700 166602
rect 679756 166546 679761 166602
rect 674946 166544 679761 166546
rect 674607 166541 674673 166544
rect 674554 166394 674560 166458
rect 674624 166456 674630 166458
rect 674946 166456 675006 166544
rect 679695 166541 679761 166544
rect 674624 166396 675006 166456
rect 675759 166456 675825 166459
rect 679791 166456 679857 166459
rect 675759 166454 679857 166456
rect 675759 166398 675764 166454
rect 675820 166398 679796 166454
rect 679852 166398 679857 166454
rect 675759 166396 679857 166398
rect 674624 166394 674630 166396
rect 675759 166393 675825 166396
rect 679791 166393 679857 166396
rect 647919 166308 647985 166311
rect 640416 166306 647985 166308
rect 640416 166250 647924 166306
rect 647980 166250 647985 166306
rect 640416 166248 647985 166250
rect 647919 166245 647985 166248
rect 647055 166012 647121 166015
rect 640386 166010 647121 166012
rect 640386 165954 647060 166010
rect 647116 165954 647121 166010
rect 640386 165952 647121 165954
rect 640386 165686 640446 165952
rect 647055 165949 647121 165952
rect 674754 165719 674814 166278
rect 674703 165714 674814 165719
rect 674703 165658 674708 165714
rect 674764 165658 674814 165714
rect 674703 165656 674814 165658
rect 674703 165653 674769 165656
rect 674362 165506 674368 165570
rect 674432 165568 674438 165570
rect 675759 165568 675825 165571
rect 674432 165566 675825 165568
rect 674432 165510 675764 165566
rect 675820 165510 675825 165566
rect 674432 165508 675825 165510
rect 674432 165506 674438 165508
rect 675759 165505 675825 165508
rect 140802 164828 140862 165316
rect 144495 164828 144561 164831
rect 140802 164826 144561 164828
rect 140802 164770 144500 164826
rect 144556 164770 144561 164826
rect 140802 164768 144561 164770
rect 144495 164765 144561 164768
rect 140802 163644 140862 164130
rect 676666 164026 676672 164090
rect 676736 164088 676742 164090
rect 677199 164088 677265 164091
rect 676736 164086 677265 164088
rect 676736 164030 677204 164086
rect 677260 164030 677265 164086
rect 676736 164028 677265 164030
rect 676736 164026 676742 164028
rect 677199 164025 677265 164028
rect 144687 163644 144753 163647
rect 140802 163642 144753 163644
rect 140802 163586 144692 163642
rect 144748 163586 144753 163642
rect 140802 163584 144753 163586
rect 144687 163581 144753 163584
rect 144015 162904 144081 162907
rect 140832 162902 144081 162904
rect 140832 162846 144020 162902
rect 144076 162846 144081 162902
rect 140832 162844 144081 162846
rect 144015 162841 144081 162844
rect 676474 162842 676480 162906
rect 676544 162904 676550 162906
rect 676911 162904 676977 162907
rect 676544 162902 676977 162904
rect 676544 162846 676916 162902
rect 676972 162846 676977 162902
rect 676544 162844 676977 162846
rect 676544 162842 676550 162844
rect 676911 162841 676977 162844
rect 140802 161424 140862 161682
rect 144783 161424 144849 161427
rect 140802 161422 144849 161424
rect 140802 161366 144788 161422
rect 144844 161366 144849 161422
rect 140802 161364 144849 161366
rect 144783 161361 144849 161364
rect 675898 161362 675904 161426
rect 675968 161424 675974 161426
rect 677007 161424 677073 161427
rect 675968 161422 677073 161424
rect 675968 161366 677012 161422
rect 677068 161366 677073 161422
rect 675968 161364 677073 161366
rect 675968 161362 675974 161364
rect 677007 161361 677073 161364
rect 140802 159944 140862 160432
rect 144111 159944 144177 159947
rect 140802 159942 144177 159944
rect 140802 159886 144116 159942
rect 144172 159886 144177 159942
rect 140802 159884 144177 159886
rect 144111 159881 144177 159884
rect 144015 159352 144081 159355
rect 140832 159350 144081 159352
rect 140832 159294 144020 159350
rect 144076 159294 144081 159350
rect 140832 159292 144081 159294
rect 144015 159289 144081 159292
rect 674746 159290 674752 159354
rect 674816 159352 674822 159354
rect 675375 159352 675441 159355
rect 674816 159350 675441 159352
rect 674816 159294 675380 159350
rect 675436 159294 675441 159350
rect 674816 159292 675441 159294
rect 674816 159290 674822 159292
rect 675375 159289 675441 159292
rect 144207 158168 144273 158171
rect 140832 158166 144273 158168
rect 140832 158110 144212 158166
rect 144268 158110 144273 158166
rect 140832 158108 144273 158110
rect 144207 158105 144273 158108
rect 675759 157724 675825 157727
rect 675898 157724 675904 157726
rect 675759 157722 675904 157724
rect 675759 157666 675764 157722
rect 675820 157666 675904 157722
rect 675759 157664 675904 157666
rect 675759 157661 675825 157664
rect 675898 157662 675904 157664
rect 675968 157662 675974 157726
rect 140802 156392 140862 156880
rect 144111 156392 144177 156395
rect 140802 156390 144177 156392
rect 140802 156334 144116 156390
rect 144172 156334 144177 156390
rect 140802 156332 144177 156334
rect 144111 156329 144177 156332
rect 144015 155800 144081 155803
rect 140802 155798 144081 155800
rect 140802 155742 144020 155798
rect 144076 155742 144081 155798
rect 140802 155740 144081 155742
rect 140802 155698 140862 155740
rect 144015 155737 144081 155740
rect 675375 154618 675441 154619
rect 675322 154554 675328 154618
rect 675392 154616 675441 154618
rect 675392 154614 675484 154616
rect 675436 154558 675484 154614
rect 675392 154556 675484 154558
rect 675392 154554 675441 154556
rect 675375 154553 675441 154554
rect 144111 154468 144177 154471
rect 140832 154466 144177 154468
rect 140832 154410 144116 154466
rect 144172 154410 144177 154466
rect 140832 154408 144177 154410
rect 144111 154405 144177 154408
rect 675375 154320 675441 154323
rect 675514 154320 675520 154322
rect 675375 154318 675520 154320
rect 675375 154262 675380 154318
rect 675436 154262 675520 154318
rect 675375 154260 675520 154262
rect 675375 154257 675441 154260
rect 675514 154258 675520 154260
rect 675584 154258 675590 154322
rect 675759 153432 675825 153435
rect 676474 153432 676480 153434
rect 675759 153430 676480 153432
rect 675759 153374 675764 153430
rect 675820 153374 676480 153430
rect 675759 153372 676480 153374
rect 675759 153369 675825 153372
rect 676474 153370 676480 153372
rect 676544 153370 676550 153434
rect 140802 152988 140862 153250
rect 144015 152988 144081 152991
rect 140802 152986 144081 152988
rect 140802 152930 144020 152986
rect 144076 152930 144081 152986
rect 140802 152928 144081 152930
rect 144015 152925 144081 152928
rect 210682 152778 210688 152842
rect 210752 152840 210758 152842
rect 210752 152780 210942 152840
rect 210752 152778 210758 152780
rect 210159 152692 210225 152695
rect 210682 152692 210688 152694
rect 210159 152690 210688 152692
rect 210159 152634 210164 152690
rect 210220 152634 210688 152690
rect 210159 152632 210688 152634
rect 210159 152629 210225 152632
rect 210682 152630 210688 152632
rect 210752 152630 210758 152694
rect 210882 152692 210942 152780
rect 211066 152692 211072 152694
rect 210882 152632 211072 152692
rect 211066 152630 211072 152632
rect 211136 152630 211142 152694
rect 140802 151656 140862 152144
rect 144111 151656 144177 151659
rect 140802 151654 144177 151656
rect 140802 151598 144116 151654
rect 144172 151598 144177 151654
rect 140802 151596 144177 151598
rect 144111 151593 144177 151596
rect 210298 151594 210304 151658
rect 210368 151656 210374 151658
rect 211066 151656 211072 151658
rect 210368 151596 211072 151656
rect 210368 151594 210374 151596
rect 211066 151594 211072 151596
rect 211136 151594 211142 151658
rect 144015 150916 144081 150919
rect 140832 150914 144081 150916
rect 140832 150858 144020 150914
rect 144076 150858 144081 150914
rect 140832 150856 144081 150858
rect 144015 150853 144081 150856
rect 149103 149732 149169 149735
rect 140832 149730 149169 149732
rect 140832 149674 149108 149730
rect 149164 149674 149169 149730
rect 140832 149672 149169 149674
rect 149103 149669 149169 149672
rect 674170 148486 674176 148550
rect 674240 148548 674246 148550
rect 675471 148548 675537 148551
rect 674240 148546 675537 148548
rect 674240 148490 675476 148546
rect 675532 148490 675537 148546
rect 674240 148488 675537 148490
rect 674240 148486 674246 148488
rect 675471 148485 675537 148488
rect 140802 147956 140862 148444
rect 674746 148338 674752 148402
rect 674816 148400 674822 148402
rect 675183 148400 675249 148403
rect 674816 148398 675249 148400
rect 674816 148342 675188 148398
rect 675244 148342 675249 148398
rect 674816 148340 675249 148342
rect 674816 148338 674822 148340
rect 675183 148337 675249 148340
rect 144495 147956 144561 147959
rect 140802 147954 144561 147956
rect 140802 147898 144500 147954
rect 144556 147898 144561 147954
rect 140802 147896 144561 147898
rect 144495 147893 144561 147896
rect 140802 147068 140862 147260
rect 144207 147068 144273 147071
rect 140802 147066 144273 147068
rect 140802 147010 144212 147066
rect 144268 147010 144273 147066
rect 140802 147008 144273 147010
rect 144207 147005 144273 147008
rect 675759 146624 675825 146627
rect 676666 146624 676672 146626
rect 675759 146622 676672 146624
rect 675759 146566 675764 146622
rect 675820 146566 676672 146622
rect 675759 146564 676672 146566
rect 675759 146561 675825 146564
rect 676666 146562 676672 146564
rect 676736 146562 676742 146626
rect 144207 146032 144273 146035
rect 140832 146030 144273 146032
rect 140832 145974 144212 146030
rect 144268 145974 144273 146030
rect 140832 145972 144273 145974
rect 144207 145969 144273 145972
rect 140802 144256 140862 144790
rect 144207 144256 144273 144259
rect 140802 144254 144273 144256
rect 140802 144198 144212 144254
rect 144268 144198 144273 144254
rect 140802 144196 144273 144198
rect 144207 144193 144273 144196
rect 140802 143220 140862 143708
rect 144207 143220 144273 143223
rect 140802 143218 144273 143220
rect 140802 143162 144212 143218
rect 144268 143162 144273 143218
rect 140802 143160 144273 143162
rect 144207 143157 144273 143160
rect 144207 142480 144273 142483
rect 140832 142478 144273 142480
rect 140832 142422 144212 142478
rect 144268 142422 144273 142478
rect 140832 142420 144273 142422
rect 144207 142417 144273 142420
rect 143919 141296 143985 141299
rect 140832 141294 143985 141296
rect 140832 141238 143924 141294
rect 143980 141238 143985 141294
rect 140832 141236 143985 141238
rect 143919 141233 143985 141236
rect 140802 139520 140862 140008
rect 144495 139520 144561 139523
rect 140802 139518 144561 139520
rect 140802 139462 144500 139518
rect 144556 139462 144561 139518
rect 140802 139460 144561 139462
rect 144495 139457 144561 139460
rect 674754 139079 674814 139342
rect 674703 139074 674814 139079
rect 674703 139018 674708 139074
rect 674764 139018 674814 139074
rect 674703 139016 674814 139018
rect 674703 139013 674769 139016
rect 140802 138336 140862 138824
rect 674415 138484 674481 138487
rect 674415 138482 674784 138484
rect 674415 138426 674420 138482
rect 674476 138426 674784 138482
rect 674415 138424 674784 138426
rect 674415 138421 674481 138424
rect 143823 138336 143889 138339
rect 140802 138334 143889 138336
rect 140802 138278 143828 138334
rect 143884 138278 143889 138334
rect 140802 138276 143889 138278
rect 143823 138273 143889 138276
rect 146895 137596 146961 137599
rect 140832 137594 146961 137596
rect 140832 137538 146900 137594
rect 146956 137538 146961 137594
rect 140832 137536 146961 137538
rect 146895 137533 146961 137536
rect 674607 137300 674673 137303
rect 674754 137300 674814 137640
rect 674607 137298 674814 137300
rect 674607 137242 674612 137298
rect 674668 137242 674814 137298
rect 674607 137240 674814 137242
rect 674607 137237 674673 137240
rect 673978 136794 673984 136858
rect 674048 136856 674054 136858
rect 674048 136796 674784 136856
rect 674048 136794 674054 136796
rect 140802 136116 140862 136522
rect 146895 136116 146961 136119
rect 140802 136114 146961 136116
rect 140802 136058 146900 136114
rect 146956 136058 146961 136114
rect 140802 136056 146961 136058
rect 146895 136053 146961 136056
rect 674754 135675 674814 136012
rect 674703 135670 674814 135675
rect 674703 135614 674708 135670
rect 674764 135614 674814 135670
rect 674703 135612 674814 135614
rect 674703 135609 674769 135612
rect 674554 135462 674560 135526
rect 674624 135462 674630 135526
rect 674562 135376 674622 135462
rect 674562 135316 674784 135376
rect 140802 134784 140862 135272
rect 673551 134932 673617 134935
rect 674554 134932 674560 134934
rect 673551 134930 674560 134932
rect 673551 134874 673556 134930
rect 673612 134874 674560 134930
rect 673551 134872 674560 134874
rect 673551 134869 673617 134872
rect 674554 134870 674560 134872
rect 674624 134870 674630 134934
rect 144207 134784 144273 134787
rect 140802 134782 144273 134784
rect 140802 134726 144212 134782
rect 144268 134726 144273 134782
rect 140802 134724 144273 134726
rect 144207 134721 144273 134724
rect 674362 134500 674368 134564
rect 674432 134562 674438 134564
rect 674432 134502 674784 134562
rect 674432 134500 674438 134502
rect 146799 134490 146865 134491
rect 146746 134488 146752 134490
rect 146708 134428 146752 134488
rect 146816 134486 146865 134490
rect 146860 134430 146865 134486
rect 146746 134426 146752 134428
rect 146816 134426 146865 134430
rect 146799 134425 146865 134426
rect 144207 134044 144273 134047
rect 140832 134042 144273 134044
rect 140832 133986 144212 134042
rect 144268 133986 144273 134042
rect 140832 133984 144273 133986
rect 144207 133981 144273 133984
rect 674170 133686 674176 133750
rect 674240 133748 674246 133750
rect 674240 133688 674784 133748
rect 674240 133686 674246 133688
rect 144495 132860 144561 132863
rect 140832 132858 144561 132860
rect 140832 132802 144500 132858
rect 144556 132802 144561 132858
rect 140832 132800 144561 132802
rect 144495 132797 144561 132800
rect 210490 132650 210496 132714
rect 210560 132712 210566 132714
rect 211066 132712 211072 132714
rect 210560 132652 211072 132712
rect 210560 132650 210566 132652
rect 211066 132650 211072 132652
rect 211136 132650 211142 132714
rect 146799 132566 146865 132567
rect 674946 132566 675006 132904
rect 146746 132564 146752 132566
rect 146708 132504 146752 132564
rect 146816 132562 146865 132566
rect 146860 132506 146865 132562
rect 146746 132502 146752 132504
rect 146816 132502 146865 132506
rect 674938 132502 674944 132566
rect 675008 132502 675014 132566
rect 146799 132501 146865 132502
rect 675522 131827 675582 132090
rect 675471 131822 675582 131827
rect 675471 131766 675476 131822
rect 675532 131766 675582 131822
rect 675471 131764 675582 131766
rect 675471 131761 675537 131764
rect 140802 131084 140862 131572
rect 675138 131087 675198 131202
rect 144495 131084 144561 131087
rect 140802 131082 144561 131084
rect 140802 131026 144500 131082
rect 144556 131026 144561 131082
rect 140802 131024 144561 131026
rect 675138 131082 675249 131087
rect 675138 131026 675188 131082
rect 675244 131026 675249 131082
rect 675138 131024 675249 131026
rect 144495 131021 144561 131024
rect 675183 131021 675249 131024
rect 140802 130048 140862 130388
rect 677058 130347 677118 130610
rect 677007 130342 677118 130347
rect 677007 130286 677012 130342
rect 677068 130286 677118 130342
rect 677007 130284 677118 130286
rect 677007 130281 677073 130284
rect 144207 130048 144273 130051
rect 140802 130046 144273 130048
rect 140802 129990 144212 130046
rect 144268 129990 144273 130046
rect 140802 129988 144273 129990
rect 144207 129985 144273 129988
rect 677058 129607 677118 129722
rect 677058 129602 677169 129607
rect 677058 129546 677108 129602
rect 677164 129546 677169 129602
rect 677058 129544 677169 129546
rect 677103 129541 677169 129544
rect 146703 129308 146769 129311
rect 140832 129306 146769 129308
rect 140832 129250 146708 129306
rect 146764 129250 146769 129306
rect 140832 129248 146769 129250
rect 146703 129245 146769 129248
rect 674754 128719 674814 128982
rect 674754 128714 674865 128719
rect 674754 128658 674804 128714
rect 674860 128658 674865 128714
rect 674754 128656 674865 128658
rect 674799 128653 674865 128656
rect 140802 127532 140862 128090
rect 675138 127979 675198 128094
rect 675087 127974 675198 127979
rect 675087 127918 675092 127974
rect 675148 127918 675198 127974
rect 675087 127916 675198 127918
rect 675087 127913 675153 127916
rect 146319 127532 146385 127535
rect 140802 127530 146385 127532
rect 140802 127474 146324 127530
rect 146380 127474 146385 127530
rect 140802 127472 146385 127474
rect 146319 127469 146385 127472
rect 674946 127091 675006 127354
rect 674895 127086 675006 127091
rect 674895 127030 674900 127086
rect 674956 127030 675006 127086
rect 674895 127028 675006 127030
rect 674895 127025 674961 127028
rect 147087 126940 147153 126943
rect 140832 126938 147153 126940
rect 140832 126882 147092 126938
rect 147148 126882 147153 126938
rect 140832 126880 147153 126882
rect 147087 126877 147153 126880
rect 146511 126794 146577 126795
rect 146511 126792 146560 126794
rect 146468 126790 146560 126792
rect 146468 126734 146516 126790
rect 146468 126732 146560 126734
rect 146511 126730 146560 126732
rect 146624 126730 146630 126794
rect 146511 126729 146577 126730
rect 676866 126351 676926 126466
rect 676866 126346 676977 126351
rect 676866 126290 676916 126346
rect 676972 126290 676977 126346
rect 676866 126288 676977 126290
rect 676911 126285 676977 126288
rect 39855 125312 39921 125315
rect 39810 125310 39921 125312
rect 39810 125254 39860 125310
rect 39916 125254 39921 125310
rect 39810 125249 39921 125254
rect 39810 124986 39870 125249
rect 140802 125164 140862 125642
rect 676866 125611 676926 125874
rect 676815 125606 676926 125611
rect 676815 125550 676820 125606
rect 676876 125550 676926 125606
rect 676815 125548 676926 125550
rect 676815 125545 676881 125548
rect 146319 125164 146385 125167
rect 140802 125162 146385 125164
rect 140802 125106 146324 125162
rect 146380 125106 146385 125162
rect 140802 125104 146385 125106
rect 146319 125101 146385 125104
rect 674511 124868 674577 124871
rect 674754 124868 674814 124986
rect 674511 124866 674814 124868
rect 674511 124810 674516 124866
rect 674572 124810 674814 124866
rect 674511 124808 674814 124810
rect 674511 124805 674577 124808
rect 146703 124424 146769 124427
rect 140832 124422 146769 124424
rect 140832 124366 146708 124422
rect 146764 124366 146769 124422
rect 140832 124364 146769 124366
rect 146703 124361 146769 124364
rect 674319 124276 674385 124279
rect 674319 124274 674784 124276
rect 674319 124218 674324 124274
rect 674380 124218 674784 124274
rect 674319 124216 674784 124218
rect 674319 124213 674385 124216
rect 210490 123918 210496 123982
rect 210560 123980 210566 123982
rect 211066 123980 211072 123982
rect 210560 123920 211072 123980
rect 210560 123918 210566 123920
rect 211066 123918 211072 123920
rect 211136 123918 211142 123982
rect 209722 123770 209728 123834
rect 209792 123832 209798 123834
rect 210874 123832 210880 123834
rect 209792 123772 210880 123832
rect 209792 123770 209798 123772
rect 210874 123770 210880 123772
rect 210944 123770 210950 123834
rect 674127 123388 674193 123391
rect 674127 123386 674784 123388
rect 674127 123330 674132 123386
rect 674188 123330 674784 123386
rect 674127 123328 674784 123330
rect 674127 123325 674193 123328
rect 140802 122648 140862 123136
rect 146703 122648 146769 122651
rect 140802 122646 146769 122648
rect 140802 122590 146708 122646
rect 146764 122590 146769 122646
rect 140802 122588 146769 122590
rect 146703 122585 146769 122588
rect 210298 122438 210304 122502
rect 210368 122500 210374 122502
rect 210874 122500 210880 122502
rect 210368 122440 210880 122500
rect 210368 122438 210374 122440
rect 210874 122438 210880 122440
rect 210944 122438 210950 122502
rect 674754 122355 674814 122544
rect 674703 122350 674814 122355
rect 674703 122294 674708 122350
rect 674764 122294 674814 122350
rect 674703 122292 674814 122294
rect 674703 122289 674769 122292
rect 140802 121464 140862 121952
rect 146895 121464 146961 121467
rect 140802 121462 146961 121464
rect 140802 121406 146900 121462
rect 146956 121406 146961 121462
rect 140802 121404 146961 121406
rect 640386 121464 640446 121730
rect 647727 121464 647793 121467
rect 640386 121462 647793 121464
rect 640386 121406 647732 121462
rect 647788 121406 647793 121462
rect 640386 121404 647793 121406
rect 146895 121401 146961 121404
rect 647727 121401 647793 121404
rect 674607 121316 674673 121319
rect 674754 121316 674814 121730
rect 674607 121314 674814 121316
rect 674607 121258 674612 121314
rect 674668 121258 674814 121314
rect 674607 121256 674814 121258
rect 674607 121253 674673 121256
rect 647823 121168 647889 121171
rect 640416 121166 647889 121168
rect 640416 121110 647828 121166
rect 647884 121110 647889 121166
rect 640416 121108 647889 121110
rect 647823 121105 647889 121108
rect 674415 121094 674481 121097
rect 674415 121092 674784 121094
rect 674415 121036 674420 121092
rect 674476 121036 674784 121092
rect 674415 121034 674784 121036
rect 674415 121031 674481 121034
rect 146703 120872 146769 120875
rect 647919 120872 647985 120875
rect 140832 120870 146769 120872
rect 140832 120814 146708 120870
rect 146764 120814 146769 120870
rect 140832 120812 146769 120814
rect 146703 120809 146769 120812
rect 640386 120870 647985 120872
rect 640386 120814 647924 120870
rect 647980 120814 647985 120870
rect 640386 120812 647985 120814
rect 640386 120546 640446 120812
rect 647919 120809 647985 120812
rect 646479 120428 646545 120431
rect 640386 120426 646545 120428
rect 640386 120370 646484 120426
rect 646540 120370 646545 120426
rect 640386 120368 646545 120370
rect 640386 120028 640446 120368
rect 646479 120365 646545 120368
rect 675898 120366 675904 120430
rect 675968 120428 675974 120430
rect 677007 120428 677073 120431
rect 675968 120426 677073 120428
rect 675968 120370 677012 120426
rect 677068 120370 677073 120426
rect 675968 120368 677073 120370
rect 675968 120366 675974 120368
rect 677007 120365 677073 120368
rect 140802 119096 140862 119630
rect 146319 119096 146385 119099
rect 140802 119094 146385 119096
rect 140802 119038 146324 119094
rect 146380 119038 146385 119094
rect 140802 119036 146385 119038
rect 146319 119033 146385 119036
rect 210159 119096 210225 119099
rect 211066 119096 211072 119098
rect 210159 119094 211072 119096
rect 210159 119038 210164 119094
rect 210220 119038 211072 119094
rect 210159 119036 211072 119038
rect 210159 119033 210225 119036
rect 211066 119034 211072 119036
rect 211136 119034 211142 119098
rect 146703 118504 146769 118507
rect 140832 118502 146769 118504
rect 140832 118446 146708 118502
rect 146764 118446 146769 118502
rect 140832 118444 146769 118446
rect 146703 118441 146769 118444
rect 209914 118442 209920 118506
rect 209984 118504 209990 118506
rect 211066 118504 211072 118506
rect 209984 118444 211072 118504
rect 209984 118442 209990 118444
rect 211066 118442 211072 118444
rect 211136 118442 211142 118506
rect 676666 117998 676672 118062
rect 676736 118060 676742 118062
rect 677103 118060 677169 118063
rect 676736 118058 677169 118060
rect 676736 118002 677108 118058
rect 677164 118002 677169 118058
rect 676736 118000 677169 118002
rect 676736 117998 676742 118000
rect 677103 117997 677169 118000
rect 140802 116728 140862 117210
rect 146703 116728 146769 116731
rect 140802 116726 146769 116728
rect 140802 116670 146708 116726
rect 146764 116670 146769 116726
rect 140802 116668 146769 116670
rect 146703 116665 146769 116668
rect 146895 115988 146961 115991
rect 140832 115986 146961 115988
rect 140832 115930 146900 115986
rect 146956 115930 146961 115986
rect 140832 115928 146961 115930
rect 146895 115925 146961 115928
rect 146511 115250 146577 115251
rect 146511 115248 146560 115250
rect 146468 115246 146560 115248
rect 146468 115190 146516 115246
rect 146468 115188 146560 115190
rect 146511 115186 146560 115188
rect 146624 115186 146630 115250
rect 146511 115185 146577 115186
rect 144303 115100 144369 115103
rect 144591 115100 144657 115103
rect 144303 115098 144657 115100
rect 144303 115042 144308 115098
rect 144364 115042 144596 115098
rect 144652 115042 144657 115098
rect 144303 115040 144657 115042
rect 144303 115037 144369 115040
rect 144591 115037 144657 115040
rect 140802 114212 140862 114762
rect 146703 114212 146769 114215
rect 140802 114210 146769 114212
rect 140802 114154 146708 114210
rect 146764 114154 146769 114210
rect 140802 114152 146769 114154
rect 146703 114149 146769 114152
rect 674170 114150 674176 114214
rect 674240 114212 674246 114214
rect 675375 114212 675441 114215
rect 674240 114210 675441 114212
rect 674240 114154 675380 114210
rect 675436 114154 675441 114210
rect 674240 114152 675441 114154
rect 674240 114150 674246 114152
rect 675375 114149 675441 114152
rect 140802 113176 140862 113664
rect 144399 113176 144465 113179
rect 140802 113174 144465 113176
rect 140802 113118 144404 113174
rect 144460 113118 144465 113174
rect 140802 113116 144465 113118
rect 144399 113113 144465 113116
rect 146703 112436 146769 112439
rect 140832 112434 146769 112436
rect 140832 112378 146708 112434
rect 146764 112378 146769 112434
rect 140832 112376 146769 112378
rect 146703 112373 146769 112376
rect 144399 111252 144465 111255
rect 140832 111250 144465 111252
rect 140832 111194 144404 111250
rect 144460 111194 144465 111250
rect 140832 111192 144465 111194
rect 144399 111189 144465 111192
rect 675375 110070 675441 110071
rect 675322 110068 675328 110070
rect 675284 110008 675328 110068
rect 675392 110066 675441 110070
rect 675436 110010 675441 110066
rect 675322 110006 675328 110008
rect 675392 110006 675441 110010
rect 675375 110005 675441 110006
rect 140802 109772 140862 109964
rect 146703 109772 146769 109775
rect 140802 109770 146769 109772
rect 140802 109714 146708 109770
rect 146764 109714 146769 109770
rect 140802 109712 146769 109714
rect 146703 109709 146769 109712
rect 674746 109266 674752 109330
rect 674816 109328 674822 109330
rect 675087 109328 675153 109331
rect 674816 109326 675153 109328
rect 674816 109270 675092 109326
rect 675148 109270 675153 109326
rect 674816 109268 675153 109270
rect 674816 109266 674822 109268
rect 675087 109265 675153 109268
rect 140802 108292 140862 108778
rect 144399 108292 144465 108295
rect 140802 108290 144465 108292
rect 140802 108234 144404 108290
rect 144460 108234 144465 108290
rect 140802 108232 144465 108234
rect 144399 108229 144465 108232
rect 675759 108144 675825 108147
rect 675898 108144 675904 108146
rect 675759 108142 675904 108144
rect 675759 108086 675764 108142
rect 675820 108086 675904 108142
rect 675759 108084 675904 108086
rect 675759 108081 675825 108084
rect 675898 108082 675904 108084
rect 675968 108082 675974 108146
rect 146703 107552 146769 107555
rect 140832 107550 146769 107552
rect 140832 107494 146708 107550
rect 146764 107494 146769 107550
rect 140832 107492 146769 107494
rect 146703 107489 146769 107492
rect 210106 106750 210112 106814
rect 210176 106812 210182 106814
rect 210874 106812 210880 106814
rect 210176 106752 210880 106812
rect 210176 106750 210182 106752
rect 210874 106750 210880 106752
rect 210944 106750 210950 106814
rect 144442 106454 144448 106518
rect 144512 106516 144518 106518
rect 144687 106516 144753 106519
rect 675087 106516 675153 106519
rect 144512 106514 144753 106516
rect 144512 106458 144692 106514
rect 144748 106458 144753 106514
rect 144512 106456 144753 106458
rect 144512 106454 144518 106456
rect 144687 106453 144753 106456
rect 665442 106514 675153 106516
rect 665442 106458 675092 106514
rect 675148 106458 675153 106514
rect 665442 106456 675153 106458
rect 140802 105924 140862 106412
rect 665442 106080 665502 106456
rect 675087 106453 675153 106456
rect 144303 105924 144369 105927
rect 140802 105922 144369 105924
rect 140802 105866 144308 105922
rect 144364 105866 144369 105922
rect 140802 105864 144369 105866
rect 144303 105861 144369 105864
rect 140802 104740 140862 105228
rect 665346 105184 665406 105359
rect 668175 105184 668241 105187
rect 665346 105182 668241 105184
rect 665346 105126 668180 105182
rect 668236 105126 668241 105182
rect 665346 105124 668241 105126
rect 668175 105121 668241 105124
rect 144111 104740 144177 104743
rect 140802 104738 144177 104740
rect 140802 104682 144116 104738
rect 144172 104682 144177 104738
rect 140802 104680 144177 104682
rect 144111 104677 144177 104680
rect 665154 104595 665214 104994
rect 665154 104590 665265 104595
rect 665154 104534 665204 104590
rect 665260 104534 665265 104590
rect 665154 104532 665265 104534
rect 665199 104529 665265 104532
rect 647919 104296 647985 104299
rect 640416 104294 647985 104296
rect 640416 104238 647924 104294
rect 647980 104238 647985 104294
rect 640416 104236 647985 104238
rect 647919 104233 647985 104236
rect 144783 104000 144849 104003
rect 140832 103998 144849 104000
rect 140832 103942 144788 103998
rect 144844 103942 144849 103998
rect 140832 103940 144849 103942
rect 144783 103937 144849 103940
rect 144303 103704 144369 103707
rect 144442 103704 144448 103706
rect 144303 103702 144448 103704
rect 144303 103646 144308 103702
rect 144364 103646 144448 103702
rect 144303 103644 144448 103646
rect 144303 103641 144369 103644
rect 144442 103642 144448 103644
rect 144512 103642 144518 103706
rect 674938 103198 674944 103262
rect 675008 103260 675014 103262
rect 675375 103260 675441 103263
rect 675008 103258 675441 103260
rect 675008 103202 675380 103258
rect 675436 103202 675441 103258
rect 675008 103200 675441 103202
rect 675008 103198 675014 103200
rect 675375 103197 675441 103200
rect 144111 102816 144177 102819
rect 140832 102814 144177 102816
rect 140832 102758 144116 102814
rect 144172 102758 144177 102814
rect 140832 102756 144177 102758
rect 144111 102753 144177 102756
rect 204495 102076 204561 102079
rect 204495 102074 210528 102076
rect 204495 102018 204500 102074
rect 204556 102018 210528 102074
rect 204495 102016 210528 102018
rect 204495 102013 204561 102016
rect 144015 101632 144081 101635
rect 140832 101630 144081 101632
rect 140832 101574 144020 101630
rect 144076 101574 144081 101630
rect 140832 101572 144081 101574
rect 144015 101569 144081 101572
rect 206703 101632 206769 101635
rect 206703 101630 210528 101632
rect 206703 101574 206708 101630
rect 206764 101574 210528 101630
rect 206703 101572 210528 101574
rect 206703 101569 206769 101572
rect 675759 101484 675825 101487
rect 676666 101484 676672 101486
rect 675759 101482 676672 101484
rect 675759 101426 675764 101482
rect 675820 101426 676672 101482
rect 675759 101424 676672 101426
rect 675759 101421 675825 101424
rect 676666 101422 676672 101424
rect 676736 101422 676742 101486
rect 206223 101040 206289 101043
rect 206223 101038 210528 101040
rect 206223 100982 206228 101038
rect 206284 100982 210528 101038
rect 206223 100980 210528 100982
rect 206223 100977 206289 100980
rect 204495 100448 204561 100451
rect 204495 100446 210528 100448
rect 204495 100390 204500 100446
rect 204556 100390 210528 100446
rect 204495 100388 210528 100390
rect 204495 100385 204561 100388
rect 140802 99856 140862 100344
rect 204591 100300 204657 100303
rect 204591 100298 210558 100300
rect 204591 100242 204596 100298
rect 204652 100242 210558 100298
rect 204591 100240 210558 100242
rect 204591 100237 204657 100240
rect 210498 99900 210558 100240
rect 144303 99856 144369 99859
rect 140802 99854 144369 99856
rect 140802 99798 144308 99854
rect 144364 99798 144369 99854
rect 140802 99796 144369 99798
rect 144303 99793 144369 99796
rect 204783 99412 204849 99415
rect 204783 99410 210528 99412
rect 204783 99354 204788 99410
rect 204844 99354 210528 99410
rect 204783 99352 210528 99354
rect 204783 99349 204849 99352
rect 144111 99116 144177 99119
rect 140832 99114 144177 99116
rect 140832 99058 144116 99114
rect 144172 99058 144177 99114
rect 140832 99056 144177 99058
rect 144111 99053 144177 99056
rect 206895 98820 206961 98823
rect 206895 98818 210528 98820
rect 206895 98762 206900 98818
rect 206956 98762 210528 98818
rect 206895 98760 210528 98762
rect 206895 98757 206961 98760
rect 204687 98672 204753 98675
rect 204687 98670 210558 98672
rect 204687 98614 204692 98670
rect 204748 98614 210558 98670
rect 204687 98612 210558 98614
rect 204687 98609 204753 98612
rect 210498 98272 210558 98612
rect 144015 98080 144081 98083
rect 140832 98078 144081 98080
rect 140832 98022 144020 98078
rect 144076 98022 144081 98078
rect 140832 98020 144081 98022
rect 144015 98017 144081 98020
rect 204495 97784 204561 97787
rect 204495 97782 210528 97784
rect 204495 97726 204500 97782
rect 204556 97726 210528 97782
rect 204495 97724 210528 97726
rect 204495 97721 204561 97724
rect 204495 97192 204561 97195
rect 204495 97190 210528 97192
rect 204495 97134 204500 97190
rect 204556 97134 210528 97190
rect 204495 97132 210528 97134
rect 204495 97129 204561 97132
rect 206127 97044 206193 97047
rect 206127 97042 210558 97044
rect 206127 96986 206132 97042
rect 206188 96986 210558 97042
rect 206127 96984 210558 96986
rect 206127 96981 206193 96984
rect 140802 96304 140862 96792
rect 210498 96644 210558 96984
rect 210682 96834 210688 96898
rect 210752 96896 210758 96898
rect 211066 96896 211072 96898
rect 210752 96836 211072 96896
rect 210752 96834 210758 96836
rect 211066 96834 211072 96836
rect 211136 96834 211142 96898
rect 144111 96304 144177 96307
rect 140802 96302 144177 96304
rect 140802 96246 144116 96302
rect 144172 96246 144177 96302
rect 140802 96244 144177 96246
rect 144111 96241 144177 96244
rect 205263 96156 205329 96159
rect 205263 96154 210528 96156
rect 205263 96098 205268 96154
rect 205324 96098 210528 96154
rect 205263 96096 210528 96098
rect 205263 96093 205329 96096
rect 210298 95798 210304 95862
rect 210368 95860 210374 95862
rect 211066 95860 211072 95862
rect 210368 95800 211072 95860
rect 210368 95798 210374 95800
rect 211066 95798 211072 95800
rect 211136 95798 211142 95862
rect 144015 95564 144081 95567
rect 140832 95562 144081 95564
rect 140832 95506 144020 95562
rect 144076 95506 144081 95562
rect 140832 95504 144081 95506
rect 144015 95501 144081 95504
rect 206511 95564 206577 95567
rect 206511 95562 210528 95564
rect 206511 95506 206516 95562
rect 206572 95506 210528 95562
rect 206511 95504 210528 95506
rect 206511 95501 206577 95504
rect 204495 94676 204561 94679
rect 210498 94676 210558 95016
rect 204495 94674 210558 94676
rect 204495 94618 204500 94674
rect 204556 94618 210558 94674
rect 204495 94616 210558 94618
rect 204495 94613 204561 94616
rect 205743 94528 205809 94531
rect 205743 94526 210528 94528
rect 205743 94470 205748 94526
rect 205804 94470 210528 94526
rect 205743 94468 210528 94470
rect 205743 94465 205809 94468
rect 144111 94380 144177 94383
rect 140832 94378 144177 94380
rect 140832 94322 144116 94378
rect 144172 94322 144177 94378
rect 140832 94320 144177 94322
rect 144111 94317 144177 94320
rect 210159 94232 210225 94235
rect 211066 94232 211072 94234
rect 210159 94230 211072 94232
rect 210159 94174 210164 94230
rect 210220 94174 211072 94230
rect 210159 94172 211072 94174
rect 210159 94169 210225 94172
rect 211066 94170 211072 94172
rect 211136 94170 211142 94234
rect 205839 93936 205905 93939
rect 205839 93934 210528 93936
rect 205839 93878 205844 93934
rect 205900 93878 210528 93934
rect 205839 93876 210528 93878
rect 205839 93873 205905 93876
rect 204591 93788 204657 93791
rect 204591 93786 210558 93788
rect 204591 93730 204596 93786
rect 204652 93730 210558 93786
rect 204591 93728 210558 93730
rect 204591 93725 204657 93728
rect 210498 93388 210558 93728
rect 210106 93134 210112 93198
rect 210176 93196 210182 93198
rect 211066 93196 211072 93198
rect 210176 93136 211072 93196
rect 210176 93134 210182 93136
rect 211066 93134 211072 93136
rect 211136 93134 211142 93198
rect 140802 92752 140862 93092
rect 210298 92986 210304 93050
rect 210368 93048 210374 93050
rect 211066 93048 211072 93050
rect 210368 92988 211072 93048
rect 210368 92986 210374 92988
rect 211066 92986 211072 92988
rect 211136 92986 211142 93050
rect 206895 92900 206961 92903
rect 206895 92898 210528 92900
rect 206895 92842 206900 92898
rect 206956 92842 210528 92898
rect 206895 92840 210528 92842
rect 206895 92837 206961 92840
rect 144015 92752 144081 92755
rect 140802 92750 144081 92752
rect 140802 92694 144020 92750
rect 144076 92694 144081 92750
rect 140802 92692 144081 92694
rect 144015 92689 144081 92692
rect 206319 92308 206385 92311
rect 206319 92306 210528 92308
rect 206319 92250 206324 92306
rect 206380 92250 210528 92306
rect 206319 92248 210528 92250
rect 206319 92245 206385 92248
rect 204591 92012 204657 92015
rect 204591 92010 210558 92012
rect 204591 91954 204596 92010
rect 204652 91954 210558 92010
rect 204591 91952 210558 91954
rect 204591 91949 204657 91952
rect 140802 91420 140862 91908
rect 210498 91760 210558 91952
rect 144111 91420 144177 91423
rect 140802 91418 144177 91420
rect 140802 91362 144116 91418
rect 144172 91362 144177 91418
rect 140802 91360 144177 91362
rect 144111 91357 144177 91360
rect 204495 91272 204561 91275
rect 204495 91270 210528 91272
rect 204495 91214 204500 91270
rect 204556 91214 210528 91270
rect 204495 91212 210528 91214
rect 204495 91209 204561 91212
rect 144303 90828 144369 90831
rect 140832 90826 144369 90828
rect 140832 90770 144308 90826
rect 144364 90770 144369 90826
rect 140832 90768 144369 90770
rect 144303 90765 144369 90768
rect 204687 90680 204753 90683
rect 204687 90678 210528 90680
rect 204687 90622 204692 90678
rect 204748 90622 210528 90678
rect 204687 90620 210528 90622
rect 204687 90617 204753 90620
rect 204591 90088 204657 90091
rect 204591 90086 210528 90088
rect 204591 90030 204596 90086
rect 204652 90030 210528 90086
rect 204591 90028 210528 90030
rect 204591 90025 204657 90028
rect 144015 89644 144081 89647
rect 140832 89642 144081 89644
rect 140832 89586 144020 89642
rect 144076 89586 144081 89642
rect 140832 89584 144081 89586
rect 144015 89581 144081 89584
rect 204783 89644 204849 89647
rect 204783 89642 210528 89644
rect 204783 89586 204788 89642
rect 204844 89586 210528 89642
rect 204783 89584 210528 89586
rect 204783 89581 204849 89584
rect 204783 89052 204849 89055
rect 647631 89052 647697 89055
rect 204783 89050 210528 89052
rect 204783 88994 204788 89050
rect 204844 88994 210528 89050
rect 204783 88992 210528 88994
rect 640416 89050 647697 89052
rect 640416 88994 647636 89050
rect 647692 88994 647697 89050
rect 640416 88992 647697 88994
rect 204783 88989 204849 88992
rect 647631 88989 647697 88992
rect 204495 88460 204561 88463
rect 204495 88458 210528 88460
rect 204495 88402 204500 88458
rect 204556 88402 210528 88458
rect 204495 88400 210528 88402
rect 204495 88397 204561 88400
rect 140802 87868 140862 88356
rect 640194 88164 640254 88430
rect 646863 88164 646929 88167
rect 640194 88162 646929 88164
rect 640194 88106 646868 88162
rect 646924 88106 646929 88162
rect 640194 88104 646929 88106
rect 646863 88101 646929 88104
rect 204591 88016 204657 88019
rect 204591 88014 210528 88016
rect 204591 87958 204596 88014
rect 204652 87958 210528 88014
rect 204591 87956 210528 87958
rect 204591 87953 204657 87956
rect 144111 87868 144177 87871
rect 140802 87866 144177 87868
rect 140802 87810 144116 87866
rect 144172 87810 144177 87866
rect 140802 87808 144177 87810
rect 144111 87805 144177 87808
rect 640386 87720 640446 87986
rect 647919 87720 647985 87723
rect 640386 87718 647985 87720
rect 640386 87662 647924 87718
rect 647980 87662 647985 87718
rect 640386 87660 647985 87662
rect 647919 87657 647985 87660
rect 205263 87424 205329 87427
rect 647439 87424 647505 87427
rect 205263 87422 210528 87424
rect 205263 87366 205268 87422
rect 205324 87366 210528 87422
rect 205263 87364 210528 87366
rect 640416 87422 647505 87424
rect 640416 87366 647444 87422
rect 647500 87366 647505 87422
rect 640416 87364 647505 87366
rect 205263 87361 205329 87364
rect 647439 87361 647505 87364
rect 146511 87128 146577 87131
rect 140832 87126 146577 87128
rect 140832 87070 146516 87126
rect 146572 87070 146577 87126
rect 140832 87068 146577 87070
rect 146511 87065 146577 87068
rect 650991 86980 651057 86983
rect 650991 86978 656736 86980
rect 650991 86922 650996 86978
rect 651052 86922 656736 86978
rect 650991 86920 656736 86922
rect 650991 86917 651057 86920
rect 204687 86832 204753 86835
rect 204687 86830 210528 86832
rect 204687 86774 204692 86830
rect 204748 86774 210528 86830
rect 204687 86772 210528 86774
rect 204687 86769 204753 86772
rect 640194 86536 640254 86802
rect 647919 86536 647985 86539
rect 640194 86534 647985 86536
rect 640194 86478 647924 86534
rect 647980 86478 647985 86534
rect 640194 86476 647985 86478
rect 647919 86473 647985 86476
rect 204495 86388 204561 86391
rect 204495 86386 210528 86388
rect 204495 86330 204500 86386
rect 204556 86330 210528 86386
rect 204495 86328 210528 86330
rect 204495 86325 204561 86328
rect 640386 86240 640446 86358
rect 647823 86240 647889 86243
rect 640386 86238 647889 86240
rect 640386 86182 647828 86238
rect 647884 86182 647889 86238
rect 640386 86180 647889 86182
rect 647823 86177 647889 86180
rect 651183 86240 651249 86243
rect 651183 86238 656736 86240
rect 651183 86182 651188 86238
rect 651244 86182 656736 86238
rect 651183 86180 656736 86182
rect 651183 86177 651249 86180
rect 146703 85944 146769 85947
rect 140832 85942 146769 85944
rect 140832 85886 146708 85942
rect 146764 85886 146769 85942
rect 140832 85884 146769 85886
rect 146703 85881 146769 85884
rect 204495 85796 204561 85799
rect 646191 85796 646257 85799
rect 204495 85794 210528 85796
rect 204495 85738 204500 85794
rect 204556 85738 210528 85794
rect 204495 85736 210528 85738
rect 640416 85794 646257 85796
rect 640416 85738 646196 85794
rect 646252 85738 646257 85794
rect 640416 85736 646257 85738
rect 204495 85733 204561 85736
rect 646191 85733 646257 85736
rect 663426 85651 663486 86210
rect 663375 85646 663486 85651
rect 663375 85590 663380 85646
rect 663436 85590 663486 85646
rect 663375 85588 663486 85590
rect 663375 85585 663441 85588
rect 647727 85500 647793 85503
rect 640386 85498 647793 85500
rect 640386 85442 647732 85498
rect 647788 85442 647793 85498
rect 640386 85440 647793 85442
rect 205551 85204 205617 85207
rect 205551 85202 210528 85204
rect 205551 85146 205556 85202
rect 205612 85146 210528 85202
rect 640386 85174 640446 85440
rect 647727 85437 647793 85440
rect 650895 85352 650961 85355
rect 650895 85350 656736 85352
rect 650895 85294 650900 85350
rect 650956 85294 656736 85350
rect 650895 85292 656736 85294
rect 650895 85289 650961 85292
rect 663279 85204 663345 85207
rect 663234 85202 663345 85204
rect 205551 85144 210528 85146
rect 663234 85146 663284 85202
rect 663340 85146 663345 85202
rect 205551 85141 205617 85144
rect 663234 85141 663345 85146
rect 646863 85056 646929 85059
rect 640194 85054 646929 85056
rect 640194 84998 646868 85054
rect 646924 84998 646929 85054
rect 640194 84996 646929 84998
rect 204591 84760 204657 84763
rect 204591 84758 210528 84760
rect 204591 84702 204596 84758
rect 204652 84702 210528 84758
rect 640194 84730 640254 84996
rect 646863 84993 646929 84996
rect 204591 84700 210528 84702
rect 204591 84697 204657 84700
rect 140802 84168 140862 84656
rect 663234 84582 663294 85141
rect 663426 84763 663486 85322
rect 663426 84758 663537 84763
rect 663426 84702 663476 84758
rect 663532 84702 663537 84758
rect 663426 84700 663537 84702
rect 663471 84697 663537 84700
rect 650991 84316 651057 84319
rect 650991 84314 656736 84316
rect 650991 84258 650996 84314
rect 651052 84258 656736 84314
rect 650991 84256 656736 84258
rect 650991 84253 651057 84256
rect 146319 84168 146385 84171
rect 140802 84166 146385 84168
rect 140802 84110 146324 84166
rect 146380 84110 146385 84166
rect 140802 84108 146385 84110
rect 146319 84105 146385 84108
rect 206607 84168 206673 84171
rect 645903 84168 645969 84171
rect 206607 84166 210528 84168
rect 206607 84110 206612 84166
rect 206668 84110 210528 84166
rect 206607 84108 210528 84110
rect 640416 84166 645969 84168
rect 640416 84110 645908 84166
rect 645964 84110 645969 84166
rect 640416 84108 645969 84110
rect 206607 84105 206673 84108
rect 645903 84105 645969 84108
rect 647247 83872 647313 83875
rect 640386 83870 647313 83872
rect 640386 83814 647252 83870
rect 647308 83814 647313 83870
rect 640386 83812 647313 83814
rect 140802 83576 140862 83618
rect 144591 83576 144657 83579
rect 140802 83574 144657 83576
rect 140802 83518 144596 83574
rect 144652 83518 144657 83574
rect 140802 83516 144657 83518
rect 144591 83513 144657 83516
rect 204687 83576 204753 83579
rect 204687 83574 210528 83576
rect 204687 83518 204692 83574
rect 204748 83518 210528 83574
rect 640386 83546 640446 83812
rect 647247 83809 647313 83812
rect 204687 83516 210528 83518
rect 204687 83513 204753 83516
rect 647919 83428 647985 83431
rect 640194 83426 647985 83428
rect 640194 83370 647924 83426
rect 647980 83370 647985 83426
rect 640194 83368 647985 83370
rect 204495 83132 204561 83135
rect 204495 83130 210528 83132
rect 204495 83074 204500 83130
rect 204556 83074 210528 83130
rect 640194 83102 640254 83368
rect 647919 83365 647985 83368
rect 651087 83428 651153 83431
rect 651087 83426 656736 83428
rect 651087 83370 651092 83426
rect 651148 83370 656736 83426
rect 651087 83368 656736 83370
rect 651087 83365 651153 83368
rect 204495 83072 210528 83074
rect 204495 83069 204561 83072
rect 663426 82839 663486 83398
rect 663375 82834 663486 82839
rect 663375 82778 663380 82834
rect 663436 82778 663486 82834
rect 663375 82776 663486 82778
rect 663375 82773 663441 82776
rect 650895 82688 650961 82691
rect 650895 82686 656736 82688
rect 650895 82630 650900 82686
rect 650956 82630 656736 82686
rect 650895 82628 656736 82630
rect 650895 82625 650961 82628
rect 205743 82540 205809 82543
rect 647919 82540 647985 82543
rect 205743 82538 210528 82540
rect 205743 82482 205748 82538
rect 205804 82482 210528 82538
rect 205743 82480 210528 82482
rect 640416 82538 647985 82540
rect 640416 82482 647924 82538
rect 647980 82482 647985 82538
rect 640416 82480 647985 82482
rect 205743 82477 205809 82480
rect 647919 82477 647985 82480
rect 146703 82392 146769 82395
rect 140832 82390 146769 82392
rect 140832 82334 146708 82390
rect 146764 82334 146769 82390
rect 140832 82332 146769 82334
rect 146703 82329 146769 82332
rect 209914 82182 209920 82246
rect 209984 82244 209990 82246
rect 210874 82244 210880 82246
rect 209984 82184 210880 82244
rect 209984 82182 209990 82184
rect 210874 82182 210880 82184
rect 210944 82182 210950 82246
rect 647535 82244 647601 82247
rect 640386 82242 647601 82244
rect 640386 82186 647540 82242
rect 647596 82186 647601 82242
rect 640386 82184 647601 82186
rect 204495 81948 204561 81951
rect 204495 81946 210528 81948
rect 204495 81890 204500 81946
rect 204556 81890 210528 81946
rect 640386 81918 640446 82184
rect 647535 82181 647601 82184
rect 663234 82099 663294 82658
rect 663234 82094 663345 82099
rect 663234 82038 663284 82094
rect 663340 82038 663345 82094
rect 663234 82036 663345 82038
rect 663279 82033 663345 82036
rect 204495 81888 210528 81890
rect 204495 81885 204561 81888
rect 206703 81504 206769 81507
rect 206703 81502 210528 81504
rect 206703 81446 206708 81502
rect 206764 81446 210528 81502
rect 206703 81444 210528 81446
rect 206703 81441 206769 81444
rect 640386 81356 640446 81474
rect 647919 81356 647985 81359
rect 640386 81354 647985 81356
rect 640386 81298 647924 81354
rect 647980 81298 647985 81354
rect 640386 81296 647985 81298
rect 647919 81293 647985 81296
rect 140802 80764 140862 81170
rect 210490 81146 210496 81210
rect 210560 81208 210566 81210
rect 211066 81208 211072 81210
rect 210560 81148 211072 81208
rect 210560 81146 210566 81148
rect 211066 81146 211072 81148
rect 211136 81146 211142 81210
rect 662895 81208 662961 81211
rect 663042 81208 663102 81770
rect 662895 81206 663102 81208
rect 662895 81150 662900 81206
rect 662956 81150 663102 81206
rect 662895 81148 663102 81150
rect 662895 81145 662961 81148
rect 206223 80912 206289 80915
rect 647343 80912 647409 80915
rect 206223 80910 210528 80912
rect 206223 80854 206228 80910
rect 206284 80854 210528 80910
rect 206223 80852 210528 80854
rect 640416 80910 647409 80912
rect 640416 80854 647348 80910
rect 647404 80854 647409 80910
rect 640416 80852 647409 80854
rect 206223 80849 206289 80852
rect 647343 80849 647409 80852
rect 144399 80764 144465 80767
rect 140802 80762 144465 80764
rect 140802 80706 144404 80762
rect 144460 80706 144465 80762
rect 140802 80704 144465 80706
rect 144399 80701 144465 80704
rect 647823 80468 647889 80471
rect 640386 80466 647889 80468
rect 640386 80410 647828 80466
rect 647884 80410 647889 80466
rect 640386 80408 647889 80410
rect 205263 80320 205329 80323
rect 205263 80318 210528 80320
rect 205263 80262 205268 80318
rect 205324 80262 210528 80318
rect 640386 80290 640446 80408
rect 647823 80405 647889 80408
rect 205263 80260 210528 80262
rect 205263 80257 205329 80260
rect 204495 80172 204561 80175
rect 647919 80172 647985 80175
rect 204495 80170 210558 80172
rect 204495 80114 204500 80170
rect 204556 80114 210558 80170
rect 204495 80112 210558 80114
rect 204495 80109 204561 80112
rect 140802 79432 140862 79920
rect 210498 79772 210558 80112
rect 640386 80170 647985 80172
rect 640386 80114 647924 80170
rect 647980 80114 647985 80170
rect 640386 80112 647985 80114
rect 640386 79772 640446 80112
rect 647919 80109 647985 80112
rect 146703 79432 146769 79435
rect 140802 79430 146769 79432
rect 140802 79374 146708 79430
rect 146764 79374 146769 79430
rect 140802 79372 146769 79374
rect 146703 79369 146769 79372
rect 204591 79284 204657 79287
rect 647919 79284 647985 79287
rect 204591 79282 210528 79284
rect 204591 79226 204596 79282
rect 204652 79226 210528 79282
rect 204591 79224 210528 79226
rect 640416 79282 647985 79284
rect 640416 79226 647924 79282
rect 647980 79226 647985 79282
rect 640416 79224 647985 79226
rect 204591 79221 204657 79224
rect 647919 79221 647985 79224
rect 647727 78988 647793 78991
rect 640386 78986 647793 78988
rect 640386 78930 647732 78986
rect 647788 78930 647793 78986
rect 640386 78928 647793 78930
rect 144303 78692 144369 78695
rect 140832 78690 144369 78692
rect 140832 78634 144308 78690
rect 144364 78634 144369 78690
rect 140832 78632 144369 78634
rect 144303 78629 144369 78632
rect 204687 78692 204753 78695
rect 204687 78690 210528 78692
rect 204687 78634 204692 78690
rect 204748 78634 210528 78690
rect 640386 78662 640446 78928
rect 647727 78925 647793 78928
rect 204687 78632 210528 78634
rect 204687 78629 204753 78632
rect 645423 78544 645489 78547
rect 640386 78542 645489 78544
rect 640386 78486 645428 78542
rect 645484 78486 645489 78542
rect 640386 78484 645489 78486
rect 210159 78174 210225 78177
rect 210159 78172 210528 78174
rect 210159 78116 210164 78172
rect 210220 78116 210528 78172
rect 640386 78144 640446 78484
rect 645423 78481 645489 78484
rect 210159 78114 210528 78116
rect 210159 78111 210225 78114
rect 209722 77742 209728 77806
rect 209792 77804 209798 77806
rect 210874 77804 210880 77806
rect 209792 77744 210880 77804
rect 209792 77742 209798 77744
rect 210874 77742 210880 77744
rect 210944 77742 210950 77806
rect 204783 77656 204849 77659
rect 647919 77656 647985 77659
rect 204783 77654 210528 77656
rect 204783 77598 204788 77654
rect 204844 77598 210528 77654
rect 204783 77596 210528 77598
rect 640416 77654 647985 77656
rect 640416 77598 647924 77654
rect 647980 77598 647985 77654
rect 640416 77596 647985 77598
rect 204783 77593 204849 77596
rect 647919 77593 647985 77596
rect 144303 77508 144369 77511
rect 140832 77506 144369 77508
rect 140832 77450 144308 77506
rect 144364 77450 144369 77506
rect 140832 77448 144369 77450
rect 144303 77445 144369 77448
rect 204591 77064 204657 77067
rect 647919 77064 647985 77067
rect 204591 77062 210528 77064
rect 204591 77006 204596 77062
rect 204652 77006 210528 77062
rect 204591 77004 210528 77006
rect 640416 77062 647985 77064
rect 640416 77006 647924 77062
rect 647980 77006 647985 77062
rect 640416 77004 647985 77006
rect 204591 77001 204657 77004
rect 647919 77001 647985 77004
rect 205935 76916 206001 76919
rect 646479 76916 646545 76919
rect 205935 76914 210558 76916
rect 205935 76858 205940 76914
rect 205996 76858 210558 76914
rect 205935 76856 210558 76858
rect 205935 76853 206001 76856
rect 210498 76516 210558 76856
rect 640386 76914 646545 76916
rect 640386 76858 646484 76914
rect 646540 76858 646545 76914
rect 640386 76856 646545 76858
rect 640386 76516 640446 76856
rect 646479 76853 646545 76856
rect 140802 75732 140862 76220
rect 204495 76028 204561 76031
rect 646479 76028 646545 76031
rect 204495 76026 210528 76028
rect 204495 75970 204500 76026
rect 204556 75970 210528 76026
rect 204495 75968 210528 75970
rect 640416 76026 646545 76028
rect 640416 75970 646484 76026
rect 646540 75970 646545 76026
rect 640416 75968 646545 75970
rect 204495 75965 204561 75968
rect 646479 75965 646545 75968
rect 146511 75732 146577 75735
rect 140802 75730 146577 75732
rect 140802 75674 146516 75730
rect 146572 75674 146577 75730
rect 140802 75672 146577 75674
rect 146511 75669 146577 75672
rect 206511 75436 206577 75439
rect 646479 75436 646545 75439
rect 206511 75434 210528 75436
rect 206511 75378 206516 75434
rect 206572 75378 210528 75434
rect 206511 75376 210528 75378
rect 640416 75434 646545 75436
rect 640416 75378 646484 75434
rect 646540 75378 646545 75434
rect 640416 75376 646545 75378
rect 206511 75373 206577 75376
rect 646479 75373 646545 75376
rect 204687 75288 204753 75291
rect 646095 75288 646161 75291
rect 204687 75286 210558 75288
rect 204687 75230 204692 75286
rect 204748 75230 210558 75286
rect 204687 75228 210558 75230
rect 204687 75225 204753 75228
rect 140802 75140 140862 75184
rect 144015 75140 144081 75143
rect 140802 75138 144081 75140
rect 140802 75082 144020 75138
rect 144076 75082 144081 75138
rect 140802 75080 144081 75082
rect 144015 75077 144081 75080
rect 144111 74992 144177 74995
rect 146511 74992 146577 74995
rect 144111 74990 146577 74992
rect 144111 74934 144116 74990
rect 144172 74934 146516 74990
rect 146572 74934 146577 74990
rect 144111 74932 146577 74934
rect 144111 74929 144177 74932
rect 146511 74929 146577 74932
rect 210498 74888 210558 75228
rect 640386 75286 646161 75288
rect 640386 75230 646100 75286
rect 646156 75230 646161 75286
rect 640386 75228 646161 75230
rect 640386 74888 640446 75228
rect 646095 75225 646161 75228
rect 204495 74400 204561 74403
rect 647247 74400 647313 74403
rect 204495 74398 210528 74400
rect 204495 74342 204500 74398
rect 204556 74342 210528 74398
rect 204495 74340 210528 74342
rect 640416 74398 647313 74400
rect 640416 74342 647252 74398
rect 647308 74342 647313 74398
rect 640416 74340 647313 74342
rect 204495 74337 204561 74340
rect 647247 74337 647313 74340
rect 146031 73956 146097 73959
rect 140832 73954 146097 73956
rect 140832 73898 146036 73954
rect 146092 73898 146097 73954
rect 140832 73896 146097 73898
rect 146031 73893 146097 73896
rect 205743 73808 205809 73811
rect 646863 73808 646929 73811
rect 205743 73806 210528 73808
rect 205743 73750 205748 73806
rect 205804 73750 210528 73806
rect 205743 73748 210528 73750
rect 640416 73806 646929 73808
rect 640416 73750 646868 73806
rect 646924 73750 646929 73806
rect 640416 73748 646929 73750
rect 205743 73745 205809 73748
rect 646863 73745 646929 73748
rect 204591 73660 204657 73663
rect 204591 73658 210558 73660
rect 204591 73602 204596 73658
rect 204652 73602 210558 73658
rect 204591 73600 210558 73602
rect 204591 73597 204657 73600
rect 210498 73260 210558 73600
rect 640386 72920 640446 73260
rect 646095 72920 646161 72923
rect 640386 72918 646161 72920
rect 640386 72862 646100 72918
rect 646156 72862 646161 72918
rect 640386 72860 646161 72862
rect 646095 72857 646161 72860
rect 144111 72772 144177 72775
rect 140832 72770 144177 72772
rect 140832 72714 144116 72770
rect 144172 72714 144177 72770
rect 140832 72712 144177 72714
rect 144111 72709 144177 72712
rect 206799 72772 206865 72775
rect 206799 72770 210528 72772
rect 206799 72714 206804 72770
rect 206860 72714 210528 72770
rect 206799 72712 210528 72714
rect 206799 72709 206865 72712
rect 640386 72624 640446 72742
rect 646671 72624 646737 72627
rect 640386 72622 646737 72624
rect 640386 72566 646676 72622
rect 646732 72566 646737 72622
rect 640386 72564 646737 72566
rect 646671 72561 646737 72564
rect 204687 72180 204753 72183
rect 646479 72180 646545 72183
rect 204687 72178 210528 72180
rect 204687 72122 204692 72178
rect 204748 72122 210528 72178
rect 204687 72120 210528 72122
rect 640416 72178 646545 72180
rect 640416 72122 646484 72178
rect 646540 72122 646545 72178
rect 640416 72120 646545 72122
rect 204687 72117 204753 72120
rect 646479 72117 646545 72120
rect 204495 71736 204561 71739
rect 204495 71734 210558 71736
rect 204495 71678 204500 71734
rect 204556 71678 210558 71734
rect 204495 71676 210558 71678
rect 204495 71673 204561 71676
rect 210498 71632 210558 71676
rect 140802 70996 140862 71484
rect 204591 71144 204657 71147
rect 204591 71142 210528 71144
rect 204591 71086 204596 71142
rect 204652 71086 210528 71142
rect 204591 71084 210528 71086
rect 204591 71081 204657 71084
rect 144015 70996 144081 70999
rect 140802 70994 144081 70996
rect 140802 70938 144020 70994
rect 144076 70938 144081 70994
rect 140802 70936 144081 70938
rect 144015 70933 144081 70936
rect 205455 70552 205521 70555
rect 205455 70550 210528 70552
rect 205455 70494 205460 70550
rect 205516 70494 210528 70550
rect 205455 70492 210528 70494
rect 205455 70489 205521 70492
rect 140802 69812 140862 70290
rect 206799 69960 206865 69963
rect 206799 69958 210528 69960
rect 206799 69902 206804 69958
rect 206860 69902 210528 69958
rect 206799 69900 210528 69902
rect 206799 69897 206865 69900
rect 144015 69812 144081 69815
rect 140802 69810 144081 69812
rect 140802 69754 144020 69810
rect 144076 69754 144081 69810
rect 140802 69752 144081 69754
rect 144015 69749 144081 69752
rect 204975 69516 205041 69519
rect 204975 69514 210528 69516
rect 204975 69458 204980 69514
rect 205036 69458 210528 69514
rect 204975 69456 210528 69458
rect 204975 69453 205041 69456
rect 146319 69072 146385 69075
rect 140832 69070 146385 69072
rect 140832 69014 146324 69070
rect 146380 69014 146385 69070
rect 140832 69012 146385 69014
rect 146319 69009 146385 69012
rect 204495 68924 204561 68927
rect 204495 68922 210528 68924
rect 204495 68866 204500 68922
rect 204556 68866 210528 68922
rect 204495 68864 210528 68866
rect 204495 68861 204561 68864
rect 206415 68332 206481 68335
rect 206415 68330 210528 68332
rect 206415 68274 206420 68330
rect 206476 68274 210528 68330
rect 206415 68272 210528 68274
rect 206415 68269 206481 68272
rect 140802 67444 140862 67932
rect 204591 67888 204657 67891
rect 204591 67886 210528 67888
rect 204591 67830 204596 67886
rect 204652 67830 210528 67886
rect 204591 67828 210528 67830
rect 204591 67825 204657 67828
rect 144111 67444 144177 67447
rect 140802 67442 144177 67444
rect 140802 67386 144116 67442
rect 144172 67386 144177 67442
rect 140802 67384 144177 67386
rect 144111 67381 144177 67384
rect 204111 67296 204177 67299
rect 204111 67294 210528 67296
rect 204111 67238 204116 67294
rect 204172 67238 210528 67294
rect 204111 67236 210528 67238
rect 204111 67233 204177 67236
rect 140802 66408 140862 66748
rect 206511 66704 206577 66707
rect 206511 66702 210528 66704
rect 206511 66646 206516 66702
rect 206572 66646 210528 66702
rect 206511 66644 210528 66646
rect 206511 66641 206577 66644
rect 146799 66408 146865 66411
rect 140802 66406 146865 66408
rect 140802 66350 146804 66406
rect 146860 66350 146865 66406
rect 140802 66348 146865 66350
rect 146799 66345 146865 66348
rect 144783 66262 144849 66263
rect 144783 66260 144832 66262
rect 144740 66258 144832 66260
rect 144740 66202 144788 66258
rect 144740 66200 144832 66202
rect 144783 66198 144832 66200
rect 144896 66198 144902 66262
rect 204495 66260 204561 66263
rect 204495 66258 210528 66260
rect 204495 66202 204500 66258
rect 204556 66202 210528 66258
rect 204495 66200 210528 66202
rect 144783 66197 144849 66198
rect 204495 66197 204561 66200
rect 206319 65668 206385 65671
rect 206319 65666 210528 65668
rect 206319 65610 206324 65666
rect 206380 65610 210528 65666
rect 206319 65608 210528 65610
rect 206319 65605 206385 65608
rect 144975 65520 145041 65523
rect 140832 65518 145041 65520
rect 140832 65462 144980 65518
rect 145036 65462 145041 65518
rect 140832 65460 145041 65462
rect 144975 65457 145041 65460
rect 205455 65076 205521 65079
rect 205455 65074 210528 65076
rect 205455 65018 205460 65074
rect 205516 65018 210528 65074
rect 205455 65016 210528 65018
rect 205455 65013 205521 65016
rect 144303 64632 144369 64635
rect 140802 64630 144369 64632
rect 140802 64574 144308 64630
rect 144364 64574 144369 64630
rect 140802 64572 144369 64574
rect 140802 64334 140862 64572
rect 144303 64569 144369 64572
rect 144826 64570 144832 64634
rect 144896 64632 144902 64634
rect 144975 64632 145041 64635
rect 144896 64630 145041 64632
rect 144896 64574 144980 64630
rect 145036 64574 145041 64630
rect 144896 64572 145041 64574
rect 144896 64570 144902 64572
rect 144975 64569 145041 64572
rect 204495 64632 204561 64635
rect 204495 64630 210528 64632
rect 204495 64574 204500 64630
rect 204556 64574 210528 64630
rect 204495 64572 210528 64574
rect 204495 64569 204561 64572
rect 204591 64040 204657 64043
rect 204591 64038 210528 64040
rect 204591 63982 204596 64038
rect 204652 63982 210528 64038
rect 204591 63980 210528 63982
rect 204591 63977 204657 63980
rect 204495 63448 204561 63451
rect 204495 63446 210528 63448
rect 204495 63390 204500 63446
rect 204556 63390 210528 63446
rect 204495 63388 210528 63390
rect 204495 63385 204561 63388
rect 140802 62856 140862 63048
rect 204591 63004 204657 63007
rect 204591 63002 210528 63004
rect 204591 62946 204596 63002
rect 204652 62946 210528 63002
rect 204591 62944 210528 62946
rect 204591 62941 204657 62944
rect 144015 62856 144081 62859
rect 140802 62854 144081 62856
rect 140802 62798 144020 62854
rect 144076 62798 144081 62854
rect 140802 62796 144081 62798
rect 144015 62793 144081 62796
rect 146895 62412 146961 62415
rect 140802 62410 146961 62412
rect 140802 62354 146900 62410
rect 146956 62354 146961 62410
rect 140802 62352 146961 62354
rect 140802 61864 140862 62352
rect 146895 62349 146961 62352
rect 204687 62412 204753 62415
rect 204687 62410 210528 62412
rect 204687 62354 204692 62410
rect 204748 62354 210528 62410
rect 204687 62352 210528 62354
rect 204687 62349 204753 62352
rect 204879 61820 204945 61823
rect 204879 61818 210528 61820
rect 204879 61762 204884 61818
rect 204940 61762 210528 61818
rect 204879 61760 210528 61762
rect 204879 61757 204945 61760
rect 204783 61376 204849 61379
rect 204783 61374 210528 61376
rect 204783 61318 204788 61374
rect 204844 61318 210528 61374
rect 204783 61316 210528 61318
rect 204783 61313 204849 61316
rect 146895 60784 146961 60787
rect 140832 60782 146961 60784
rect 140832 60726 146900 60782
rect 146956 60726 146961 60782
rect 140832 60724 146961 60726
rect 146895 60721 146961 60724
rect 204495 60784 204561 60787
rect 204495 60782 210528 60784
rect 204495 60726 204500 60782
rect 204556 60726 210528 60782
rect 204495 60724 210528 60726
rect 204495 60721 204561 60724
rect 204495 60192 204561 60195
rect 204495 60190 210528 60192
rect 204495 60134 204500 60190
rect 204556 60134 210528 60190
rect 204495 60132 210528 60134
rect 204495 60129 204561 60132
rect 206799 60044 206865 60047
rect 206799 60042 210558 60044
rect 206799 59986 206804 60042
rect 206860 59986 210558 60042
rect 206799 59984 210558 59986
rect 206799 59981 206865 59984
rect 210498 59644 210558 59984
rect 144015 59600 144081 59603
rect 140832 59598 144081 59600
rect 140832 59542 144020 59598
rect 144076 59542 144081 59598
rect 140832 59540 144081 59542
rect 144015 59537 144081 59540
rect 204591 59156 204657 59159
rect 204591 59154 210528 59156
rect 204591 59098 204596 59154
rect 204652 59098 210528 59154
rect 204591 59096 210528 59098
rect 204591 59093 204657 59096
rect 144015 58712 144081 58715
rect 140802 58710 144081 58712
rect 140802 58654 144020 58710
rect 144076 58654 144081 58710
rect 140802 58652 144081 58654
rect 140802 58322 140862 58652
rect 144015 58649 144081 58652
rect 211074 58270 211134 58534
rect 211066 58206 211072 58270
rect 211136 58206 211142 58270
rect 207279 57676 207345 57679
rect 210498 57676 210558 58016
rect 207279 57674 210558 57676
rect 207279 57618 207284 57674
rect 207340 57618 210558 57674
rect 207279 57616 210558 57618
rect 207279 57613 207345 57616
rect 209199 57232 209265 57235
rect 210498 57232 210558 57498
rect 209199 57230 210558 57232
rect 209199 57174 209204 57230
rect 209260 57174 210558 57230
rect 209199 57172 210558 57174
rect 209199 57169 209265 57172
rect 144015 57084 144081 57087
rect 140832 57082 144081 57084
rect 140832 57026 144020 57082
rect 144076 57026 144081 57082
rect 140832 57024 144081 57026
rect 144015 57021 144081 57024
rect 209295 56640 209361 56643
rect 210498 56640 210558 56906
rect 209295 56638 210558 56640
rect 209295 56582 209300 56638
rect 209356 56582 210558 56638
rect 209295 56580 210558 56582
rect 209295 56577 209361 56580
rect 144015 56196 144081 56199
rect 140802 56194 144081 56196
rect 140802 56138 144020 56194
rect 144076 56138 144081 56194
rect 140802 56136 144081 56138
rect 140802 55874 140862 56136
rect 144015 56133 144081 56136
rect 209967 56048 210033 56051
rect 210498 56048 210558 56388
rect 209967 56046 210558 56048
rect 209967 55990 209972 56046
rect 210028 55990 210558 56046
rect 209967 55988 210558 55990
rect 209967 55985 210033 55988
rect 206895 55900 206961 55903
rect 206895 55898 210528 55900
rect 206895 55842 206900 55898
rect 206956 55842 210528 55898
rect 206895 55840 210528 55842
rect 206895 55837 206961 55840
rect 210255 55012 210321 55015
rect 210498 55012 210558 55278
rect 210255 55010 210558 55012
rect 210255 54954 210260 55010
rect 210316 54954 210558 55010
rect 210255 54952 210558 54954
rect 210255 54949 210321 54952
rect 209967 54790 210033 54793
rect 209967 54788 210528 54790
rect 209967 54732 209972 54788
rect 210028 54732 210528 54788
rect 209967 54730 210528 54732
rect 209967 54727 210033 54730
rect 144015 54716 144081 54719
rect 140832 54714 144081 54716
rect 140832 54658 144020 54714
rect 144076 54658 144081 54714
rect 140832 54656 144081 54658
rect 144015 54653 144081 54656
rect 210874 54210 210880 54274
rect 210944 54272 210950 54274
rect 212367 54272 212433 54275
rect 210944 54270 212433 54272
rect 210944 54214 212372 54270
rect 212428 54214 212433 54270
rect 210944 54212 212433 54214
rect 210944 54210 210950 54212
rect 212367 54209 212433 54212
rect 212602 54210 212608 54274
rect 212672 54272 212678 54274
rect 214383 54272 214449 54275
rect 212672 54270 214449 54272
rect 212672 54214 214388 54270
rect 214444 54214 214449 54270
rect 212672 54212 214449 54214
rect 212672 54210 212678 54212
rect 214383 54209 214449 54212
rect 211258 54062 211264 54126
rect 211328 54124 211334 54126
rect 214767 54124 214833 54127
rect 211328 54122 214833 54124
rect 211328 54066 214772 54122
rect 214828 54066 214833 54122
rect 211328 54064 214833 54066
rect 211328 54062 211334 54064
rect 214767 54061 214833 54064
rect 212218 53914 212224 53978
rect 212288 53976 212294 53978
rect 216591 53976 216657 53979
rect 212288 53974 216657 53976
rect 212288 53918 216596 53974
rect 216652 53918 216657 53974
rect 212288 53916 216657 53918
rect 212288 53914 212294 53916
rect 216591 53913 216657 53916
rect 144015 53828 144081 53831
rect 140802 53826 144081 53828
rect 140802 53770 144020 53826
rect 144076 53770 144081 53826
rect 140802 53768 144081 53770
rect 140802 53576 140862 53768
rect 144015 53765 144081 53768
rect 210682 53766 210688 53830
rect 210752 53828 210758 53830
rect 216975 53828 217041 53831
rect 210752 53826 217041 53828
rect 210752 53770 216980 53826
rect 217036 53770 217041 53826
rect 210752 53768 217041 53770
rect 210752 53766 210758 53768
rect 216975 53765 217041 53768
rect 211834 53618 211840 53682
rect 211904 53680 211910 53682
rect 211904 53620 215982 53680
rect 211904 53618 211910 53620
rect 215922 53535 215982 53620
rect 213039 53534 213105 53535
rect 212986 53470 212992 53534
rect 213056 53532 213105 53534
rect 213056 53530 213148 53532
rect 213100 53474 213148 53530
rect 213056 53472 213148 53474
rect 215919 53530 215985 53535
rect 215919 53474 215924 53530
rect 215980 53474 215985 53530
rect 213056 53470 213105 53472
rect 213039 53469 213105 53470
rect 215919 53469 215985 53474
rect 216783 53532 216849 53535
rect 219999 53532 220065 53535
rect 216783 53530 220065 53532
rect 216783 53474 216788 53530
rect 216844 53474 220004 53530
rect 220060 53474 220065 53530
rect 216783 53472 220065 53474
rect 216783 53469 216849 53472
rect 219999 53469 220065 53472
rect 212410 53322 212416 53386
rect 212480 53384 212486 53386
rect 215247 53384 215313 53387
rect 212480 53382 215313 53384
rect 212480 53326 215252 53382
rect 215308 53326 215313 53382
rect 212480 53324 215313 53326
rect 212480 53322 212486 53324
rect 215247 53321 215313 53324
rect 207087 53236 207153 53239
rect 220335 53236 220401 53239
rect 207087 53234 220401 53236
rect 207087 53178 207092 53234
rect 207148 53178 220340 53234
rect 220396 53178 220401 53234
rect 207087 53176 220401 53178
rect 207087 53173 207153 53176
rect 220335 53173 220401 53176
rect 211066 53026 211072 53090
rect 211136 53088 211142 53090
rect 216015 53088 216081 53091
rect 211136 53086 216081 53088
rect 211136 53030 216020 53086
rect 216076 53030 216081 53086
rect 211136 53028 216081 53030
rect 211136 53026 211142 53028
rect 216015 53025 216081 53028
rect 161295 52200 161361 52203
rect 181359 52200 181425 52203
rect 161295 52198 181425 52200
rect 161295 52142 161300 52198
rect 161356 52142 181364 52198
rect 181420 52142 181425 52198
rect 161295 52140 181425 52142
rect 161295 52137 161361 52140
rect 181359 52137 181425 52140
rect 222543 52200 222609 52203
rect 637882 52200 637888 52202
rect 222543 52198 637888 52200
rect 222543 52142 222548 52198
rect 222604 52142 637888 52198
rect 222543 52140 637888 52142
rect 222543 52137 222609 52140
rect 637882 52138 637888 52140
rect 637952 52138 637958 52202
rect 212655 52052 212721 52055
rect 637498 52052 637504 52054
rect 212655 52050 637504 52052
rect 212655 51994 212660 52050
rect 212716 51994 637504 52050
rect 212655 51992 637504 51994
rect 212655 51989 212721 51992
rect 637498 51990 637504 51992
rect 637568 51990 637574 52054
rect 211887 51904 211953 51907
rect 637690 51904 637696 51906
rect 211887 51902 637696 51904
rect 211887 51846 211892 51902
rect 211948 51846 637696 51902
rect 211887 51844 637696 51846
rect 211887 51841 211953 51844
rect 637690 51842 637696 51844
rect 637760 51842 637766 51906
rect 221871 51756 221937 51759
rect 637306 51756 637312 51758
rect 221871 51754 637312 51756
rect 221871 51698 221876 51754
rect 221932 51698 637312 51754
rect 221871 51696 637312 51698
rect 221871 51693 221937 51696
rect 637306 51694 637312 51696
rect 637376 51694 637382 51758
rect 223311 51608 223377 51611
rect 637114 51608 637120 51610
rect 223311 51606 637120 51608
rect 223311 51550 223316 51606
rect 223372 51550 637120 51606
rect 223311 51548 637120 51550
rect 223311 51545 223377 51548
rect 637114 51546 637120 51548
rect 637184 51546 637190 51610
rect 145402 51398 145408 51462
rect 145472 51460 145478 51462
rect 243375 51460 243441 51463
rect 145472 51458 243441 51460
rect 145472 51402 243380 51458
rect 243436 51402 243441 51458
rect 145472 51400 243441 51402
rect 145472 51398 145478 51400
rect 243375 51397 243441 51400
rect 145594 51250 145600 51314
rect 145664 51312 145670 51314
rect 238191 51312 238257 51315
rect 145664 51310 238257 51312
rect 145664 51254 238196 51310
rect 238252 51254 238257 51310
rect 145664 51252 238257 51254
rect 145664 51250 145670 51252
rect 238191 51249 238257 51252
rect 229647 50424 229713 50427
rect 636922 50424 636928 50426
rect 229647 50422 636928 50424
rect 229647 50366 229652 50422
rect 229708 50366 636928 50422
rect 229647 50364 636928 50366
rect 229647 50361 229713 50364
rect 636922 50362 636928 50364
rect 636992 50362 636998 50426
rect 209487 48944 209553 48947
rect 220719 48944 220785 48947
rect 209487 48942 220785 48944
rect 209487 48886 209492 48942
rect 209548 48886 220724 48942
rect 220780 48886 220785 48942
rect 209487 48884 220785 48886
rect 209487 48881 209553 48884
rect 220719 48881 220785 48884
rect 171279 48648 171345 48651
rect 242031 48648 242097 48651
rect 171279 48646 242097 48648
rect 171279 48590 171284 48646
rect 171340 48590 242036 48646
rect 242092 48590 242097 48646
rect 171279 48588 242097 48590
rect 171279 48585 171345 48588
rect 242031 48585 242097 48588
rect 174159 48500 174225 48503
rect 242991 48500 243057 48503
rect 174159 48498 243057 48500
rect 174159 48442 174164 48498
rect 174220 48442 242996 48498
rect 243052 48442 243057 48498
rect 174159 48440 243057 48442
rect 174159 48437 174225 48440
rect 242991 48437 243057 48440
rect 177039 48352 177105 48355
rect 243759 48352 243825 48355
rect 177039 48350 243825 48352
rect 177039 48294 177044 48350
rect 177100 48294 243764 48350
rect 243820 48294 243825 48350
rect 177039 48292 243825 48294
rect 177039 48289 177105 48292
rect 243759 48289 243825 48292
rect 165519 48204 165585 48207
rect 241935 48204 242001 48207
rect 165519 48202 242001 48204
rect 165519 48146 165524 48202
rect 165580 48146 241940 48202
rect 241996 48146 242001 48202
rect 165519 48144 242001 48146
rect 165519 48141 165585 48144
rect 241935 48141 242001 48144
rect 168399 47908 168465 47911
rect 242607 47908 242673 47911
rect 168399 47906 242673 47908
rect 168399 47850 168404 47906
rect 168460 47850 242612 47906
rect 242668 47850 242673 47906
rect 168399 47848 242673 47850
rect 168399 47845 168465 47848
rect 242607 47845 242673 47848
rect 466575 46132 466641 46135
rect 471034 46132 471040 46134
rect 466575 46130 471040 46132
rect 466575 46074 466580 46130
rect 466636 46074 471040 46130
rect 466575 46072 471040 46074
rect 466575 46069 466641 46072
rect 471034 46070 471040 46072
rect 471104 46070 471110 46134
rect 212079 45096 212145 45099
rect 302458 45096 302464 45098
rect 212079 45094 302464 45096
rect 212079 45038 212084 45094
rect 212140 45038 302464 45094
rect 212079 45036 302464 45038
rect 212079 45033 212145 45036
rect 302458 45034 302464 45036
rect 302528 45034 302534 45098
rect 212847 44948 212913 44951
rect 414778 44948 414784 44950
rect 212847 44946 414784 44948
rect 212847 44890 212852 44946
rect 212908 44890 414784 44946
rect 212847 44888 414784 44890
rect 212847 44885 212913 44888
rect 414778 44886 414784 44888
rect 414848 44886 414854 44950
rect 302511 43322 302577 43323
rect 302458 43320 302464 43322
rect 302420 43260 302464 43320
rect 302528 43318 302577 43322
rect 302572 43262 302577 43318
rect 302458 43258 302464 43260
rect 302528 43258 302577 43262
rect 414778 43258 414784 43322
rect 414848 43320 414854 43322
rect 416559 43320 416625 43323
rect 414848 43318 416625 43320
rect 414848 43262 416564 43318
rect 416620 43262 416625 43318
rect 414848 43260 416625 43262
rect 414848 43258 414854 43260
rect 302511 43257 302577 43258
rect 416559 43257 416625 43260
rect 517839 43320 517905 43323
rect 520623 43320 520689 43323
rect 517839 43318 520689 43320
rect 517839 43262 517844 43318
rect 517900 43262 520628 43318
rect 520684 43262 520689 43318
rect 517839 43260 520689 43262
rect 517839 43257 517905 43260
rect 520623 43257 520689 43260
rect 461103 43172 461169 43175
rect 465615 43172 465681 43175
rect 461103 43170 465681 43172
rect 461103 43114 461108 43170
rect 461164 43114 465620 43170
rect 465676 43114 465681 43170
rect 461103 43112 465681 43114
rect 461103 43109 461169 43112
rect 465615 43109 465681 43112
rect 302319 42136 302385 42139
rect 306735 42136 306801 42139
rect 471087 42138 471153 42139
rect 302319 42134 306801 42136
rect 302319 42078 302324 42134
rect 302380 42078 306740 42134
rect 306796 42078 306801 42134
rect 302319 42076 306801 42078
rect 302319 42073 302385 42076
rect 306735 42073 306801 42076
rect 471034 42074 471040 42138
rect 471104 42136 471153 42138
rect 526959 42136 527025 42139
rect 528975 42136 529041 42139
rect 471104 42134 471196 42136
rect 471148 42078 471196 42134
rect 471104 42076 471196 42078
rect 526959 42134 529041 42136
rect 526959 42078 526964 42134
rect 527020 42078 528980 42134
rect 529036 42078 529041 42134
rect 526959 42076 529041 42078
rect 471104 42074 471153 42076
rect 471087 42073 471153 42074
rect 526959 42073 527025 42076
rect 528975 42073 529041 42076
rect 187599 41840 187665 41843
rect 189946 41840 189952 41842
rect 187599 41838 189952 41840
rect 187599 41782 187604 41838
rect 187660 41782 189952 41838
rect 187599 41780 189952 41782
rect 187599 41777 187665 41780
rect 189946 41778 189952 41780
rect 190016 41778 190022 41842
rect 194319 41840 194385 41843
rect 194938 41840 194944 41842
rect 194319 41838 194944 41840
rect 194319 41782 194324 41838
rect 194380 41782 194944 41838
rect 194319 41780 194944 41782
rect 194319 41777 194385 41780
rect 194938 41778 194944 41780
rect 195008 41778 195014 41842
rect 360058 41778 360064 41842
rect 360128 41840 360134 41842
rect 361455 41840 361521 41843
rect 360128 41838 361521 41840
rect 360128 41782 361460 41838
rect 361516 41782 361521 41838
rect 360128 41780 361521 41782
rect 360128 41778 360134 41780
rect 361455 41777 361521 41780
rect 362938 41778 362944 41842
rect 363008 41840 363014 41842
rect 364623 41840 364689 41843
rect 363008 41838 364689 41840
rect 363008 41782 364628 41838
rect 364684 41782 364689 41838
rect 363008 41780 364689 41782
rect 363008 41778 363014 41780
rect 364623 41777 364689 41780
rect 459322 41778 459328 41842
rect 459392 41840 459398 41842
rect 463695 41840 463761 41843
rect 459392 41838 463761 41840
rect 459392 41782 463700 41838
rect 463756 41782 463761 41838
rect 459392 41780 463761 41782
rect 459392 41778 459398 41780
rect 463695 41777 463761 41780
rect 328047 40952 328113 40955
rect 360058 40952 360064 40954
rect 328047 40950 360064 40952
rect 328047 40894 328052 40950
rect 328108 40894 360064 40950
rect 328047 40892 360064 40894
rect 328047 40889 328113 40892
rect 360058 40890 360064 40892
rect 360128 40890 360134 40954
rect 189946 40742 189952 40806
rect 190016 40804 190022 40806
rect 210735 40804 210801 40807
rect 190016 40802 210801 40804
rect 190016 40746 210740 40802
rect 210796 40746 210801 40802
rect 190016 40744 210801 40746
rect 190016 40742 190022 40744
rect 210735 40741 210801 40744
rect 327279 40804 327345 40807
rect 362938 40804 362944 40806
rect 327279 40802 362944 40804
rect 327279 40746 327284 40802
rect 327340 40746 362944 40802
rect 327279 40744 362944 40746
rect 327279 40741 327345 40744
rect 362938 40742 362944 40744
rect 363008 40742 363014 40806
rect 194938 40594 194944 40658
rect 195008 40656 195014 40658
rect 640719 40656 640785 40659
rect 195008 40654 640785 40656
rect 195008 40598 640724 40654
rect 640780 40598 640785 40654
rect 195008 40596 640785 40598
rect 195008 40594 195014 40596
rect 640719 40593 640785 40596
rect 454959 40360 455025 40363
rect 455098 40360 455104 40362
rect 454959 40358 455104 40360
rect 454959 40302 454964 40358
rect 455020 40302 455104 40358
rect 454959 40300 455104 40302
rect 454959 40297 455025 40300
rect 455098 40298 455104 40300
rect 455168 40298 455174 40362
rect 136527 40212 136593 40215
rect 136527 40210 141822 40212
rect 136527 40154 136532 40210
rect 136588 40154 141822 40210
rect 136527 40152 141822 40154
rect 136527 40149 136593 40152
rect 141762 39886 141822 40152
<< via3 >>
rect 83392 993626 83456 993630
rect 83392 993570 83444 993626
rect 83444 993570 83456 993626
rect 83392 993566 83456 993570
rect 83392 992086 83456 992150
rect 40960 968702 41024 968766
rect 675328 967370 675392 967434
rect 40576 967074 40640 967138
rect 676672 966334 676736 966398
rect 675712 965802 675776 965806
rect 675712 965746 675724 965802
rect 675724 965746 675776 965802
rect 675712 965742 675776 965746
rect 40768 965002 40832 965066
rect 675136 964914 675200 964918
rect 675136 964858 675188 964914
rect 675188 964858 675200 964914
rect 675136 964854 675200 964858
rect 40384 963966 40448 964030
rect 41536 963226 41600 963290
rect 676480 963226 676544 963290
rect 42304 962782 42368 962846
rect 674368 962486 674432 962550
rect 42112 962250 42176 962254
rect 42112 962194 42124 962250
rect 42124 962194 42176 962250
rect 42112 962190 42176 962194
rect 43072 962190 43136 962254
rect 674560 962190 674624 962254
rect 42880 962042 42944 962106
rect 674176 961450 674240 961514
rect 675328 961362 675392 961366
rect 675328 961306 675380 961362
rect 675380 961306 675392 961362
rect 675328 961302 675392 961306
rect 675520 960178 675584 960182
rect 675520 960122 675532 960178
rect 675532 960122 675584 960178
rect 675520 960118 675584 960122
rect 42688 959526 42752 959590
rect 41728 959142 41792 959146
rect 41728 959086 41780 959142
rect 41780 959086 41792 959142
rect 41728 959082 41792 959086
rect 676096 959082 676160 959146
rect 41920 958402 41984 958406
rect 41920 958346 41972 958402
rect 41972 958346 41984 958402
rect 41920 958342 41984 958346
rect 42496 957750 42560 957814
rect 674752 957750 674816 957814
rect 41152 956566 41216 956630
rect 674944 955974 675008 956038
rect 677056 953458 677120 953522
rect 676864 953310 676928 953374
rect 41152 944430 41216 944494
rect 40576 943690 40640 943754
rect 42496 941618 42560 941682
rect 42112 941174 42176 941238
rect 675136 940878 675200 940942
rect 40960 940582 41024 940646
rect 676672 939250 676736 939314
rect 41920 938806 41984 938870
rect 41728 938066 41792 938130
rect 676480 938066 676544 938130
rect 40768 937326 40832 937390
rect 676096 937326 676160 937390
rect 41536 936438 41600 936502
rect 675712 935846 675776 935910
rect 42688 935254 42752 935318
rect 42304 934958 42368 935022
rect 674368 934662 674432 934726
rect 674560 934514 674624 934578
rect 40384 934070 40448 934134
rect 674944 933330 675008 933394
rect 674752 932886 674816 932950
rect 674176 931554 674240 931618
rect 677056 931406 677120 931470
rect 676864 930222 676928 930286
rect 676096 876942 676160 877006
rect 673984 876498 674048 876562
rect 674752 875906 674816 875970
rect 675328 875758 675392 875822
rect 675520 875610 675584 875674
rect 674560 873982 674624 874046
rect 674176 873390 674240 873454
rect 674944 869838 675008 869902
rect 676672 864658 676736 864722
rect 675328 862942 675392 862946
rect 675328 862886 675380 862942
rect 675380 862886 675392 862942
rect 675328 862882 675392 862886
rect 41344 818630 41408 818694
rect 41536 802202 41600 802266
rect 42688 802202 42752 802266
rect 41152 802054 41216 802118
rect 41728 801906 41792 801970
rect 42304 800426 42368 800490
rect 41920 800278 41984 800342
rect 42112 800338 42176 800342
rect 42112 800282 42124 800338
rect 42124 800282 42176 800338
rect 42112 800278 42176 800282
rect 42496 799746 42560 799750
rect 42496 799690 42508 799746
rect 42508 799690 42560 799746
rect 42496 799686 42560 799690
rect 42688 798354 42752 798418
rect 41920 794270 41984 794274
rect 41920 794214 41932 794270
rect 41932 794214 41984 794270
rect 41920 794210 41984 794214
rect 42112 793826 42176 793830
rect 42112 793770 42124 793826
rect 42124 793770 42176 793826
rect 42112 793766 42176 793770
rect 42496 792494 42560 792498
rect 42496 792438 42508 792494
rect 42508 792438 42560 792494
rect 42496 792434 42560 792438
rect 42304 792286 42368 792350
rect 41536 791842 41600 791906
rect 42112 791694 42176 791758
rect 42112 791162 42176 791166
rect 42112 791106 42124 791162
rect 42124 791106 42176 791162
rect 42112 791102 42176 791106
rect 43072 791102 43136 791166
rect 41536 790954 41600 791018
rect 42880 790954 42944 791018
rect 41728 790510 41792 790574
rect 42304 788586 42368 788650
rect 675712 788054 675776 788058
rect 675712 787998 675724 788054
rect 675724 787998 675776 788054
rect 675712 787994 675776 787998
rect 675520 787166 675584 787170
rect 675520 787110 675532 787166
rect 675532 787110 675584 787166
rect 675520 787106 675584 787110
rect 676480 786662 676544 786726
rect 675904 784738 675968 784802
rect 674368 780594 674432 780658
rect 676864 779114 676928 779178
rect 677056 777486 677120 777550
rect 677056 777338 677120 777402
rect 41152 776746 41216 776810
rect 41536 775858 41600 775922
rect 676288 775414 676352 775478
rect 41344 775118 41408 775182
rect 675136 773638 675200 773702
rect 677824 773046 677888 773110
rect 42496 764018 42560 764082
rect 674752 762390 674816 762454
rect 676672 761650 676736 761714
rect 42880 760466 42944 760530
rect 676096 760466 676160 760530
rect 41152 760170 41216 760234
rect 674560 760022 674624 760086
rect 674944 759134 675008 759198
rect 40768 758690 40832 758754
rect 675328 758542 675392 758606
rect 42688 758394 42752 758458
rect 43072 757358 43136 757422
rect 40960 757210 41024 757274
rect 42112 757210 42176 757274
rect 41728 757122 41792 757126
rect 41728 757066 41780 757122
rect 41780 757066 41792 757122
rect 41728 757062 41792 757066
rect 42112 757122 42176 757126
rect 42112 757066 42124 757122
rect 42124 757066 42176 757122
rect 42112 757062 42176 757066
rect 673984 757062 674048 757126
rect 674176 756322 674240 756386
rect 677824 755286 677888 755350
rect 677248 754398 677312 754462
rect 42112 753126 42176 753130
rect 42112 753070 42124 753126
rect 42124 753070 42176 753126
rect 42112 753066 42176 753070
rect 42496 751734 42560 751798
rect 43072 751734 43136 751798
rect 42688 750994 42752 751058
rect 40960 748626 41024 748690
rect 41920 748626 41984 748690
rect 41728 747502 41792 747506
rect 41728 747446 41780 747502
rect 41780 747446 41792 747502
rect 41728 747442 41792 747446
rect 41728 747294 41792 747358
rect 42112 747294 42176 747358
rect 40768 747146 40832 747210
rect 41152 746702 41216 746766
rect 42880 745962 42944 746026
rect 674560 743150 674624 743214
rect 676672 742410 676736 742474
rect 676096 741670 676160 741734
rect 674944 740338 675008 740402
rect 674752 739302 674816 739366
rect 675328 738622 675392 738626
rect 675328 738566 675380 738622
rect 675380 738566 675392 738622
rect 675328 738562 675392 738566
rect 41536 733826 41600 733890
rect 41344 733086 41408 733150
rect 42112 732198 42176 732262
rect 677056 731754 677120 731818
rect 43072 729534 43136 729598
rect 677824 728054 677888 728118
rect 677056 727906 677120 727970
rect 41152 726278 41216 726342
rect 42112 725538 42176 725602
rect 43456 725538 43520 725602
rect 41920 722430 41984 722494
rect 42496 722430 42560 722494
rect 43264 721394 43328 721458
rect 673984 717014 674048 717018
rect 676480 717102 676544 717166
rect 673984 716958 673996 717014
rect 673996 716958 674048 717014
rect 673984 716954 674048 716958
rect 676288 716658 676352 716722
rect 675712 715770 675776 715834
rect 675904 715030 675968 715094
rect 41920 714290 41984 714354
rect 41344 714202 41408 714206
rect 41344 714146 41396 714202
rect 41396 714146 41408 714202
rect 41344 714142 41408 714146
rect 42880 714142 42944 714206
rect 41728 713906 41792 713910
rect 41728 713850 41780 713906
rect 41780 713850 41792 713906
rect 41728 713846 41792 713850
rect 42688 713846 42752 713910
rect 674368 713698 674432 713762
rect 675136 713550 675200 713614
rect 675520 712662 675584 712726
rect 41344 711034 41408 711098
rect 677824 710294 677888 710358
rect 42688 709702 42752 709766
rect 676864 709406 676928 709470
rect 43264 708518 43328 708582
rect 41920 707986 41984 707990
rect 41920 707930 41932 707986
rect 41932 707930 41984 707986
rect 41920 707926 41984 707930
rect 42880 707926 42944 707990
rect 41728 706802 41792 706806
rect 41728 706746 41780 706802
rect 41780 706746 41792 706802
rect 41728 706742 41792 706746
rect 43456 705854 43520 705918
rect 42304 705706 42368 705770
rect 41152 705410 41216 705474
rect 42112 704730 42176 704734
rect 42112 704674 42124 704730
rect 42124 704674 42176 704730
rect 42112 704670 42176 704674
rect 42496 704670 42560 704734
rect 41728 704138 41792 704142
rect 41728 704082 41780 704138
rect 41780 704082 41792 704138
rect 41728 704078 41792 704082
rect 43072 702806 43136 702810
rect 43072 702750 43084 702806
rect 43084 702750 43136 702806
rect 43072 702746 43136 702750
rect 675520 697922 675584 697926
rect 675520 697866 675532 697922
rect 675532 697866 675584 697922
rect 675520 697862 675584 697866
rect 676480 697270 676544 697334
rect 675904 697122 675968 697186
rect 675712 694814 675776 694818
rect 675712 694758 675724 694814
rect 675724 694758 675776 694814
rect 675712 694754 675776 694758
rect 674176 694310 674240 694374
rect 674368 693422 674432 693486
rect 676288 691646 676352 691710
rect 41536 690314 41600 690378
rect 42112 689574 42176 689638
rect 675136 689130 675200 689194
rect 42304 688686 42368 688750
rect 676864 687502 676928 687566
rect 41920 675366 41984 675430
rect 42880 675366 42944 675430
rect 40768 673886 40832 673950
rect 673984 672998 674048 673062
rect 40576 672554 40640 672618
rect 676096 672258 676160 672322
rect 41728 670926 41792 670990
rect 42688 670926 42752 670990
rect 43072 670986 43136 670990
rect 43072 670930 43124 670986
rect 43124 670930 43136 670986
rect 43072 670926 43136 670930
rect 41920 670838 41984 670842
rect 41920 670782 41972 670838
rect 41972 670782 41984 670838
rect 41920 670778 41984 670782
rect 42496 670778 42560 670842
rect 674560 670482 674624 670546
rect 674944 669742 675008 669806
rect 676672 667522 676736 667586
rect 674752 666634 674816 666698
rect 675328 665894 675392 665958
rect 43072 665302 43136 665366
rect 677056 663526 677120 663590
rect 42688 663378 42752 663442
rect 42496 662846 42560 662850
rect 42496 662790 42508 662846
rect 42508 662790 42560 662846
rect 42496 662786 42560 662790
rect 40768 662342 40832 662406
rect 42496 661454 42560 661518
rect 41152 660714 41216 660778
rect 41728 660330 41792 660334
rect 41728 660274 41780 660330
rect 41780 660274 41792 660330
rect 41728 660270 41792 660274
rect 41728 660122 41792 660186
rect 41920 659146 41984 659150
rect 41920 659090 41932 659146
rect 41932 659090 41984 659146
rect 41920 659086 41984 659090
rect 41920 658938 41984 659002
rect 42496 658938 42560 659002
rect 40576 656570 40640 656634
rect 676288 653610 676352 653674
rect 675328 652634 675392 652638
rect 675328 652578 675380 652634
rect 675380 652578 675392 652634
rect 675328 652574 675392 652578
rect 674560 652130 674624 652194
rect 674944 651390 675008 651454
rect 676672 649762 676736 649826
rect 674752 648874 674816 648938
rect 42112 647394 42176 647458
rect 42304 646654 42368 646718
rect 676096 645322 676160 645386
rect 673984 640290 674048 640354
rect 675904 639846 675968 639910
rect 675712 639402 675776 639466
rect 42688 638884 42752 638948
rect 675520 638662 675584 638726
rect 675520 638574 675584 638578
rect 675520 638518 675532 638574
rect 675532 638518 675584 638574
rect 675520 638514 675584 638518
rect 675712 630878 675776 630882
rect 675712 630822 675764 630878
rect 675764 630822 675776 630878
rect 675712 630818 675776 630822
rect 675904 630818 675968 630882
rect 675712 630434 675776 630438
rect 675712 630378 675764 630434
rect 675764 630378 675776 630434
rect 675712 630374 675776 630378
rect 40768 628154 40832 628218
rect 40576 627858 40640 627922
rect 41344 627770 41408 627774
rect 41344 627714 41356 627770
rect 41356 627714 41408 627770
rect 41344 627710 41408 627714
rect 41728 627710 41792 627774
rect 41920 627562 41984 627626
rect 42112 627474 42176 627478
rect 42112 627418 42124 627474
rect 42124 627418 42176 627474
rect 42112 627414 42176 627418
rect 676288 627266 676352 627330
rect 675904 625638 675968 625702
rect 42688 625046 42752 625110
rect 42304 624898 42368 624962
rect 42496 624750 42560 624814
rect 675712 624750 675776 624814
rect 676480 622086 676544 622150
rect 42112 621702 42176 621706
rect 42112 621646 42124 621702
rect 42124 621646 42176 621702
rect 42112 621642 42176 621646
rect 674176 621050 674240 621114
rect 41920 620814 41984 620818
rect 41920 620758 41972 620814
rect 41972 620758 41984 620814
rect 41920 620754 41984 620758
rect 674368 620310 674432 620374
rect 675136 619126 675200 619190
rect 41536 618238 41600 618302
rect 41920 618150 41984 618154
rect 41920 618094 41972 618150
rect 41972 618094 41984 618150
rect 41920 618090 41984 618094
rect 42496 618090 42560 618154
rect 41728 617854 41792 617858
rect 41728 617798 41780 617854
rect 41780 617798 41792 617854
rect 41728 617794 41792 617798
rect 676864 617794 676928 617858
rect 41344 616462 41408 616526
rect 40768 613354 40832 613418
rect 673984 613354 674048 613418
rect 676288 613354 676352 613418
rect 40576 612762 40640 612826
rect 673984 607730 674048 607794
rect 674368 607138 674432 607202
rect 675712 606458 675776 606462
rect 675712 606402 675724 606458
rect 675724 606402 675776 606458
rect 675712 606398 675776 606402
rect 41920 604918 41984 604982
rect 42112 604770 42176 604834
rect 675136 604770 675200 604834
rect 674176 600182 674240 600246
rect 40960 599886 41024 599950
rect 40768 596778 40832 596842
rect 41152 594410 41216 594474
rect 43072 593670 43136 593734
rect 675904 593522 675968 593586
rect 676672 593522 676736 593586
rect 676864 593374 676928 593438
rect 41344 585974 41408 586038
rect 42112 585974 42176 586038
rect 42496 584790 42560 584854
rect 42304 584642 42368 584706
rect 42880 584642 42944 584706
rect 41728 584494 41792 584558
rect 41920 584406 41984 584410
rect 41920 584350 41932 584406
rect 41932 584350 41984 584406
rect 41920 584346 41984 584350
rect 42112 584258 42176 584262
rect 42112 584202 42124 584258
rect 42124 584202 42176 584258
rect 42112 584198 42176 584202
rect 42688 583754 42752 583818
rect 41920 582038 41984 582042
rect 41920 581982 41972 582038
rect 41972 581982 41984 582038
rect 41920 581978 41984 581982
rect 674944 581682 675008 581746
rect 43072 581386 43136 581450
rect 676480 581238 676544 581302
rect 675328 580350 675392 580414
rect 41152 580202 41216 580266
rect 675904 579610 675968 579674
rect 42688 578870 42752 578934
rect 674176 578870 674240 578934
rect 675904 578870 675968 578934
rect 676288 578722 676352 578786
rect 42880 578338 42944 578342
rect 42880 578282 42932 578338
rect 42932 578282 42944 578338
rect 42880 578278 42944 578282
rect 675520 578130 675584 578194
rect 42496 577538 42560 577602
rect 674560 577242 674624 577306
rect 41728 577006 41792 577010
rect 41728 576950 41780 577006
rect 41780 576950 41792 577006
rect 41728 576946 41792 576950
rect 42304 576354 42368 576418
rect 674752 576058 674816 576122
rect 41344 575910 41408 575974
rect 41920 575910 41984 575974
rect 41536 575022 41600 575086
rect 42112 574638 42176 574642
rect 42112 574582 42164 574638
rect 42164 574582 42176 574638
rect 42112 574578 42176 574582
rect 40768 573986 40832 574050
rect 40960 573098 41024 573162
rect 41920 572950 41984 573014
rect 43072 572950 43136 573014
rect 674944 568718 675008 568722
rect 674944 568662 674956 568718
rect 674956 568662 675008 568718
rect 674944 568658 675008 568662
rect 675328 562442 675392 562506
rect 674176 561998 674240 562062
rect 675520 561762 675584 561766
rect 675520 561706 675532 561762
rect 675532 561706 675584 561762
rect 675520 561702 675584 561706
rect 674944 558890 675008 558954
rect 674944 558742 675008 558806
rect 676288 558742 676352 558806
rect 674560 558150 674624 558214
rect 676864 557558 676928 557622
rect 40768 556670 40832 556734
rect 41344 555990 41408 555994
rect 41344 555934 41396 555990
rect 41396 555934 41408 555990
rect 41344 555930 41408 555934
rect 674752 554450 674816 554514
rect 40960 553562 41024 553626
rect 41344 553030 41408 553034
rect 41344 552974 41396 553030
rect 41396 552974 41408 553030
rect 41344 552970 41408 552974
rect 676480 550158 676544 550222
rect 676672 549862 676736 549926
rect 40576 544830 40640 544894
rect 41344 544830 41408 544894
rect 41152 544090 41216 544154
rect 41344 541278 41408 541342
rect 42304 541278 42368 541342
rect 42880 541130 42944 541194
rect 41920 541042 41984 541046
rect 41920 540986 41932 541042
rect 41932 540986 41984 541042
rect 41920 540982 41984 540986
rect 42112 541042 42176 541046
rect 42112 540986 42164 541042
rect 42164 540986 42176 541042
rect 42112 540982 42176 540986
rect 41152 538910 41216 538974
rect 42112 537046 42176 537050
rect 42112 536990 42124 537046
rect 42124 536990 42176 537046
rect 42112 536986 42176 536990
rect 675712 536986 675776 537050
rect 676288 536246 676352 536310
rect 40576 535654 40640 535718
rect 41536 535654 41600 535718
rect 673984 535358 674048 535422
rect 42880 535210 42944 535274
rect 675136 534618 675200 534682
rect 42304 534470 42368 534534
rect 41920 533790 41984 533794
rect 41920 533734 41972 533790
rect 41972 533734 41984 533790
rect 41920 533730 41984 533734
rect 675904 533730 675968 533794
rect 42112 532754 42176 532758
rect 42112 532698 42164 532754
rect 42164 532698 42176 532754
rect 42112 532694 42176 532698
rect 43072 532694 43136 532758
rect 676672 532694 676736 532758
rect 41536 531806 41600 531870
rect 674368 531658 674432 531722
rect 41344 531362 41408 531426
rect 40960 530030 41024 530094
rect 40768 526478 40832 526542
rect 41536 524170 41600 524174
rect 41536 524114 41588 524170
rect 41588 524114 41600 524170
rect 41536 524110 41600 524114
rect 42112 510110 42176 510114
rect 42112 510054 42164 510110
rect 42164 510054 42176 510110
rect 42112 510050 42176 510054
rect 41728 503982 41792 504046
rect 42112 504042 42176 504046
rect 42112 503986 42164 504042
rect 42164 503986 42176 504042
rect 42112 503982 42176 503986
rect 675520 492734 675584 492798
rect 675328 491402 675392 491466
rect 41728 491018 41792 491022
rect 41728 490962 41780 491018
rect 41780 490962 41792 491018
rect 41728 490958 41792 490962
rect 42112 489626 42176 489690
rect 42304 489330 42368 489394
rect 674176 487702 674240 487766
rect 674944 487406 675008 487470
rect 674560 486666 674624 486730
rect 676864 484002 676928 484066
rect 42304 483706 42368 483770
rect 42688 483706 42752 483770
rect 674752 483558 674816 483622
rect 41920 481042 41984 481106
rect 41920 463874 41984 463938
rect 41728 463726 41792 463790
rect 40384 432646 40448 432710
rect 40576 431906 40640 431970
rect 40768 430722 40832 430786
rect 40960 429390 41024 429454
rect 41344 428354 41408 428418
rect 42112 427614 42176 427678
rect 41152 426282 41216 426346
rect 41536 425098 41600 425162
rect 42112 423174 42176 423238
rect 42112 423026 42176 423090
rect 676480 412134 676544 412138
rect 676480 412078 676532 412134
rect 676532 412078 676544 412134
rect 676480 412074 676544 412078
rect 676672 411986 676736 411990
rect 676672 411930 676684 411986
rect 676684 411930 676736 411986
rect 676672 411926 676736 411930
rect 42304 409114 42368 409178
rect 42496 408818 42560 408882
rect 42112 406362 42176 406366
rect 42112 406306 42124 406362
rect 42124 406306 42176 406362
rect 42112 406302 42176 406306
rect 676480 406154 676544 406218
rect 674176 405858 674240 405922
rect 675328 405266 675392 405330
rect 676672 405266 676736 405330
rect 42496 405118 42560 405182
rect 41728 403698 41792 403702
rect 41728 403642 41780 403698
rect 41780 403642 41792 403698
rect 41728 403638 41792 403642
rect 41920 403194 41984 403258
rect 674944 403194 675008 403258
rect 41536 402602 41600 402666
rect 41344 401862 41408 401926
rect 674560 400530 674624 400594
rect 674368 400382 674432 400446
rect 40768 400086 40832 400150
rect 41152 399494 41216 399558
rect 40960 398754 41024 398818
rect 40384 390170 40448 390234
rect 40576 389134 40640 389198
rect 40768 387506 40832 387570
rect 40960 386026 41024 386090
rect 41344 385138 41408 385202
rect 42112 384398 42176 384462
rect 41152 383066 41216 383130
rect 41536 381882 41600 381946
rect 674560 378774 674624 378838
rect 675520 374482 675584 374546
rect 675712 374038 675776 374102
rect 674944 373890 675008 373954
rect 674368 371966 674432 372030
rect 42304 370486 42368 370550
rect 42112 362850 42176 362854
rect 42112 362794 42124 362850
rect 42124 362794 42176 362850
rect 42112 362790 42176 362794
rect 41920 361962 41984 361966
rect 41920 361906 41932 361962
rect 41932 361906 41984 361962
rect 41920 361902 41984 361906
rect 674368 361384 674432 361448
rect 674176 360718 674240 360782
rect 41728 360630 41792 360634
rect 41728 360574 41780 360630
rect 41780 360574 41792 360630
rect 41728 360570 41792 360574
rect 42304 360186 42368 360190
rect 42304 360130 42316 360186
rect 42316 360130 42368 360186
rect 42304 360126 42368 360130
rect 675328 360126 675392 360190
rect 673984 359978 674048 360042
rect 41536 359386 41600 359450
rect 41344 358646 41408 358710
rect 40768 356870 40832 356934
rect 41152 356426 41216 356490
rect 40960 355538 41024 355602
rect 40384 346806 40448 346870
rect 40576 346214 40640 346278
rect 676480 345474 676544 345538
rect 676288 345326 676352 345390
rect 676672 345178 676736 345242
rect 40960 344290 41024 344354
rect 40768 342810 40832 342874
rect 41152 341922 41216 341986
rect 42112 341182 42176 341246
rect 41344 338666 41408 338730
rect 41536 336446 41600 336510
rect 675520 335174 675584 335178
rect 675520 335118 675532 335174
rect 675532 335118 675584 335174
rect 675520 335114 675584 335118
rect 675328 333782 675392 333846
rect 676288 333486 676352 333550
rect 675520 329490 675584 329554
rect 676480 328010 676544 328074
rect 676672 326826 676736 326890
rect 42112 319782 42176 319786
rect 42112 319726 42124 319782
rect 42124 319726 42176 319782
rect 42112 319722 42176 319726
rect 41920 318746 41984 318750
rect 41920 318690 41932 318746
rect 41932 318690 41984 318746
rect 41920 318686 41984 318690
rect 41728 317858 41792 317862
rect 41728 317802 41780 317858
rect 41780 317802 41792 317858
rect 41728 317798 41792 317802
rect 674368 317206 674432 317270
rect 41344 316022 41408 316086
rect 674944 315874 675008 315938
rect 674176 315726 674240 315790
rect 41152 315430 41216 315494
rect 673984 314838 674048 314902
rect 674560 314246 674624 314310
rect 40960 313654 41024 313718
rect 41536 313210 41600 313274
rect 674368 313210 674432 313274
rect 40768 312322 40832 312386
rect 40384 303738 40448 303802
rect 42304 303146 42368 303210
rect 40576 302998 40640 303062
rect 42112 302258 42176 302322
rect 40768 301074 40832 301138
rect 40960 299594 41024 299658
rect 675904 299446 675968 299510
rect 676672 299298 676736 299362
rect 41152 298706 41216 298770
rect 40384 297966 40448 298030
rect 41536 295450 41600 295514
rect 41344 292342 41408 292406
rect 675520 289738 675584 289742
rect 675520 289682 675532 289738
rect 675532 289682 675584 289738
rect 675520 289678 675584 289682
rect 675328 289590 675392 289594
rect 675328 289534 675380 289590
rect 675380 289534 675392 289590
rect 675328 289530 675392 289534
rect 674752 284942 674816 285006
rect 675904 284794 675968 284858
rect 40576 284114 40640 284118
rect 40576 284058 40588 284114
rect 40588 284058 40640 284114
rect 40576 284054 40640 284058
rect 674368 283610 674432 283674
rect 42304 283374 42368 283378
rect 42304 283318 42316 283374
rect 42316 283318 42368 283374
rect 42304 283314 42368 283318
rect 42688 282426 42752 282490
rect 676672 281834 676736 281898
rect 40576 279762 40640 279826
rect 40384 276506 40448 276570
rect 41920 275530 41984 275534
rect 41920 275474 41972 275530
rect 41972 275474 41984 275530
rect 41920 275470 41984 275474
rect 42880 275470 42944 275534
rect 41728 274938 41792 274942
rect 41728 274882 41780 274938
rect 41780 274882 41792 274938
rect 41728 274878 41792 274882
rect 378496 274878 378560 274942
rect 42688 274138 42752 274202
rect 42304 273754 42368 273758
rect 42304 273698 42316 273754
rect 42316 273698 42368 273754
rect 42304 273694 42368 273698
rect 368512 273546 368576 273610
rect 378112 273606 378176 273610
rect 378112 273550 378164 273606
rect 378164 273550 378176 273606
rect 378112 273546 378176 273550
rect 378112 273250 378176 273314
rect 41536 272954 41600 273018
rect 384640 273102 384704 273166
rect 379648 272954 379712 273018
rect 197440 272658 197504 272722
rect 674944 272806 675008 272870
rect 405376 272362 405440 272426
rect 41152 272214 41216 272278
rect 379456 272214 379520 272278
rect 404224 271770 404288 271834
rect 324160 271622 324224 271686
rect 379072 271622 379136 271686
rect 403840 271622 403904 271686
rect 356992 271474 357056 271538
rect 197056 271030 197120 271094
rect 331072 271178 331136 271242
rect 387136 270882 387200 270946
rect 673984 270882 674048 270946
rect 384064 270734 384128 270798
rect 404032 270734 404096 270798
rect 40768 270586 40832 270650
rect 41728 270438 41792 270502
rect 41344 269994 41408 270058
rect 138112 269846 138176 269910
rect 674176 270142 674240 270206
rect 323008 269698 323072 269762
rect 342592 269698 342656 269762
rect 399040 269698 399104 269762
rect 138112 269550 138176 269614
rect 674560 269698 674624 269762
rect 675136 269698 675200 269762
rect 106432 269402 106496 269466
rect 106624 269402 106688 269466
rect 40960 269106 41024 269170
rect 371008 268514 371072 268578
rect 398656 268514 398720 268578
rect 389248 268366 389312 268430
rect 401152 268426 401216 268430
rect 401152 268370 401164 268426
rect 401164 268370 401216 268426
rect 401152 268366 401216 268370
rect 389248 268070 389312 268134
rect 328576 267774 328640 267838
rect 372928 267922 372992 267986
rect 377152 267982 377216 267986
rect 377152 267926 377164 267982
rect 377164 267926 377216 267982
rect 377152 267922 377216 267926
rect 396736 267922 396800 267986
rect 400384 267922 400448 267986
rect 674944 267922 675008 267986
rect 389248 267774 389312 267838
rect 267520 267626 267584 267690
rect 378688 267538 378752 267542
rect 378688 267482 378740 267538
rect 378740 267482 378752 267538
rect 378688 267478 378752 267482
rect 379072 267478 379136 267542
rect 389056 267478 389120 267542
rect 267712 267330 267776 267394
rect 396736 267390 396800 267394
rect 396736 267334 396788 267390
rect 396788 267334 396800 267390
rect 396736 267330 396800 267334
rect 374464 267242 374528 267246
rect 374464 267186 374476 267242
rect 374476 267186 374528 267242
rect 374464 267182 374528 267186
rect 328384 267094 328448 267098
rect 328384 267038 328396 267094
rect 328396 267038 328448 267094
rect 328384 267034 328448 267038
rect 328576 267034 328640 267098
rect 368512 267034 368576 267098
rect 388096 267034 388160 267098
rect 388288 267034 388352 267098
rect 389440 266886 389504 266950
rect 328384 266738 328448 266802
rect 328768 266738 328832 266802
rect 389056 266738 389120 266802
rect 389632 266738 389696 266802
rect 368512 266590 368576 266654
rect 389440 266590 389504 266654
rect 400000 266590 400064 266654
rect 400192 266650 400256 266654
rect 400192 266594 400204 266650
rect 400204 266594 400256 266650
rect 400192 266590 400256 266594
rect 400576 266590 400640 266654
rect 401344 266590 401408 266654
rect 401536 266590 401600 266654
rect 403264 266650 403328 266654
rect 403264 266594 403276 266650
rect 403276 266594 403328 266650
rect 403264 266590 403328 266594
rect 404608 266590 404672 266654
rect 404800 266650 404864 266654
rect 404800 266594 404812 266650
rect 404812 266594 404864 266650
rect 404800 266590 404864 266594
rect 405184 266650 405248 266654
rect 405184 266594 405236 266650
rect 405236 266594 405248 266650
rect 405184 266590 405248 266594
rect 406144 266650 406208 266654
rect 406144 266594 406196 266650
rect 406196 266594 406208 266650
rect 406144 266590 406208 266594
rect 406528 266650 406592 266654
rect 406528 266594 406580 266650
rect 406580 266594 406592 266650
rect 406528 266590 406592 266594
rect 406912 266650 406976 266654
rect 406912 266594 406924 266650
rect 406924 266594 406976 266650
rect 406912 266590 406976 266594
rect 407104 266650 407168 266654
rect 407104 266594 407156 266650
rect 407156 266594 407168 266650
rect 407104 266590 407168 266594
rect 409024 266650 409088 266654
rect 409024 266594 409076 266650
rect 409076 266594 409088 266650
rect 409024 266590 409088 266594
rect 409408 266650 409472 266654
rect 409408 266594 409460 266650
rect 409460 266594 409472 266650
rect 409408 266590 409472 266594
rect 674560 265406 674624 265470
rect 325504 264985 325568 264989
rect 325504 264929 325516 264985
rect 325516 264929 325568 264985
rect 325504 264925 325568 264929
rect 365056 264985 365120 264989
rect 365056 264929 365068 264985
rect 365068 264929 365120 264985
rect 365056 264925 365120 264929
rect 400768 264925 400832 264989
rect 42496 260374 42560 260438
rect 42112 259486 42176 259550
rect 41536 257858 41600 257922
rect 40384 256230 40448 256294
rect 40960 255638 41024 255702
rect 41152 254750 41216 254814
rect 40768 253418 40832 253482
rect 675712 253418 675776 253482
rect 41344 252678 41408 252742
rect 404800 247498 404864 247562
rect 42112 247114 42176 247118
rect 42112 247058 42164 247114
rect 42164 247058 42176 247114
rect 42112 247054 42176 247058
rect 42880 246758 42944 246822
rect 247552 246758 247616 246822
rect 360064 246758 360128 246822
rect 360448 246758 360512 246822
rect 367744 246758 367808 246822
rect 406336 247350 406400 247414
rect 407104 247202 407168 247266
rect 368512 246758 368576 246822
rect 369280 246758 369344 246822
rect 401344 247054 401408 247118
rect 401536 247054 401600 247118
rect 406144 247054 406208 247118
rect 404416 246906 404480 246970
rect 674752 246758 674816 246822
rect 674752 245930 674816 245934
rect 674752 245874 674804 245930
rect 674804 245874 674816 245930
rect 674752 245870 674816 245874
rect 210304 245130 210368 245194
rect 675520 245190 675584 245194
rect 675520 245134 675532 245190
rect 675532 245134 675584 245190
rect 675520 245130 675584 245134
rect 388864 244982 388928 245046
rect 401344 244982 401408 245046
rect 401920 244982 401984 245046
rect 404224 244982 404288 245046
rect 404992 244982 405056 245046
rect 406912 244982 406976 245046
rect 409024 244982 409088 245046
rect 409408 244982 409472 245046
rect 42112 244834 42176 244898
rect 247360 244686 247424 244750
rect 400768 244686 400832 244750
rect 401152 244686 401216 244750
rect 404032 244686 404096 244750
rect 404608 244686 404672 244750
rect 674176 244686 674240 244750
rect 328384 244538 328448 244602
rect 369280 244538 369344 244602
rect 400000 244538 400064 244602
rect 403840 244598 403904 244602
rect 403840 244542 403852 244598
rect 403852 244542 403904 244598
rect 403840 244538 403904 244542
rect 675136 244538 675200 244602
rect 368704 244390 368768 244454
rect 400192 244390 400256 244454
rect 367744 244242 367808 244306
rect 400576 244242 400640 244306
rect 400384 244094 400448 244158
rect 388864 243946 388928 244010
rect 403264 243946 403328 244010
rect 328576 243502 328640 243566
rect 674560 243502 674624 243566
rect 41920 242614 41984 242678
rect 42880 242614 42944 242678
rect 41728 242022 41792 242086
rect 40384 241874 40448 241938
rect 42304 241874 42368 241938
rect 675328 241874 675392 241938
rect 383104 241786 383168 241790
rect 383104 241730 383116 241786
rect 383116 241730 383168 241786
rect 383104 241726 383168 241730
rect 145408 239802 145472 239866
rect 383104 239122 383168 239126
rect 383104 239066 383116 239122
rect 383116 239066 383168 239122
rect 383104 239062 383168 239066
rect 675520 238914 675584 238978
rect 674944 238618 675008 238682
rect 212992 237582 213056 237646
rect 675712 236902 675776 236906
rect 675712 236846 675764 236902
rect 675764 236846 675776 236902
rect 675712 236842 675776 236846
rect 212992 236546 213056 236610
rect 210304 236250 210368 236314
rect 211456 234622 211520 234686
rect 212032 233734 212096 233798
rect 637312 233734 637376 233798
rect 211072 233646 211136 233650
rect 211072 233590 211084 233646
rect 211084 233590 211136 233646
rect 211072 233586 211136 233590
rect 211648 233646 211712 233650
rect 211648 233590 211700 233646
rect 211700 233590 211712 233646
rect 211648 233586 211712 233590
rect 212224 233646 212288 233650
rect 212224 233590 212236 233646
rect 212236 233590 212288 233646
rect 212224 233586 212288 233590
rect 212416 233586 212480 233650
rect 212992 233586 213056 233650
rect 636928 233586 636992 233650
rect 637504 233586 637568 233650
rect 212992 233438 213056 233502
rect 637120 233438 637184 233502
rect 637888 233498 637952 233502
rect 637888 233442 637940 233498
rect 637940 233442 637952 233498
rect 637888 233438 637952 233442
rect 41152 233290 41216 233354
rect 210880 233290 210944 233354
rect 637696 233290 637760 233354
rect 210304 232846 210368 232910
rect 212416 232846 212480 232910
rect 41920 231722 41984 231726
rect 41920 231666 41972 231722
rect 41972 231666 41984 231722
rect 41920 231662 41984 231666
rect 42112 230922 42176 230986
rect 41728 230390 41792 230394
rect 41728 230334 41780 230390
rect 41780 230334 41792 230390
rect 41728 230330 41792 230334
rect 41728 230182 41792 230246
rect 41344 229738 41408 229802
rect 40960 228998 41024 229062
rect 673984 227370 674048 227434
rect 41536 227222 41600 227286
rect 40768 226630 40832 226694
rect 42304 226186 42368 226250
rect 673984 226186 674048 226250
rect 210496 223078 210560 223142
rect 211072 223078 211136 223142
rect 674368 223078 674432 223142
rect 145600 221746 145664 221810
rect 40384 214642 40448 214706
rect 40576 213162 40640 213226
rect 40960 212422 41024 212486
rect 41152 211534 41216 211598
rect 40768 210350 40832 210414
rect 207232 210262 207296 210266
rect 207232 210206 207244 210262
rect 207244 210206 207296 210262
rect 207232 210202 207296 210206
rect 676480 210202 676544 210266
rect 676672 210054 676736 210118
rect 675904 207686 675968 207750
rect 676288 207538 676352 207602
rect 676096 207390 676160 207454
rect 210304 200582 210368 200646
rect 211072 200582 211136 200646
rect 675328 199310 675392 199314
rect 675328 199254 675380 199310
rect 675380 199254 675392 199310
rect 675328 199250 675392 199254
rect 210496 198954 210560 199018
rect 211072 198806 211136 198870
rect 41344 198658 41408 198722
rect 675520 198718 675584 198722
rect 675520 198662 675532 198718
rect 675532 198662 675584 198718
rect 675520 198658 675584 198662
rect 675904 198362 675968 198426
rect 42304 197474 42368 197538
rect 42304 195166 42368 195170
rect 42304 195110 42356 195166
rect 42356 195110 42368 195166
rect 42304 195106 42368 195110
rect 676096 195254 676160 195318
rect 674368 193478 674432 193542
rect 676288 191554 676352 191618
rect 41344 190962 41408 191026
rect 41152 190074 41216 190138
rect 207232 190134 207296 190138
rect 207232 190078 207284 190134
rect 207284 190078 207296 190134
rect 207232 190074 207296 190078
rect 41920 189098 41984 189102
rect 41920 189042 41972 189098
rect 41972 189042 41984 189098
rect 41920 189038 41984 189042
rect 41728 188358 41792 188362
rect 41728 188302 41780 188358
rect 41780 188302 41792 188358
rect 41728 188298 41792 188302
rect 40960 185930 41024 185994
rect 40384 184154 40448 184218
rect 40768 183562 40832 183626
rect 40576 182822 40640 182886
rect 673984 182526 674048 182590
rect 673984 181194 674048 181258
rect 676480 180898 676544 180962
rect 676672 179418 676736 179482
rect 674752 178530 674816 178594
rect 674176 178086 674240 178150
rect 211072 172758 211136 172822
rect 210880 172610 210944 172674
rect 210304 172462 210368 172526
rect 674560 166394 674624 166458
rect 674368 165506 674432 165570
rect 676672 164026 676736 164090
rect 676480 162842 676544 162906
rect 675904 161362 675968 161426
rect 674752 159290 674816 159354
rect 675904 157662 675968 157726
rect 675328 154614 675392 154618
rect 675328 154558 675380 154614
rect 675380 154558 675392 154614
rect 675328 154554 675392 154558
rect 675520 154258 675584 154322
rect 676480 153370 676544 153434
rect 210688 152778 210752 152842
rect 210688 152630 210752 152694
rect 211072 152630 211136 152694
rect 210304 151594 210368 151658
rect 211072 151594 211136 151658
rect 674176 148486 674240 148550
rect 674752 148338 674816 148402
rect 676672 146562 676736 146626
rect 673984 136794 674048 136858
rect 674560 135462 674624 135526
rect 674560 134870 674624 134934
rect 674368 134500 674432 134564
rect 146752 134486 146816 134490
rect 146752 134430 146804 134486
rect 146804 134430 146816 134486
rect 146752 134426 146816 134430
rect 674176 133686 674240 133750
rect 210496 132650 210560 132714
rect 211072 132650 211136 132714
rect 146752 132562 146816 132566
rect 146752 132506 146804 132562
rect 146804 132506 146816 132562
rect 146752 132502 146816 132506
rect 674944 132502 675008 132566
rect 146560 126790 146624 126794
rect 146560 126734 146572 126790
rect 146572 126734 146624 126790
rect 146560 126730 146624 126734
rect 210496 123918 210560 123982
rect 211072 123918 211136 123982
rect 209728 123770 209792 123834
rect 210880 123770 210944 123834
rect 210304 122438 210368 122502
rect 210880 122438 210944 122502
rect 675904 120366 675968 120430
rect 211072 119034 211136 119098
rect 209920 118442 209984 118506
rect 211072 118442 211136 118506
rect 676672 117998 676736 118062
rect 146560 115246 146624 115250
rect 146560 115190 146572 115246
rect 146572 115190 146624 115246
rect 146560 115186 146624 115190
rect 674176 114150 674240 114214
rect 675328 110066 675392 110070
rect 675328 110010 675380 110066
rect 675380 110010 675392 110066
rect 675328 110006 675392 110010
rect 674752 109266 674816 109330
rect 675904 108082 675968 108146
rect 210112 106750 210176 106814
rect 210880 106750 210944 106814
rect 144448 106454 144512 106518
rect 144448 103642 144512 103706
rect 674944 103198 675008 103262
rect 676672 101422 676736 101486
rect 210688 96834 210752 96898
rect 211072 96834 211136 96898
rect 210304 95798 210368 95862
rect 211072 95798 211136 95862
rect 211072 94170 211136 94234
rect 210112 93134 210176 93198
rect 211072 93134 211136 93198
rect 210304 92986 210368 93050
rect 211072 92986 211136 93050
rect 209920 82182 209984 82246
rect 210880 82182 210944 82246
rect 210496 81146 210560 81210
rect 211072 81146 211136 81210
rect 209728 77742 209792 77806
rect 210880 77742 210944 77806
rect 144832 66258 144896 66262
rect 144832 66202 144844 66258
rect 144844 66202 144896 66258
rect 144832 66198 144896 66202
rect 144832 64570 144896 64634
rect 211072 58206 211136 58270
rect 210880 54210 210944 54274
rect 212608 54210 212672 54274
rect 211264 54062 211328 54126
rect 212224 53914 212288 53978
rect 210688 53766 210752 53830
rect 211840 53618 211904 53682
rect 212992 53530 213056 53534
rect 212992 53474 213044 53530
rect 213044 53474 213056 53530
rect 212992 53470 213056 53474
rect 212416 53322 212480 53386
rect 211072 53026 211136 53090
rect 637888 52138 637952 52202
rect 637504 51990 637568 52054
rect 637696 51842 637760 51906
rect 637312 51694 637376 51758
rect 637120 51546 637184 51610
rect 145408 51398 145472 51462
rect 145600 51250 145664 51314
rect 636928 50362 636992 50426
rect 471040 46070 471104 46134
rect 302464 45034 302528 45098
rect 414784 44886 414848 44950
rect 302464 43318 302528 43322
rect 302464 43262 302516 43318
rect 302516 43262 302528 43318
rect 302464 43258 302528 43262
rect 414784 43258 414848 43322
rect 471040 42134 471104 42138
rect 471040 42078 471092 42134
rect 471092 42078 471104 42134
rect 471040 42074 471104 42078
rect 189952 41778 190016 41842
rect 194944 41778 195008 41842
rect 360064 41778 360128 41842
rect 362944 41778 363008 41842
rect 459328 41778 459392 41842
rect 360064 40890 360128 40954
rect 189952 40742 190016 40806
rect 362944 40742 363008 40806
rect 194944 40594 195008 40658
rect 455104 40298 455168 40362
<< metal4 >>
rect 83391 993630 83457 993631
rect 83391 993566 83392 993630
rect 83456 993566 83457 993630
rect 83391 993565 83457 993566
rect 83394 992151 83454 993565
rect 83391 992150 83457 992151
rect 83391 992086 83392 992150
rect 83456 992086 83457 992150
rect 83391 992085 83457 992086
rect 40959 968766 41025 968767
rect 40959 968702 40960 968766
rect 41024 968702 41025 968766
rect 40959 968701 41025 968702
rect 40575 967138 40641 967139
rect 40575 967074 40576 967138
rect 40640 967074 40641 967138
rect 40575 967073 40641 967074
rect 40383 964030 40449 964031
rect 40383 963966 40384 964030
rect 40448 963966 40449 964030
rect 40383 963965 40449 963966
rect 40386 934135 40446 963965
rect 40578 943755 40638 967073
rect 40767 965066 40833 965067
rect 40767 965002 40768 965066
rect 40832 965002 40833 965066
rect 40767 965001 40833 965002
rect 40575 943754 40641 943755
rect 40575 943690 40576 943754
rect 40640 943690 40641 943754
rect 40575 943689 40641 943690
rect 40770 937391 40830 965001
rect 40962 940647 41022 968701
rect 675327 967434 675393 967435
rect 675327 967370 675328 967434
rect 675392 967370 675393 967434
rect 675327 967369 675393 967370
rect 675135 964918 675201 964919
rect 675135 964854 675136 964918
rect 675200 964854 675201 964918
rect 675135 964853 675201 964854
rect 41535 963290 41601 963291
rect 41535 963226 41536 963290
rect 41600 963226 41601 963290
rect 41535 963225 41601 963226
rect 41151 956630 41217 956631
rect 41151 956566 41152 956630
rect 41216 956566 41217 956630
rect 41151 956565 41217 956566
rect 41154 944495 41214 956565
rect 41151 944494 41217 944495
rect 41151 944430 41152 944494
rect 41216 944430 41217 944494
rect 41151 944429 41217 944430
rect 40959 940646 41025 940647
rect 40959 940582 40960 940646
rect 41024 940582 41025 940646
rect 40959 940581 41025 940582
rect 40767 937390 40833 937391
rect 40767 937326 40768 937390
rect 40832 937326 40833 937390
rect 40767 937325 40833 937326
rect 41538 936503 41598 963225
rect 42303 962846 42369 962847
rect 42303 962782 42304 962846
rect 42368 962782 42369 962846
rect 42303 962781 42369 962782
rect 42111 962254 42177 962255
rect 42111 962190 42112 962254
rect 42176 962190 42177 962254
rect 42111 962189 42177 962190
rect 41727 959146 41793 959147
rect 41727 959082 41728 959146
rect 41792 959082 41793 959146
rect 41727 959081 41793 959082
rect 41730 938131 41790 959081
rect 41919 958406 41985 958407
rect 41919 958342 41920 958406
rect 41984 958342 41985 958406
rect 41919 958341 41985 958342
rect 41922 938871 41982 958341
rect 42114 941239 42174 962189
rect 42111 941238 42177 941239
rect 42111 941174 42112 941238
rect 42176 941174 42177 941238
rect 42111 941173 42177 941174
rect 41919 938870 41985 938871
rect 41919 938806 41920 938870
rect 41984 938806 41985 938870
rect 41919 938805 41985 938806
rect 41727 938130 41793 938131
rect 41727 938066 41728 938130
rect 41792 938066 41793 938130
rect 41727 938065 41793 938066
rect 41535 936502 41601 936503
rect 41535 936438 41536 936502
rect 41600 936438 41601 936502
rect 41535 936437 41601 936438
rect 42306 935023 42366 962781
rect 674367 962550 674433 962551
rect 674367 962486 674368 962550
rect 674432 962486 674433 962550
rect 674367 962485 674433 962486
rect 43071 962254 43137 962255
rect 43071 962190 43072 962254
rect 43136 962190 43137 962254
rect 43071 962189 43137 962190
rect 42879 962106 42945 962107
rect 42879 962042 42880 962106
rect 42944 962042 42945 962106
rect 42879 962041 42945 962042
rect 42687 959590 42753 959591
rect 42687 959526 42688 959590
rect 42752 959526 42753 959590
rect 42687 959525 42753 959526
rect 42495 957814 42561 957815
rect 42495 957750 42496 957814
rect 42560 957750 42561 957814
rect 42495 957749 42561 957750
rect 42498 941683 42558 957749
rect 42495 941682 42561 941683
rect 42495 941618 42496 941682
rect 42560 941618 42561 941682
rect 42495 941617 42561 941618
rect 42690 935319 42750 959525
rect 42687 935318 42753 935319
rect 42687 935254 42688 935318
rect 42752 935254 42753 935318
rect 42687 935253 42753 935254
rect 42303 935022 42369 935023
rect 42303 934958 42304 935022
rect 42368 934958 42369 935022
rect 42303 934957 42369 934958
rect 40383 934134 40449 934135
rect 40383 934070 40384 934134
rect 40448 934070 40449 934134
rect 40383 934069 40449 934070
rect 41343 818694 41409 818695
rect 41343 818630 41344 818694
rect 41408 818630 41409 818694
rect 41343 818629 41409 818630
rect 41151 802118 41217 802119
rect 41151 802054 41152 802118
rect 41216 802054 41217 802118
rect 41151 802053 41217 802054
rect 41154 776811 41214 802053
rect 41151 776810 41217 776811
rect 41151 776746 41152 776810
rect 41216 776746 41217 776810
rect 41151 776745 41217 776746
rect 41346 775183 41406 818629
rect 41535 802266 41601 802267
rect 41535 802202 41536 802266
rect 41600 802202 41601 802266
rect 41535 802201 41601 802202
rect 42687 802266 42753 802267
rect 42687 802202 42688 802266
rect 42752 802202 42753 802266
rect 42687 802201 42753 802202
rect 41538 791907 41598 802201
rect 41727 801970 41793 801971
rect 41727 801906 41728 801970
rect 41792 801906 41793 801970
rect 41727 801905 41793 801906
rect 41535 791906 41601 791907
rect 41535 791842 41536 791906
rect 41600 791842 41601 791906
rect 41535 791841 41601 791842
rect 41535 791018 41601 791019
rect 41535 790954 41536 791018
rect 41600 790954 41601 791018
rect 41535 790953 41601 790954
rect 41538 790239 41598 790953
rect 41730 790575 41790 801905
rect 42303 800490 42369 800491
rect 42303 800426 42304 800490
rect 42368 800426 42369 800490
rect 42303 800425 42369 800426
rect 41919 800342 41985 800343
rect 41919 800278 41920 800342
rect 41984 800278 41985 800342
rect 41919 800277 41985 800278
rect 42111 800342 42177 800343
rect 42111 800278 42112 800342
rect 42176 800278 42177 800342
rect 42111 800277 42177 800278
rect 41922 794275 41982 800277
rect 41919 794274 41985 794275
rect 41919 794210 41920 794274
rect 41984 794210 41985 794274
rect 41919 794209 41985 794210
rect 42114 793831 42174 800277
rect 42111 793830 42177 793831
rect 42111 793766 42112 793830
rect 42176 793766 42177 793830
rect 42111 793765 42177 793766
rect 42306 793569 42366 800425
rect 42495 799750 42561 799751
rect 42495 799686 42496 799750
rect 42560 799686 42561 799750
rect 42495 799685 42561 799686
rect 42114 793509 42366 793569
rect 42114 791759 42174 793509
rect 42498 792499 42558 799685
rect 42690 798419 42750 802201
rect 42687 798418 42753 798419
rect 42687 798354 42688 798418
rect 42752 798354 42753 798418
rect 42687 798353 42753 798354
rect 42495 792498 42561 792499
rect 42495 792434 42496 792498
rect 42560 792434 42561 792498
rect 42495 792433 42561 792434
rect 42303 792350 42369 792351
rect 42303 792286 42304 792350
rect 42368 792286 42369 792350
rect 42303 792285 42369 792286
rect 42111 791758 42177 791759
rect 42111 791694 42112 791758
rect 42176 791694 42177 791758
rect 42111 791693 42177 791694
rect 42111 791166 42177 791167
rect 42111 791102 42112 791166
rect 42176 791102 42177 791166
rect 42111 791101 42177 791102
rect 41727 790574 41793 790575
rect 41727 790510 41728 790574
rect 41792 790510 41793 790574
rect 41727 790509 41793 790510
rect 41538 790179 41790 790239
rect 41535 775922 41601 775923
rect 41535 775858 41536 775922
rect 41600 775858 41601 775922
rect 41535 775857 41601 775858
rect 41343 775182 41409 775183
rect 41343 775118 41344 775182
rect 41408 775118 41409 775182
rect 41343 775117 41409 775118
rect 41151 760234 41217 760235
rect 41151 760170 41152 760234
rect 41216 760170 41217 760234
rect 41151 760169 41217 760170
rect 40767 758754 40833 758755
rect 40767 758690 40768 758754
rect 40832 758690 40833 758754
rect 40767 758689 40833 758690
rect 40770 747211 40830 758689
rect 40959 757274 41025 757275
rect 40959 757210 40960 757274
rect 41024 757210 41025 757274
rect 40959 757209 41025 757210
rect 40962 748691 41022 757209
rect 40959 748690 41025 748691
rect 40959 748626 40960 748690
rect 41024 748626 41025 748690
rect 40959 748625 41025 748626
rect 40767 747210 40833 747211
rect 40767 747146 40768 747210
rect 40832 747146 40833 747210
rect 40767 747145 40833 747146
rect 41154 746767 41214 760169
rect 41151 746766 41217 746767
rect 41151 746702 41152 746766
rect 41216 746702 41217 746766
rect 41151 746701 41217 746702
rect 41346 733151 41406 775117
rect 41538 733891 41598 775857
rect 41730 761601 41790 790179
rect 41730 761541 41982 761601
rect 41727 757126 41793 757127
rect 41727 757062 41728 757126
rect 41792 757062 41793 757126
rect 41727 757061 41793 757062
rect 41730 747507 41790 757061
rect 41922 752943 41982 761541
rect 42114 757275 42174 791101
rect 42306 788651 42366 792285
rect 42882 791019 42942 962041
rect 43074 791167 43134 962189
rect 674175 961514 674241 961515
rect 674175 961450 674176 961514
rect 674240 961450 674241 961514
rect 674175 961449 674241 961450
rect 674178 931619 674238 961449
rect 674370 934727 674430 962485
rect 674559 962254 674625 962255
rect 674559 962190 674560 962254
rect 674624 962190 674625 962254
rect 674559 962189 674625 962190
rect 674367 934726 674433 934727
rect 674367 934662 674368 934726
rect 674432 934662 674433 934726
rect 674367 934661 674433 934662
rect 674562 934579 674622 962189
rect 674751 957814 674817 957815
rect 674751 957750 674752 957814
rect 674816 957750 674817 957814
rect 674751 957749 674817 957750
rect 674559 934578 674625 934579
rect 674559 934514 674560 934578
rect 674624 934514 674625 934578
rect 674559 934513 674625 934514
rect 674754 932951 674814 957749
rect 674943 956038 675009 956039
rect 674943 955974 674944 956038
rect 675008 955974 675009 956038
rect 674943 955973 675009 955974
rect 674946 933395 675006 955973
rect 675138 940943 675198 964853
rect 675330 961367 675390 967369
rect 676671 966398 676737 966399
rect 676671 966334 676672 966398
rect 676736 966334 676737 966398
rect 676671 966333 676737 966334
rect 675711 965806 675777 965807
rect 675711 965742 675712 965806
rect 675776 965742 675777 965806
rect 675711 965741 675777 965742
rect 675327 961366 675393 961367
rect 675327 961302 675328 961366
rect 675392 961302 675393 961366
rect 675327 961301 675393 961302
rect 675135 940942 675201 940943
rect 675135 940878 675136 940942
rect 675200 940878 675201 940942
rect 675135 940877 675201 940878
rect 674943 933394 675009 933395
rect 674943 933330 674944 933394
rect 675008 933330 675009 933394
rect 674943 933329 675009 933330
rect 674751 932950 674817 932951
rect 674751 932886 674752 932950
rect 674816 932886 674817 932950
rect 674751 932885 674817 932886
rect 674175 931618 674241 931619
rect 674175 931554 674176 931618
rect 674240 931554 674241 931618
rect 674175 931553 674241 931554
rect 673983 876562 674049 876563
rect 673983 876498 673984 876562
rect 674048 876498 674049 876562
rect 673983 876497 674049 876498
rect 43071 791166 43137 791167
rect 43071 791102 43072 791166
rect 43136 791102 43137 791166
rect 43071 791101 43137 791102
rect 42879 791018 42945 791019
rect 42879 790954 42880 791018
rect 42944 790954 42945 791018
rect 42879 790953 42945 790954
rect 42303 788650 42369 788651
rect 42303 788586 42304 788650
rect 42368 788586 42369 788650
rect 42303 788585 42369 788586
rect 42495 764082 42561 764083
rect 42495 764018 42496 764082
rect 42560 764018 42561 764082
rect 42495 764017 42561 764018
rect 42111 757274 42177 757275
rect 42111 757210 42112 757274
rect 42176 757210 42177 757274
rect 42111 757209 42177 757210
rect 42111 757126 42177 757127
rect 42111 757062 42112 757126
rect 42176 757062 42177 757126
rect 42111 757061 42177 757062
rect 42114 753131 42174 757061
rect 42111 753130 42177 753131
rect 42111 753066 42112 753130
rect 42176 753066 42177 753130
rect 42111 753065 42177 753066
rect 41922 752883 42174 752943
rect 41919 748690 41985 748691
rect 41919 748626 41920 748690
rect 41984 748626 41985 748690
rect 41919 748625 41985 748626
rect 41727 747506 41793 747507
rect 41727 747442 41728 747506
rect 41792 747442 41793 747506
rect 41727 747441 41793 747442
rect 41727 747358 41793 747359
rect 41727 747294 41728 747358
rect 41792 747294 41793 747358
rect 41727 747293 41793 747294
rect 41535 733890 41601 733891
rect 41535 733826 41536 733890
rect 41600 733826 41601 733890
rect 41535 733825 41601 733826
rect 41343 733150 41409 733151
rect 41343 733086 41344 733150
rect 41408 733086 41409 733150
rect 41343 733085 41409 733086
rect 41151 726342 41217 726343
rect 41151 726278 41152 726342
rect 41216 726278 41217 726342
rect 41151 726277 41217 726278
rect 41154 705475 41214 726277
rect 41343 714206 41409 714207
rect 41343 714142 41344 714206
rect 41408 714142 41409 714206
rect 41343 714141 41409 714142
rect 41346 711099 41406 714141
rect 41343 711098 41409 711099
rect 41343 711034 41344 711098
rect 41408 711034 41409 711098
rect 41343 711033 41409 711034
rect 41151 705474 41217 705475
rect 41151 705410 41152 705474
rect 41216 705410 41217 705474
rect 41151 705409 41217 705410
rect 41538 690379 41598 733825
rect 41730 715647 41790 747293
rect 41922 722495 41982 748625
rect 42114 747359 42174 752883
rect 42498 751799 42558 764017
rect 42879 760530 42945 760531
rect 42879 760466 42880 760530
rect 42944 760466 42945 760530
rect 42879 760465 42945 760466
rect 42687 758458 42753 758459
rect 42687 758394 42688 758458
rect 42752 758394 42753 758458
rect 42687 758393 42753 758394
rect 42495 751798 42561 751799
rect 42495 751734 42496 751798
rect 42560 751734 42561 751798
rect 42495 751733 42561 751734
rect 42690 751059 42750 758393
rect 42687 751058 42753 751059
rect 42687 750994 42688 751058
rect 42752 750994 42753 751058
rect 42687 750993 42753 750994
rect 42111 747358 42177 747359
rect 42111 747294 42112 747358
rect 42176 747294 42177 747358
rect 42111 747293 42177 747294
rect 42882 746027 42942 760465
rect 43071 757422 43137 757423
rect 43071 757358 43072 757422
rect 43136 757358 43137 757422
rect 43071 757357 43137 757358
rect 43074 751799 43134 757357
rect 673986 757127 674046 876497
rect 674751 875970 674817 875971
rect 674751 875906 674752 875970
rect 674816 875906 674817 875970
rect 674751 875905 674817 875906
rect 674559 874046 674625 874047
rect 674559 873982 674560 874046
rect 674624 873982 674625 874046
rect 674559 873981 674625 873982
rect 674175 873454 674241 873455
rect 674175 873390 674176 873454
rect 674240 873390 674241 873454
rect 674175 873389 674241 873390
rect 673983 757126 674049 757127
rect 673983 757062 673984 757126
rect 674048 757062 674049 757126
rect 673983 757061 674049 757062
rect 674178 756387 674238 873389
rect 674367 780658 674433 780659
rect 674367 780594 674368 780658
rect 674432 780594 674433 780658
rect 674367 780593 674433 780594
rect 674175 756386 674241 756387
rect 674175 756322 674176 756386
rect 674240 756322 674241 756386
rect 674175 756321 674241 756322
rect 43071 751798 43137 751799
rect 43071 751734 43072 751798
rect 43136 751734 43137 751798
rect 43071 751733 43137 751734
rect 42879 746026 42945 746027
rect 42879 745962 42880 746026
rect 42944 745962 42945 746026
rect 42879 745961 42945 745962
rect 42111 732262 42177 732263
rect 42111 732198 42112 732262
rect 42176 732198 42177 732262
rect 42111 732197 42177 732198
rect 42114 725603 42174 732197
rect 43071 729598 43137 729599
rect 43071 729534 43072 729598
rect 43136 729534 43137 729598
rect 43071 729533 43137 729534
rect 42111 725602 42177 725603
rect 42111 725538 42112 725602
rect 42176 725538 42177 725602
rect 42111 725537 42177 725538
rect 41919 722494 41985 722495
rect 41919 722430 41920 722494
rect 41984 722430 41985 722494
rect 41919 722429 41985 722430
rect 42495 722494 42561 722495
rect 42495 722430 42496 722494
rect 42560 722430 42561 722494
rect 42495 722429 42561 722430
rect 41730 715587 42174 715647
rect 41919 714354 41985 714355
rect 41919 714290 41920 714354
rect 41984 714290 41985 714354
rect 41919 714289 41985 714290
rect 41727 713910 41793 713911
rect 41727 713846 41728 713910
rect 41792 713846 41793 713910
rect 41727 713845 41793 713846
rect 41730 706807 41790 713845
rect 41922 707991 41982 714289
rect 41919 707990 41985 707991
rect 41919 707926 41920 707990
rect 41984 707926 41985 707990
rect 41919 707925 41985 707926
rect 41727 706806 41793 706807
rect 41727 706742 41728 706806
rect 41792 706742 41793 706806
rect 41727 706741 41793 706742
rect 42114 704991 42174 715587
rect 42303 705770 42369 705771
rect 42303 705706 42304 705770
rect 42368 705706 42369 705770
rect 42303 705705 42369 705706
rect 41730 704931 42174 704991
rect 41730 704143 41790 704931
rect 42111 704734 42177 704735
rect 42111 704670 42112 704734
rect 42176 704670 42177 704734
rect 42111 704669 42177 704670
rect 41727 704142 41793 704143
rect 41727 704078 41728 704142
rect 41792 704078 41793 704142
rect 41727 704077 41793 704078
rect 41535 690378 41601 690379
rect 41535 690314 41536 690378
rect 41600 690314 41601 690378
rect 41535 690313 41601 690314
rect 41730 675687 41790 704077
rect 42114 702327 42174 704669
rect 41538 675627 41790 675687
rect 41922 702267 42174 702327
rect 40767 673950 40833 673951
rect 40767 673886 40768 673950
rect 40832 673886 40833 673950
rect 40767 673885 40833 673886
rect 40575 672618 40641 672619
rect 40575 672554 40576 672618
rect 40640 672554 40641 672618
rect 40575 672553 40641 672554
rect 40578 656635 40638 672553
rect 40770 662407 40830 673885
rect 41538 663033 41598 675627
rect 41922 675431 41982 702267
rect 42111 689638 42177 689639
rect 42111 689574 42112 689638
rect 42176 689574 42177 689638
rect 42111 689573 42177 689574
rect 41919 675430 41985 675431
rect 41919 675366 41920 675430
rect 41984 675366 41985 675430
rect 41919 675365 41985 675366
rect 41727 670990 41793 670991
rect 41727 670926 41728 670990
rect 41792 670926 41793 670990
rect 41727 670925 41793 670926
rect 41154 662973 41598 663033
rect 40767 662406 40833 662407
rect 40767 662342 40768 662406
rect 40832 662342 40833 662406
rect 40767 662341 40833 662342
rect 41154 660779 41214 662973
rect 41151 660778 41217 660779
rect 41151 660714 41152 660778
rect 41216 660714 41217 660778
rect 41151 660713 41217 660714
rect 41730 660335 41790 670925
rect 41919 670842 41985 670843
rect 41919 670778 41920 670842
rect 41984 670778 41985 670842
rect 41919 670777 41985 670778
rect 41727 660334 41793 660335
rect 41727 660270 41728 660334
rect 41792 660270 41793 660334
rect 41727 660269 41793 660270
rect 41727 660186 41793 660187
rect 41727 660122 41728 660186
rect 41792 660122 41793 660186
rect 41727 660121 41793 660122
rect 40575 656634 40641 656635
rect 40575 656570 40576 656634
rect 40640 656570 40641 656634
rect 40575 656569 40641 656570
rect 41730 628401 41790 660121
rect 41922 659151 41982 670777
rect 41919 659150 41985 659151
rect 41919 659086 41920 659150
rect 41984 659086 41985 659150
rect 41919 659085 41985 659086
rect 41919 659002 41985 659003
rect 41919 658938 41920 659002
rect 41984 658938 41985 659002
rect 41919 658937 41985 658938
rect 41922 635061 41982 658937
rect 42114 647459 42174 689573
rect 42306 688751 42366 705705
rect 42498 704735 42558 722429
rect 42879 714206 42945 714207
rect 42879 714142 42880 714206
rect 42944 714142 42945 714206
rect 42879 714141 42945 714142
rect 42687 713910 42753 713911
rect 42687 713846 42688 713910
rect 42752 713846 42753 713910
rect 42687 713845 42753 713846
rect 42690 709767 42750 713845
rect 42687 709766 42753 709767
rect 42687 709702 42688 709766
rect 42752 709702 42753 709766
rect 42687 709701 42753 709702
rect 42882 707991 42942 714141
rect 42879 707990 42945 707991
rect 42879 707926 42880 707990
rect 42944 707926 42945 707990
rect 42879 707925 42945 707926
rect 42495 704734 42561 704735
rect 42495 704670 42496 704734
rect 42560 704670 42561 704734
rect 42495 704669 42561 704670
rect 43074 702811 43134 729533
rect 43455 725602 43521 725603
rect 43455 725538 43456 725602
rect 43520 725538 43521 725602
rect 43455 725537 43521 725538
rect 43263 721458 43329 721459
rect 43263 721394 43264 721458
rect 43328 721394 43329 721458
rect 43263 721393 43329 721394
rect 43266 708583 43326 721393
rect 43263 708582 43329 708583
rect 43263 708518 43264 708582
rect 43328 708518 43329 708582
rect 43263 708517 43329 708518
rect 43458 705919 43518 725537
rect 673983 717018 674049 717019
rect 673983 716954 673984 717018
rect 674048 716954 674049 717018
rect 673983 716953 674049 716954
rect 43455 705918 43521 705919
rect 43455 705854 43456 705918
rect 43520 705854 43521 705918
rect 43455 705853 43521 705854
rect 43071 702810 43137 702811
rect 43071 702746 43072 702810
rect 43136 702746 43137 702810
rect 43071 702745 43137 702746
rect 42303 688750 42369 688751
rect 42303 688686 42304 688750
rect 42368 688686 42369 688750
rect 42303 688685 42369 688686
rect 42111 647458 42177 647459
rect 42111 647394 42112 647458
rect 42176 647394 42177 647458
rect 42111 647393 42177 647394
rect 42306 646719 42366 688685
rect 42879 675430 42945 675431
rect 42879 675366 42880 675430
rect 42944 675366 42945 675430
rect 42879 675365 42945 675366
rect 42687 670990 42753 670991
rect 42687 670926 42688 670990
rect 42752 670926 42753 670990
rect 42687 670925 42753 670926
rect 42495 670842 42561 670843
rect 42495 670778 42496 670842
rect 42560 670778 42561 670842
rect 42495 670777 42561 670778
rect 42498 662851 42558 670777
rect 42690 663443 42750 670925
rect 42687 663442 42753 663443
rect 42687 663378 42688 663442
rect 42752 663378 42753 663442
rect 42687 663377 42753 663378
rect 42495 662850 42561 662851
rect 42495 662786 42496 662850
rect 42560 662786 42561 662850
rect 42495 662785 42561 662786
rect 42882 662367 42942 675365
rect 673986 673063 674046 716953
rect 674370 713763 674430 780593
rect 674562 760087 674622 873981
rect 674754 762455 674814 875905
rect 675330 875823 675390 961301
rect 675519 960182 675585 960183
rect 675519 960118 675520 960182
rect 675584 960118 675585 960182
rect 675519 960117 675585 960118
rect 675327 875822 675393 875823
rect 675327 875758 675328 875822
rect 675392 875758 675393 875822
rect 675327 875757 675393 875758
rect 675522 875675 675582 960117
rect 675714 935911 675774 965741
rect 676479 963290 676545 963291
rect 676479 963226 676480 963290
rect 676544 963226 676545 963290
rect 676479 963225 676545 963226
rect 676095 959146 676161 959147
rect 676095 959082 676096 959146
rect 676160 959082 676161 959146
rect 676095 959081 676161 959082
rect 676098 937391 676158 959081
rect 676482 938131 676542 963225
rect 676674 939315 676734 966333
rect 677055 953522 677121 953523
rect 677055 953458 677056 953522
rect 677120 953458 677121 953522
rect 677055 953457 677121 953458
rect 676863 953374 676929 953375
rect 676863 953310 676864 953374
rect 676928 953310 676929 953374
rect 676863 953309 676929 953310
rect 676671 939314 676737 939315
rect 676671 939250 676672 939314
rect 676736 939250 676737 939314
rect 676671 939249 676737 939250
rect 676479 938130 676545 938131
rect 676479 938066 676480 938130
rect 676544 938066 676545 938130
rect 676479 938065 676545 938066
rect 676095 937390 676161 937391
rect 676095 937326 676096 937390
rect 676160 937326 676161 937390
rect 676095 937325 676161 937326
rect 675711 935910 675777 935911
rect 675711 935846 675712 935910
rect 675776 935846 675777 935910
rect 675711 935845 675777 935846
rect 676866 930287 676926 953309
rect 677058 931471 677118 953457
rect 677055 931470 677121 931471
rect 677055 931406 677056 931470
rect 677120 931406 677121 931470
rect 677055 931405 677121 931406
rect 676863 930286 676929 930287
rect 676863 930222 676864 930286
rect 676928 930222 676929 930286
rect 676863 930221 676929 930222
rect 676095 877006 676161 877007
rect 676095 876942 676096 877006
rect 676160 876942 676161 877006
rect 676095 876941 676161 876942
rect 675519 875674 675585 875675
rect 675519 875610 675520 875674
rect 675584 875610 675585 875674
rect 675519 875609 675585 875610
rect 674943 869902 675009 869903
rect 674943 869838 674944 869902
rect 675008 869838 675009 869902
rect 674943 869837 675009 869838
rect 674751 762454 674817 762455
rect 674751 762390 674752 762454
rect 674816 762390 674817 762454
rect 674751 762389 674817 762390
rect 674559 760086 674625 760087
rect 674559 760022 674560 760086
rect 674624 760022 674625 760086
rect 674559 760021 674625 760022
rect 674946 759199 675006 869837
rect 675327 862946 675393 862947
rect 675327 862882 675328 862946
rect 675392 862882 675393 862946
rect 675327 862881 675393 862882
rect 675135 773702 675201 773703
rect 675135 773638 675136 773702
rect 675200 773638 675201 773702
rect 675135 773637 675201 773638
rect 674943 759198 675009 759199
rect 674943 759134 674944 759198
rect 675008 759134 675009 759198
rect 674943 759133 675009 759134
rect 674559 743214 674625 743215
rect 674559 743150 674560 743214
rect 674624 743150 674625 743214
rect 674559 743149 674625 743150
rect 674367 713762 674433 713763
rect 674367 713698 674368 713762
rect 674432 713698 674433 713762
rect 674367 713697 674433 713698
rect 674175 694374 674241 694375
rect 674175 694310 674176 694374
rect 674240 694310 674241 694374
rect 674175 694309 674241 694310
rect 673983 673062 674049 673063
rect 673983 672998 673984 673062
rect 674048 672998 674049 673062
rect 673983 672997 674049 672998
rect 43071 670990 43137 670991
rect 43071 670926 43072 670990
rect 43136 670926 43137 670990
rect 43071 670925 43137 670926
rect 43074 665367 43134 670925
rect 43071 665366 43137 665367
rect 43071 665302 43072 665366
rect 43136 665302 43137 665366
rect 43071 665301 43137 665302
rect 42498 662307 42942 662367
rect 42498 661519 42558 662307
rect 42495 661518 42561 661519
rect 42495 661454 42496 661518
rect 42560 661454 42561 661518
rect 42495 661453 42561 661454
rect 42498 659003 42558 661453
rect 42495 659002 42561 659003
rect 42495 658938 42496 659002
rect 42560 658938 42561 659002
rect 42495 658937 42561 658938
rect 42303 646718 42369 646719
rect 42303 646654 42304 646718
rect 42368 646654 42369 646718
rect 42303 646653 42369 646654
rect 673983 640354 674049 640355
rect 673983 640290 673984 640354
rect 674048 640290 674049 640354
rect 673983 640289 674049 640290
rect 42687 638948 42753 638949
rect 42687 638884 42688 638948
rect 42752 638884 42753 638948
rect 42687 638883 42753 638884
rect 41922 635001 42366 635061
rect 41538 628341 41790 628401
rect 40767 628218 40833 628219
rect 40767 628154 40768 628218
rect 40832 628154 40833 628218
rect 40767 628153 40833 628154
rect 40575 627922 40641 627923
rect 40575 627858 40576 627922
rect 40640 627858 40641 627922
rect 40575 627857 40641 627858
rect 40578 612827 40638 627857
rect 40770 613419 40830 628153
rect 41343 627774 41409 627775
rect 41343 627710 41344 627774
rect 41408 627710 41409 627774
rect 41343 627709 41409 627710
rect 41346 616527 41406 627709
rect 41538 618303 41598 628341
rect 41727 627774 41793 627775
rect 41727 627710 41728 627774
rect 41792 627710 41793 627774
rect 41727 627709 41793 627710
rect 41535 618302 41601 618303
rect 41535 618238 41536 618302
rect 41600 618238 41601 618302
rect 41535 618237 41601 618238
rect 41538 617079 41598 618237
rect 41730 617859 41790 627709
rect 41919 627626 41985 627627
rect 41919 627562 41920 627626
rect 41984 627562 41985 627626
rect 41919 627561 41985 627562
rect 41922 620819 41982 627561
rect 42111 627478 42177 627479
rect 42111 627414 42112 627478
rect 42176 627414 42177 627478
rect 42111 627413 42177 627414
rect 42114 621707 42174 627413
rect 42306 624963 42366 635001
rect 42690 625111 42750 638883
rect 42687 625110 42753 625111
rect 42687 625046 42688 625110
rect 42752 625046 42753 625110
rect 42687 625045 42753 625046
rect 42303 624962 42369 624963
rect 42303 624898 42304 624962
rect 42368 624898 42369 624962
rect 42303 624897 42369 624898
rect 42495 624814 42561 624815
rect 42495 624750 42496 624814
rect 42560 624750 42561 624814
rect 42495 624749 42561 624750
rect 42111 621706 42177 621707
rect 42111 621642 42112 621706
rect 42176 621642 42177 621706
rect 42111 621641 42177 621642
rect 41919 620818 41985 620819
rect 41919 620754 41920 620818
rect 41984 620754 41985 620818
rect 41919 620753 41985 620754
rect 42498 618155 42558 624749
rect 41919 618154 41985 618155
rect 41919 618090 41920 618154
rect 41984 618090 41985 618154
rect 41919 618089 41985 618090
rect 42495 618154 42561 618155
rect 42495 618090 42496 618154
rect 42560 618090 42561 618154
rect 42495 618089 42561 618090
rect 41727 617858 41793 617859
rect 41727 617794 41728 617858
rect 41792 617794 41793 617858
rect 41727 617793 41793 617794
rect 41538 617019 41790 617079
rect 41343 616526 41409 616527
rect 41343 616462 41344 616526
rect 41408 616462 41409 616526
rect 41343 616461 41409 616462
rect 40767 613418 40833 613419
rect 40767 613354 40768 613418
rect 40832 613354 40833 613418
rect 40767 613353 40833 613354
rect 40575 612826 40641 612827
rect 40575 612762 40576 612826
rect 40640 612762 40641 612826
rect 40575 612761 40641 612762
rect 40959 599950 41025 599951
rect 40959 599886 40960 599950
rect 41024 599886 41025 599950
rect 40959 599885 41025 599886
rect 40767 596842 40833 596843
rect 40767 596778 40768 596842
rect 40832 596778 40833 596842
rect 40767 596777 40833 596778
rect 40770 574051 40830 596777
rect 40767 574050 40833 574051
rect 40767 573986 40768 574050
rect 40832 573986 40833 574050
rect 40767 573985 40833 573986
rect 40962 573163 41022 599885
rect 41151 594474 41217 594475
rect 41151 594410 41152 594474
rect 41216 594410 41217 594474
rect 41151 594409 41217 594410
rect 41154 580267 41214 594409
rect 41730 591105 41790 617019
rect 41922 604983 41982 618089
rect 673986 613419 674046 640289
rect 674178 621115 674238 694309
rect 674367 693486 674433 693487
rect 674367 693422 674368 693486
rect 674432 693422 674433 693486
rect 674367 693421 674433 693422
rect 674175 621114 674241 621115
rect 674175 621050 674176 621114
rect 674240 621050 674241 621114
rect 674175 621049 674241 621050
rect 674370 620375 674430 693421
rect 674562 670547 674622 743149
rect 674943 740402 675009 740403
rect 674943 740338 674944 740402
rect 675008 740338 675009 740402
rect 674943 740337 675009 740338
rect 674751 739366 674817 739367
rect 674751 739302 674752 739366
rect 674816 739302 674817 739366
rect 674751 739301 674817 739302
rect 674559 670546 674625 670547
rect 674559 670482 674560 670546
rect 674624 670482 674625 670546
rect 674559 670481 674625 670482
rect 674754 666699 674814 739301
rect 674946 669807 675006 740337
rect 675138 713615 675198 773637
rect 675330 758607 675390 862881
rect 675711 788058 675777 788059
rect 675711 787994 675712 788058
rect 675776 787994 675777 788058
rect 675711 787993 675777 787994
rect 675519 787170 675585 787171
rect 675519 787106 675520 787170
rect 675584 787106 675585 787170
rect 675519 787105 675585 787106
rect 675327 758606 675393 758607
rect 675327 758542 675328 758606
rect 675392 758542 675393 758606
rect 675327 758541 675393 758542
rect 675327 738626 675393 738627
rect 675327 738562 675328 738626
rect 675392 738562 675393 738626
rect 675327 738561 675393 738562
rect 675135 713614 675201 713615
rect 675135 713550 675136 713614
rect 675200 713550 675201 713614
rect 675135 713549 675201 713550
rect 675135 689194 675201 689195
rect 675135 689130 675136 689194
rect 675200 689130 675201 689194
rect 675135 689129 675201 689130
rect 674943 669806 675009 669807
rect 674943 669742 674944 669806
rect 675008 669742 675009 669806
rect 674943 669741 675009 669742
rect 674751 666698 674817 666699
rect 674751 666634 674752 666698
rect 674816 666634 674817 666698
rect 674751 666633 674817 666634
rect 674559 652194 674625 652195
rect 674559 652130 674560 652194
rect 674624 652130 674625 652194
rect 674559 652129 674625 652130
rect 674367 620374 674433 620375
rect 674367 620310 674368 620374
rect 674432 620310 674433 620374
rect 674367 620309 674433 620310
rect 673983 613418 674049 613419
rect 673983 613354 673984 613418
rect 674048 613354 674049 613418
rect 673983 613353 674049 613354
rect 673983 607794 674049 607795
rect 673983 607730 673984 607794
rect 674048 607730 674049 607794
rect 673983 607729 674049 607730
rect 41919 604982 41985 604983
rect 41919 604918 41920 604982
rect 41984 604918 41985 604982
rect 41919 604917 41985 604918
rect 42111 604834 42177 604835
rect 42111 604770 42112 604834
rect 42176 604770 42177 604834
rect 42111 604769 42177 604770
rect 41730 591045 41982 591105
rect 41343 586038 41409 586039
rect 41343 585974 41344 586038
rect 41408 585974 41409 586038
rect 41343 585973 41409 585974
rect 41151 580266 41217 580267
rect 41151 580202 41152 580266
rect 41216 580202 41217 580266
rect 41151 580201 41217 580202
rect 41346 575975 41406 585973
rect 41922 584852 41982 591045
rect 42114 586039 42174 604769
rect 43071 593734 43137 593735
rect 43071 593670 43072 593734
rect 43136 593670 43137 593734
rect 43071 593669 43137 593670
rect 42111 586038 42177 586039
rect 42111 585974 42112 586038
rect 42176 585974 42177 586038
rect 42111 585973 42177 585974
rect 41586 584792 41982 584852
rect 42495 584854 42561 584855
rect 41586 584704 41646 584792
rect 42495 584790 42496 584854
rect 42560 584790 42561 584854
rect 42495 584789 42561 584790
rect 41538 584644 41646 584704
rect 42303 584706 42369 584707
rect 41343 575974 41409 575975
rect 41343 575910 41344 575974
rect 41408 575910 41409 575974
rect 41343 575909 41409 575910
rect 41538 575087 41598 584644
rect 42303 584642 42304 584706
rect 42368 584642 42369 584706
rect 42303 584641 42369 584642
rect 41727 584558 41793 584559
rect 41727 584494 41728 584558
rect 41792 584494 41793 584558
rect 41727 584493 41793 584494
rect 41730 577011 41790 584493
rect 41919 584410 41985 584411
rect 41919 584346 41920 584410
rect 41984 584346 41985 584410
rect 41919 584345 41985 584346
rect 41922 582043 41982 584345
rect 42111 584262 42177 584263
rect 42111 584198 42112 584262
rect 42176 584198 42177 584262
rect 42111 584197 42177 584198
rect 41919 582042 41985 582043
rect 41919 581978 41920 582042
rect 41984 581978 41985 582042
rect 41919 581977 41985 581978
rect 41727 577010 41793 577011
rect 41727 576946 41728 577010
rect 41792 576946 41793 577010
rect 41727 576945 41793 576946
rect 41919 575974 41985 575975
rect 41919 575910 41920 575974
rect 41984 575910 41985 575974
rect 41919 575909 41985 575910
rect 41535 575086 41601 575087
rect 41535 575022 41536 575086
rect 41600 575022 41601 575086
rect 41535 575021 41601 575022
rect 40959 573162 41025 573163
rect 40959 573098 40960 573162
rect 41024 573098 41025 573162
rect 40959 573097 41025 573098
rect 41538 570459 41598 575021
rect 41922 573015 41982 575909
rect 42114 574643 42174 584197
rect 42306 576419 42366 584641
rect 42498 577603 42558 584789
rect 42879 584706 42945 584707
rect 42879 584642 42880 584706
rect 42944 584642 42945 584706
rect 42879 584641 42945 584642
rect 42687 583818 42753 583819
rect 42687 583754 42688 583818
rect 42752 583754 42753 583818
rect 42687 583753 42753 583754
rect 42690 578935 42750 583753
rect 42687 578934 42753 578935
rect 42687 578870 42688 578934
rect 42752 578870 42753 578934
rect 42687 578869 42753 578870
rect 42882 578343 42942 584641
rect 43074 581451 43134 593669
rect 43071 581450 43137 581451
rect 43071 581386 43072 581450
rect 43136 581386 43137 581450
rect 43071 581385 43137 581386
rect 42879 578342 42945 578343
rect 42879 578278 42880 578342
rect 42944 578278 42945 578342
rect 42879 578277 42945 578278
rect 42495 577602 42561 577603
rect 42495 577538 42496 577602
rect 42560 577538 42561 577602
rect 42495 577537 42561 577538
rect 42303 576418 42369 576419
rect 42303 576354 42304 576418
rect 42368 576354 42369 576418
rect 42303 576353 42369 576354
rect 42111 574642 42177 574643
rect 42111 574578 42112 574642
rect 42176 574578 42177 574642
rect 42111 574577 42177 574578
rect 41919 573014 41985 573015
rect 41919 572950 41920 573014
rect 41984 572950 41985 573014
rect 41919 572949 41985 572950
rect 43071 573014 43137 573015
rect 43071 572950 43072 573014
rect 43136 572950 43137 573014
rect 43071 572949 43137 572950
rect 41346 570399 41598 570459
rect 40767 556734 40833 556735
rect 40767 556670 40768 556734
rect 40832 556670 40833 556734
rect 40767 556669 40833 556670
rect 40575 544894 40641 544895
rect 40575 544830 40576 544894
rect 40640 544830 40641 544894
rect 40575 544829 40641 544830
rect 40578 535719 40638 544829
rect 40575 535718 40641 535719
rect 40575 535654 40576 535718
rect 40640 535654 40641 535718
rect 40575 535653 40641 535654
rect 40770 526543 40830 556669
rect 41346 555995 41406 570399
rect 41343 555994 41409 555995
rect 41343 555930 41344 555994
rect 41408 555930 41409 555994
rect 41343 555929 41409 555930
rect 40959 553626 41025 553627
rect 40959 553562 40960 553626
rect 41024 553562 41025 553626
rect 40959 553561 41025 553562
rect 40962 530095 41022 553561
rect 41343 553034 41409 553035
rect 41343 552970 41344 553034
rect 41408 552970 41409 553034
rect 41343 552969 41409 552970
rect 41346 544895 41406 552969
rect 41343 544894 41409 544895
rect 41343 544830 41344 544894
rect 41408 544830 41409 544894
rect 41343 544829 41409 544830
rect 41151 544154 41217 544155
rect 41151 544090 41152 544154
rect 41216 544090 41217 544154
rect 41151 544089 41217 544090
rect 41154 538975 41214 544089
rect 41343 541342 41409 541343
rect 41343 541278 41344 541342
rect 41408 541278 41409 541342
rect 41343 541277 41409 541278
rect 42303 541342 42369 541343
rect 42303 541278 42304 541342
rect 42368 541278 42369 541342
rect 42303 541277 42369 541278
rect 41151 538974 41217 538975
rect 41151 538910 41152 538974
rect 41216 538910 41217 538974
rect 41151 538909 41217 538910
rect 41346 531427 41406 541277
rect 41919 541046 41985 541047
rect 41919 540982 41920 541046
rect 41984 540982 41985 541046
rect 41919 540981 41985 540982
rect 42111 541046 42177 541047
rect 42111 540982 42112 541046
rect 42176 540982 42177 541046
rect 42111 540981 42177 540982
rect 41535 535718 41601 535719
rect 41535 535654 41536 535718
rect 41600 535654 41601 535718
rect 41535 535653 41601 535654
rect 41538 531871 41598 535653
rect 41922 533795 41982 540981
rect 42114 537051 42174 540981
rect 42111 537050 42177 537051
rect 42111 536986 42112 537050
rect 42176 536986 42177 537050
rect 42111 536985 42177 536986
rect 42306 534535 42366 541277
rect 42879 541194 42945 541195
rect 42879 541130 42880 541194
rect 42944 541130 42945 541194
rect 42879 541129 42945 541130
rect 42882 535275 42942 541129
rect 42879 535274 42945 535275
rect 42879 535210 42880 535274
rect 42944 535210 42945 535274
rect 42879 535209 42945 535210
rect 42303 534534 42369 534535
rect 42303 534470 42304 534534
rect 42368 534470 42369 534534
rect 42303 534469 42369 534470
rect 41919 533794 41985 533795
rect 41919 533730 41920 533794
rect 41984 533730 41985 533794
rect 41919 533729 41985 533730
rect 43074 532759 43134 572949
rect 673986 535423 674046 607729
rect 674367 607202 674433 607203
rect 674367 607138 674368 607202
rect 674432 607138 674433 607202
rect 674367 607137 674433 607138
rect 674175 600246 674241 600247
rect 674175 600182 674176 600246
rect 674240 600182 674241 600246
rect 674175 600181 674241 600182
rect 674178 578935 674238 600181
rect 674175 578934 674241 578935
rect 674175 578870 674176 578934
rect 674240 578870 674241 578934
rect 674175 578869 674241 578870
rect 674175 562062 674241 562063
rect 674175 561998 674176 562062
rect 674240 561998 674241 562062
rect 674175 561997 674241 561998
rect 673983 535422 674049 535423
rect 673983 535358 673984 535422
rect 674048 535358 674049 535422
rect 673983 535357 674049 535358
rect 42111 532758 42177 532759
rect 42111 532694 42112 532758
rect 42176 532694 42177 532758
rect 42111 532693 42177 532694
rect 43071 532758 43137 532759
rect 43071 532694 43072 532758
rect 43136 532694 43137 532758
rect 43071 532693 43137 532694
rect 41535 531870 41601 531871
rect 41535 531806 41536 531870
rect 41600 531806 41601 531870
rect 41535 531805 41601 531806
rect 41343 531426 41409 531427
rect 41343 531362 41344 531426
rect 41408 531362 41409 531426
rect 41343 531361 41409 531362
rect 40959 530094 41025 530095
rect 40959 530030 40960 530094
rect 41024 530030 41025 530094
rect 40959 530029 41025 530030
rect 40767 526542 40833 526543
rect 40767 526478 40768 526542
rect 40832 526478 40833 526542
rect 40767 526477 40833 526478
rect 41538 524175 41598 531805
rect 41535 524174 41601 524175
rect 41535 524110 41536 524174
rect 41600 524110 41601 524174
rect 41535 524109 41601 524110
rect 42114 510115 42174 532693
rect 42111 510114 42177 510115
rect 42111 510050 42112 510114
rect 42176 510050 42177 510114
rect 42111 510049 42177 510050
rect 41727 504046 41793 504047
rect 41727 503982 41728 504046
rect 41792 503982 41793 504046
rect 41727 503981 41793 503982
rect 42111 504046 42177 504047
rect 42111 503982 42112 504046
rect 42176 503982 42177 504046
rect 42111 503981 42177 503982
rect 41730 491023 41790 503981
rect 41727 491022 41793 491023
rect 41727 490958 41728 491022
rect 41792 490958 41793 491022
rect 41727 490957 41793 490958
rect 42114 489691 42174 503981
rect 42111 489690 42177 489691
rect 42111 489626 42112 489690
rect 42176 489626 42177 489690
rect 42111 489625 42177 489626
rect 42303 489394 42369 489395
rect 42303 489330 42304 489394
rect 42368 489330 42369 489394
rect 42303 489329 42369 489330
rect 42306 483771 42366 489329
rect 674178 487767 674238 561997
rect 674370 531723 674430 607137
rect 674562 577307 674622 652129
rect 674943 651454 675009 651455
rect 674943 651390 674944 651454
rect 675008 651390 675009 651454
rect 674943 651389 675009 651390
rect 674751 648938 674817 648939
rect 674751 648874 674752 648938
rect 674816 648874 674817 648938
rect 674751 648873 674817 648874
rect 674559 577306 674625 577307
rect 674559 577242 674560 577306
rect 674624 577242 674625 577306
rect 674559 577241 674625 577242
rect 674754 576123 674814 648873
rect 674946 581747 675006 651389
rect 675138 619191 675198 689129
rect 675330 665959 675390 738561
rect 675522 712727 675582 787105
rect 675714 715835 675774 787993
rect 675903 784802 675969 784803
rect 675903 784738 675904 784802
rect 675968 784738 675969 784802
rect 675903 784737 675969 784738
rect 675711 715834 675777 715835
rect 675711 715770 675712 715834
rect 675776 715770 675777 715834
rect 675711 715769 675777 715770
rect 675906 715095 675966 784737
rect 676098 760531 676158 876941
rect 676671 864722 676737 864723
rect 676671 864658 676672 864722
rect 676736 864658 676737 864722
rect 676671 864657 676737 864658
rect 676479 786726 676545 786727
rect 676479 786662 676480 786726
rect 676544 786662 676545 786726
rect 676479 786661 676545 786662
rect 676287 775478 676353 775479
rect 676287 775414 676288 775478
rect 676352 775414 676353 775478
rect 676287 775413 676353 775414
rect 676095 760530 676161 760531
rect 676095 760466 676096 760530
rect 676160 760466 676161 760530
rect 676095 760465 676161 760466
rect 676095 741734 676161 741735
rect 676095 741670 676096 741734
rect 676160 741670 676161 741734
rect 676095 741669 676161 741670
rect 675903 715094 675969 715095
rect 675903 715030 675904 715094
rect 675968 715030 675969 715094
rect 675903 715029 675969 715030
rect 675519 712726 675585 712727
rect 675519 712662 675520 712726
rect 675584 712662 675585 712726
rect 675519 712661 675585 712662
rect 675519 697926 675585 697927
rect 675519 697862 675520 697926
rect 675584 697862 675585 697926
rect 675519 697861 675585 697862
rect 675327 665958 675393 665959
rect 675327 665894 675328 665958
rect 675392 665894 675393 665958
rect 675327 665893 675393 665894
rect 675327 652638 675393 652639
rect 675327 652574 675328 652638
rect 675392 652574 675393 652638
rect 675327 652573 675393 652574
rect 675135 619190 675201 619191
rect 675135 619126 675136 619190
rect 675200 619126 675201 619190
rect 675135 619125 675201 619126
rect 675135 604834 675201 604835
rect 675135 604770 675136 604834
rect 675200 604770 675201 604834
rect 675135 604769 675201 604770
rect 674943 581746 675009 581747
rect 674943 581682 674944 581746
rect 675008 581682 675009 581746
rect 674943 581681 675009 581682
rect 674751 576122 674817 576123
rect 674751 576058 674752 576122
rect 674816 576058 674817 576122
rect 674751 576057 674817 576058
rect 674943 568722 675009 568723
rect 674943 568658 674944 568722
rect 675008 568658 675009 568722
rect 674943 568657 675009 568658
rect 674946 558955 675006 568657
rect 674943 558954 675009 558955
rect 674943 558890 674944 558954
rect 675008 558890 675009 558954
rect 674943 558889 675009 558890
rect 674943 558806 675009 558807
rect 674943 558742 674944 558806
rect 675008 558742 675009 558806
rect 674943 558741 675009 558742
rect 674559 558214 674625 558215
rect 674559 558150 674560 558214
rect 674624 558150 674625 558214
rect 674559 558149 674625 558150
rect 674367 531722 674433 531723
rect 674367 531658 674368 531722
rect 674432 531658 674433 531722
rect 674367 531657 674433 531658
rect 674175 487766 674241 487767
rect 674175 487702 674176 487766
rect 674240 487702 674241 487766
rect 674175 487701 674241 487702
rect 674562 486731 674622 558149
rect 674751 554514 674817 554515
rect 674751 554450 674752 554514
rect 674816 554450 674817 554514
rect 674751 554449 674817 554450
rect 674559 486730 674625 486731
rect 674559 486666 674560 486730
rect 674624 486666 674625 486730
rect 674559 486665 674625 486666
rect 42303 483770 42369 483771
rect 42303 483706 42304 483770
rect 42368 483706 42369 483770
rect 42303 483705 42369 483706
rect 42687 483770 42753 483771
rect 42687 483706 42688 483770
rect 42752 483706 42753 483770
rect 42687 483705 42753 483706
rect 41919 481106 41985 481107
rect 41919 481042 41920 481106
rect 41984 481042 41985 481106
rect 41919 481041 41985 481042
rect 41922 463939 41982 481041
rect 42690 468561 42750 483705
rect 674754 483623 674814 554449
rect 674946 487471 675006 558741
rect 675138 534683 675198 604769
rect 675330 580415 675390 652573
rect 675522 638727 675582 697861
rect 675903 697186 675969 697187
rect 675903 697122 675904 697186
rect 675968 697122 675969 697186
rect 675903 697121 675969 697122
rect 675711 694818 675777 694819
rect 675711 694754 675712 694818
rect 675776 694754 675777 694818
rect 675711 694753 675777 694754
rect 675714 641055 675774 694753
rect 675906 645717 675966 697121
rect 676098 672323 676158 741669
rect 676290 716723 676350 775413
rect 676482 717167 676542 786661
rect 676674 761715 676734 864657
rect 676863 779178 676929 779179
rect 676863 779114 676864 779178
rect 676928 779114 676929 779178
rect 676863 779113 676929 779114
rect 676671 761714 676737 761715
rect 676671 761650 676672 761714
rect 676736 761650 676737 761714
rect 676671 761649 676737 761650
rect 676671 742474 676737 742475
rect 676671 742410 676672 742474
rect 676736 742410 676737 742474
rect 676671 742409 676737 742410
rect 676479 717166 676545 717167
rect 676479 717102 676480 717166
rect 676544 717102 676545 717166
rect 676479 717101 676545 717102
rect 676287 716722 676353 716723
rect 676287 716658 676288 716722
rect 676352 716658 676353 716722
rect 676287 716657 676353 716658
rect 676479 697334 676545 697335
rect 676479 697270 676480 697334
rect 676544 697270 676545 697334
rect 676479 697269 676545 697270
rect 676287 691710 676353 691711
rect 676287 691646 676288 691710
rect 676352 691646 676353 691710
rect 676287 691645 676353 691646
rect 676095 672322 676161 672323
rect 676095 672258 676096 672322
rect 676160 672258 676161 672322
rect 676095 672257 676161 672258
rect 676290 653675 676350 691645
rect 676287 653674 676353 653675
rect 676287 653610 676288 653674
rect 676352 653610 676353 653674
rect 676287 653609 676353 653610
rect 675906 645657 676350 645717
rect 676095 645386 676161 645387
rect 676095 645322 676096 645386
rect 676160 645322 676161 645386
rect 676095 645321 676161 645322
rect 675714 640995 675966 641055
rect 675906 639911 675966 640995
rect 675903 639910 675969 639911
rect 675903 639846 675904 639910
rect 675968 639846 675969 639910
rect 675903 639845 675969 639846
rect 675711 639466 675777 639467
rect 675711 639402 675712 639466
rect 675776 639402 675777 639466
rect 675711 639401 675777 639402
rect 675519 638726 675585 638727
rect 675519 638662 675520 638726
rect 675584 638662 675585 638726
rect 675519 638661 675585 638662
rect 675519 638578 675585 638579
rect 675519 638514 675520 638578
rect 675584 638514 675585 638578
rect 675519 638513 675585 638514
rect 675327 580414 675393 580415
rect 675327 580350 675328 580414
rect 675392 580350 675393 580414
rect 675327 580349 675393 580350
rect 675522 578195 675582 638513
rect 675714 630883 675774 639401
rect 675711 630882 675777 630883
rect 675711 630818 675712 630882
rect 675776 630818 675777 630882
rect 675711 630817 675777 630818
rect 675903 630882 675969 630883
rect 675903 630818 675904 630882
rect 675968 630818 675969 630882
rect 675903 630817 675969 630818
rect 675711 630438 675777 630439
rect 675711 630374 675712 630438
rect 675776 630374 675777 630438
rect 675711 630373 675777 630374
rect 675714 624815 675774 630373
rect 675906 625703 675966 630817
rect 675903 625702 675969 625703
rect 675903 625638 675904 625702
rect 675968 625638 675969 625702
rect 675903 625637 675969 625638
rect 675711 624814 675777 624815
rect 675711 624750 675712 624814
rect 675776 624750 675777 624814
rect 675711 624749 675777 624750
rect 675711 606462 675777 606463
rect 675711 606398 675712 606462
rect 675776 606398 675777 606462
rect 675711 606397 675777 606398
rect 675519 578194 675585 578195
rect 675519 578130 675520 578194
rect 675584 578130 675585 578194
rect 675519 578129 675585 578130
rect 675327 562506 675393 562507
rect 675327 562442 675328 562506
rect 675392 562442 675393 562506
rect 675327 562441 675393 562442
rect 675135 534682 675201 534683
rect 675135 534618 675136 534682
rect 675200 534618 675201 534682
rect 675135 534617 675201 534618
rect 675330 491467 675390 562441
rect 675519 561766 675585 561767
rect 675519 561702 675520 561766
rect 675584 561702 675585 561766
rect 675519 561701 675585 561702
rect 675522 492799 675582 561701
rect 675714 537051 675774 606397
rect 676098 595767 676158 645321
rect 676290 627331 676350 645657
rect 676287 627330 676353 627331
rect 676287 627266 676288 627330
rect 676352 627266 676353 627330
rect 676287 627265 676353 627266
rect 676482 622151 676542 697269
rect 676674 667587 676734 742409
rect 676866 709471 676926 779113
rect 677058 777551 677310 777585
rect 677055 777550 677310 777551
rect 677055 777486 677056 777550
rect 677120 777525 677310 777550
rect 677120 777486 677121 777525
rect 677055 777485 677121 777486
rect 677055 777402 677121 777403
rect 677055 777338 677056 777402
rect 677120 777338 677121 777402
rect 677055 777337 677121 777338
rect 677058 731819 677118 777337
rect 677250 754463 677310 777525
rect 677823 773110 677889 773111
rect 677823 773046 677824 773110
rect 677888 773046 677889 773110
rect 677823 773045 677889 773046
rect 677826 755351 677886 773045
rect 677823 755350 677889 755351
rect 677823 755286 677824 755350
rect 677888 755286 677889 755350
rect 677823 755285 677889 755286
rect 677247 754462 677313 754463
rect 677247 754398 677248 754462
rect 677312 754398 677313 754462
rect 677247 754397 677313 754398
rect 677055 731818 677121 731819
rect 677055 731754 677056 731818
rect 677120 731754 677121 731818
rect 677055 731753 677121 731754
rect 677823 728118 677889 728119
rect 677823 728054 677824 728118
rect 677888 728054 677889 728118
rect 677823 728053 677889 728054
rect 677055 727970 677121 727971
rect 677055 727906 677056 727970
rect 677120 727906 677121 727970
rect 677055 727905 677121 727906
rect 676863 709470 676929 709471
rect 676863 709406 676864 709470
rect 676928 709406 676929 709470
rect 676863 709405 676929 709406
rect 676863 687566 676929 687567
rect 676863 687502 676864 687566
rect 676928 687502 676929 687566
rect 676863 687501 676929 687502
rect 676671 667586 676737 667587
rect 676671 667522 676672 667586
rect 676736 667522 676737 667586
rect 676671 667521 676737 667522
rect 676671 649826 676737 649827
rect 676671 649762 676672 649826
rect 676736 649762 676737 649826
rect 676671 649761 676737 649762
rect 676479 622150 676545 622151
rect 676479 622086 676480 622150
rect 676544 622086 676545 622150
rect 676479 622085 676545 622086
rect 676287 613418 676353 613419
rect 676287 613354 676288 613418
rect 676352 613354 676353 613418
rect 676287 613353 676353 613354
rect 676290 596433 676350 613353
rect 676290 596373 676542 596433
rect 676098 595707 676350 595767
rect 675903 593586 675969 593587
rect 675903 593522 675904 593586
rect 675968 593522 675969 593586
rect 675903 593521 675969 593522
rect 675906 579675 675966 593521
rect 675903 579674 675969 579675
rect 675903 579610 675904 579674
rect 675968 579610 675969 579674
rect 675903 579609 675969 579610
rect 675903 578934 675969 578935
rect 675903 578870 675904 578934
rect 675968 578870 675969 578934
rect 675903 578869 675969 578870
rect 675711 537050 675777 537051
rect 675711 536986 675712 537050
rect 675776 536986 675777 537050
rect 675711 536985 675777 536986
rect 675906 533795 675966 578869
rect 676290 578787 676350 595707
rect 676482 581303 676542 596373
rect 676674 593587 676734 649761
rect 676866 617859 676926 687501
rect 677058 663591 677118 727905
rect 677826 710359 677886 728053
rect 677823 710358 677889 710359
rect 677823 710294 677824 710358
rect 677888 710294 677889 710358
rect 677823 710293 677889 710294
rect 677055 663590 677121 663591
rect 677055 663526 677056 663590
rect 677120 663526 677121 663590
rect 677055 663525 677121 663526
rect 676863 617858 676929 617859
rect 676863 617794 676864 617858
rect 676928 617794 676929 617858
rect 676863 617793 676929 617794
rect 676671 593586 676737 593587
rect 676671 593522 676672 593586
rect 676736 593522 676737 593586
rect 676671 593521 676737 593522
rect 676863 593438 676929 593439
rect 676863 593374 676864 593438
rect 676928 593374 676929 593438
rect 676863 593373 676929 593374
rect 676479 581302 676545 581303
rect 676479 581238 676480 581302
rect 676544 581238 676545 581302
rect 676479 581237 676545 581238
rect 676866 581115 676926 593373
rect 676482 581055 676926 581115
rect 676287 578786 676353 578787
rect 676287 578722 676288 578786
rect 676352 578722 676353 578786
rect 676287 578721 676353 578722
rect 676287 558806 676353 558807
rect 676287 558742 676288 558806
rect 676352 558742 676353 558806
rect 676287 558741 676353 558742
rect 676290 536311 676350 558741
rect 676482 550223 676542 581055
rect 676863 557622 676929 557623
rect 676863 557558 676864 557622
rect 676928 557558 676929 557622
rect 676863 557557 676929 557558
rect 676479 550222 676545 550223
rect 676479 550158 676480 550222
rect 676544 550158 676545 550222
rect 676479 550157 676545 550158
rect 676671 549926 676737 549927
rect 676671 549862 676672 549926
rect 676736 549862 676737 549926
rect 676671 549861 676737 549862
rect 676287 536310 676353 536311
rect 676287 536246 676288 536310
rect 676352 536246 676353 536310
rect 676287 536245 676353 536246
rect 675903 533794 675969 533795
rect 675903 533730 675904 533794
rect 675968 533730 675969 533794
rect 675903 533729 675969 533730
rect 676674 532759 676734 549861
rect 676671 532758 676737 532759
rect 676671 532694 676672 532758
rect 676736 532694 676737 532758
rect 676671 532693 676737 532694
rect 675519 492798 675585 492799
rect 675519 492734 675520 492798
rect 675584 492734 675585 492798
rect 675519 492733 675585 492734
rect 675327 491466 675393 491467
rect 675327 491402 675328 491466
rect 675392 491402 675393 491466
rect 675327 491401 675393 491402
rect 674943 487470 675009 487471
rect 674943 487406 674944 487470
rect 675008 487406 675009 487470
rect 674943 487405 675009 487406
rect 676866 484067 676926 557557
rect 676863 484066 676929 484067
rect 676863 484002 676864 484066
rect 676928 484002 676929 484066
rect 676863 484001 676929 484002
rect 674751 483622 674817 483623
rect 674751 483558 674752 483622
rect 674816 483558 674817 483622
rect 674751 483557 674817 483558
rect 42306 468501 42750 468561
rect 41919 463938 41985 463939
rect 41919 463874 41920 463938
rect 41984 463874 41985 463938
rect 41919 463873 41985 463874
rect 41727 463790 41793 463791
rect 41727 463726 41728 463790
rect 41792 463726 41793 463790
rect 41727 463725 41793 463726
rect 40383 432710 40449 432711
rect 40383 432646 40384 432710
rect 40448 432646 40449 432710
rect 40383 432645 40449 432646
rect 40386 390235 40446 432645
rect 40575 431970 40641 431971
rect 40575 431906 40576 431970
rect 40640 431906 40641 431970
rect 40575 431905 40641 431906
rect 40383 390234 40449 390235
rect 40383 390170 40384 390234
rect 40448 390170 40449 390234
rect 40383 390169 40449 390170
rect 40386 346871 40446 390169
rect 40578 389199 40638 431905
rect 40767 430786 40833 430787
rect 40767 430722 40768 430786
rect 40832 430722 40833 430786
rect 40767 430721 40833 430722
rect 40770 400151 40830 430721
rect 40959 429454 41025 429455
rect 40959 429390 40960 429454
rect 41024 429390 41025 429454
rect 40959 429389 41025 429390
rect 40767 400150 40833 400151
rect 40767 400086 40768 400150
rect 40832 400086 40833 400150
rect 40767 400085 40833 400086
rect 40962 398819 41022 429389
rect 41343 428418 41409 428419
rect 41343 428354 41344 428418
rect 41408 428354 41409 428418
rect 41343 428353 41409 428354
rect 41151 426346 41217 426347
rect 41151 426282 41152 426346
rect 41216 426282 41217 426346
rect 41151 426281 41217 426282
rect 41154 399559 41214 426281
rect 41346 401927 41406 428353
rect 41535 425162 41601 425163
rect 41535 425098 41536 425162
rect 41600 425098 41601 425162
rect 41535 425097 41601 425098
rect 41538 402667 41598 425097
rect 41730 403703 41790 463725
rect 42306 448581 42366 468501
rect 41922 448521 42366 448581
rect 41922 427935 41982 448521
rect 41922 427875 42366 427935
rect 42111 427678 42177 427679
rect 42111 427614 42112 427678
rect 42176 427614 42177 427678
rect 42111 427613 42177 427614
rect 42114 423239 42174 427613
rect 42111 423238 42177 423239
rect 42111 423174 42112 423238
rect 42176 423174 42177 423238
rect 42111 423173 42177 423174
rect 42111 423090 42177 423091
rect 42111 423026 42112 423090
rect 42176 423026 42177 423090
rect 42111 423025 42177 423026
rect 42114 406367 42174 423025
rect 42306 409179 42366 427875
rect 676479 412138 676545 412139
rect 676479 412074 676480 412138
rect 676544 412074 676545 412138
rect 676479 412073 676545 412074
rect 42303 409178 42369 409179
rect 42303 409114 42304 409178
rect 42368 409114 42369 409178
rect 42303 409113 42369 409114
rect 42495 408882 42561 408883
rect 42495 408818 42496 408882
rect 42560 408818 42561 408882
rect 42495 408817 42561 408818
rect 42111 406366 42177 406367
rect 42111 406302 42112 406366
rect 42176 406302 42177 406366
rect 42111 406301 42177 406302
rect 42498 405183 42558 408817
rect 676482 406219 676542 412073
rect 676671 411990 676737 411991
rect 676671 411926 676672 411990
rect 676736 411926 676737 411990
rect 676671 411925 676737 411926
rect 676479 406218 676545 406219
rect 676479 406154 676480 406218
rect 676544 406154 676545 406218
rect 676479 406153 676545 406154
rect 674175 405922 674241 405923
rect 674175 405858 674176 405922
rect 674240 405858 674241 405922
rect 674175 405857 674241 405858
rect 42495 405182 42561 405183
rect 42495 405118 42496 405182
rect 42560 405118 42561 405182
rect 42495 405117 42561 405118
rect 41727 403702 41793 403703
rect 41727 403638 41728 403702
rect 41792 403638 41793 403702
rect 41727 403637 41793 403638
rect 41535 402666 41601 402667
rect 41535 402602 41536 402666
rect 41600 402602 41601 402666
rect 41535 402601 41601 402602
rect 41343 401926 41409 401927
rect 41343 401862 41344 401926
rect 41408 401862 41409 401926
rect 41343 401861 41409 401862
rect 41151 399558 41217 399559
rect 41151 399494 41152 399558
rect 41216 399494 41217 399558
rect 41151 399493 41217 399494
rect 40959 398818 41025 398819
rect 40959 398754 40960 398818
rect 41024 398754 41025 398818
rect 40959 398753 41025 398754
rect 40575 389198 40641 389199
rect 40575 389134 40576 389198
rect 40640 389134 40641 389198
rect 40575 389133 40641 389134
rect 40383 346870 40449 346871
rect 40383 346806 40384 346870
rect 40448 346806 40449 346870
rect 40383 346805 40449 346806
rect 40386 303803 40446 346805
rect 40578 346279 40638 389133
rect 40767 387570 40833 387571
rect 40767 387506 40768 387570
rect 40832 387506 40833 387570
rect 40767 387505 40833 387506
rect 40770 356935 40830 387505
rect 40959 386090 41025 386091
rect 40959 386026 40960 386090
rect 41024 386026 41025 386090
rect 40959 386025 41025 386026
rect 40767 356934 40833 356935
rect 40767 356870 40768 356934
rect 40832 356870 40833 356934
rect 40767 356869 40833 356870
rect 40962 355603 41022 386025
rect 41343 385202 41409 385203
rect 41343 385138 41344 385202
rect 41408 385138 41409 385202
rect 41343 385137 41409 385138
rect 41151 383130 41217 383131
rect 41151 383066 41152 383130
rect 41216 383066 41217 383130
rect 41151 383065 41217 383066
rect 41154 356491 41214 383065
rect 41346 358711 41406 385137
rect 41535 381946 41601 381947
rect 41535 381882 41536 381946
rect 41600 381882 41601 381946
rect 41535 381881 41601 381882
rect 41538 359451 41598 381881
rect 41730 360635 41790 403637
rect 41919 403258 41985 403259
rect 41919 403194 41920 403258
rect 41984 403194 41985 403258
rect 41919 403193 41985 403194
rect 41922 361967 41982 403193
rect 42111 384462 42177 384463
rect 42111 384398 42112 384462
rect 42176 384398 42177 384462
rect 42111 384397 42177 384398
rect 42114 362855 42174 384397
rect 42303 370550 42369 370551
rect 42303 370486 42304 370550
rect 42368 370486 42369 370550
rect 42303 370485 42369 370486
rect 42111 362854 42177 362855
rect 42111 362790 42112 362854
rect 42176 362790 42177 362854
rect 42111 362789 42177 362790
rect 41919 361966 41985 361967
rect 41919 361902 41920 361966
rect 41984 361902 41985 361966
rect 41919 361901 41985 361902
rect 41727 360634 41793 360635
rect 41727 360570 41728 360634
rect 41792 360570 41793 360634
rect 41727 360569 41793 360570
rect 41535 359450 41601 359451
rect 41535 359386 41536 359450
rect 41600 359386 41601 359450
rect 41535 359385 41601 359386
rect 41343 358710 41409 358711
rect 41343 358646 41344 358710
rect 41408 358646 41409 358710
rect 41343 358645 41409 358646
rect 41151 356490 41217 356491
rect 41151 356426 41152 356490
rect 41216 356426 41217 356490
rect 41151 356425 41217 356426
rect 40959 355602 41025 355603
rect 40959 355538 40960 355602
rect 41024 355538 41025 355602
rect 40959 355537 41025 355538
rect 40575 346278 40641 346279
rect 40575 346214 40576 346278
rect 40640 346214 40641 346278
rect 40575 346213 40641 346214
rect 40383 303802 40449 303803
rect 40383 303738 40384 303802
rect 40448 303738 40449 303802
rect 40383 303737 40449 303738
rect 40578 303063 40638 346213
rect 40959 344354 41025 344355
rect 40959 344290 40960 344354
rect 41024 344290 41025 344354
rect 40959 344289 41025 344290
rect 40767 342874 40833 342875
rect 40767 342810 40768 342874
rect 40832 342810 40833 342874
rect 40767 342809 40833 342810
rect 40770 312387 40830 342809
rect 40962 313719 41022 344289
rect 41151 341986 41217 341987
rect 41151 341922 41152 341986
rect 41216 341922 41217 341986
rect 41151 341921 41217 341922
rect 41154 315495 41214 341921
rect 41343 338730 41409 338731
rect 41343 338666 41344 338730
rect 41408 338666 41409 338730
rect 41343 338665 41409 338666
rect 41346 316087 41406 338665
rect 41535 336510 41601 336511
rect 41535 336446 41536 336510
rect 41600 336446 41601 336510
rect 41535 336445 41601 336446
rect 41343 316086 41409 316087
rect 41343 316022 41344 316086
rect 41408 316022 41409 316086
rect 41343 316021 41409 316022
rect 41151 315494 41217 315495
rect 41151 315430 41152 315494
rect 41216 315430 41217 315494
rect 41151 315429 41217 315430
rect 40959 313718 41025 313719
rect 40959 313654 40960 313718
rect 41024 313654 41025 313718
rect 40959 313653 41025 313654
rect 41538 313275 41598 336445
rect 41730 317863 41790 360569
rect 41922 318751 41982 361901
rect 42306 360191 42366 370485
rect 674178 360783 674238 405857
rect 676674 405331 676734 411925
rect 675327 405330 675393 405331
rect 675327 405266 675328 405330
rect 675392 405266 675393 405330
rect 675327 405265 675393 405266
rect 676671 405330 676737 405331
rect 676671 405266 676672 405330
rect 676736 405266 676737 405330
rect 676671 405265 676737 405266
rect 674943 403258 675009 403259
rect 674943 403194 674944 403258
rect 675008 403194 675009 403258
rect 674943 403193 675009 403194
rect 674559 400594 674625 400595
rect 674559 400530 674560 400594
rect 674624 400530 674625 400594
rect 674559 400529 674625 400530
rect 674367 400446 674433 400447
rect 674367 400382 674368 400446
rect 674432 400382 674433 400446
rect 674367 400381 674433 400382
rect 674370 372031 674430 400381
rect 674562 378839 674622 400529
rect 674559 378838 674625 378839
rect 674559 378774 674560 378838
rect 674624 378774 674625 378838
rect 674559 378773 674625 378774
rect 674946 373955 675006 403193
rect 674943 373954 675009 373955
rect 674943 373890 674944 373954
rect 675008 373890 675009 373954
rect 674943 373889 675009 373890
rect 674367 372030 674433 372031
rect 674367 371966 674368 372030
rect 674432 371966 674433 372030
rect 674367 371965 674433 371966
rect 674367 361448 674433 361449
rect 674367 361384 674368 361448
rect 674432 361384 674433 361448
rect 674367 361383 674433 361384
rect 674175 360782 674241 360783
rect 674175 360718 674176 360782
rect 674240 360718 674241 360782
rect 674175 360717 674241 360718
rect 42303 360190 42369 360191
rect 42303 360126 42304 360190
rect 42368 360126 42369 360190
rect 42303 360125 42369 360126
rect 673983 360042 674049 360043
rect 673983 359978 673984 360042
rect 674048 359978 674049 360042
rect 673983 359977 674049 359978
rect 42111 341246 42177 341247
rect 42111 341182 42112 341246
rect 42176 341182 42177 341246
rect 42111 341181 42177 341182
rect 42114 319787 42174 341181
rect 42111 319786 42177 319787
rect 42111 319722 42112 319786
rect 42176 319722 42177 319786
rect 42111 319721 42177 319722
rect 41919 318750 41985 318751
rect 41919 318686 41920 318750
rect 41984 318686 41985 318750
rect 41919 318685 41985 318686
rect 41727 317862 41793 317863
rect 41727 317798 41728 317862
rect 41792 317798 41793 317862
rect 41727 317797 41793 317798
rect 41535 313274 41601 313275
rect 41535 313210 41536 313274
rect 41600 313210 41601 313274
rect 41535 313209 41601 313210
rect 40767 312386 40833 312387
rect 40767 312322 40768 312386
rect 40832 312322 40833 312386
rect 40767 312321 40833 312322
rect 40575 303062 40641 303063
rect 40575 302998 40576 303062
rect 40640 302998 40641 303062
rect 40575 302997 40641 302998
rect 40767 301138 40833 301139
rect 40767 301074 40768 301138
rect 40832 301074 40833 301138
rect 40767 301073 40833 301074
rect 40383 298030 40449 298031
rect 40383 297966 40384 298030
rect 40448 297966 40449 298030
rect 40383 297965 40449 297966
rect 40386 276571 40446 297965
rect 40575 284118 40641 284119
rect 40575 284054 40576 284118
rect 40640 284054 40641 284118
rect 40575 284053 40641 284054
rect 40578 279827 40638 284053
rect 40575 279826 40641 279827
rect 40575 279762 40576 279826
rect 40640 279762 40641 279826
rect 40575 279761 40641 279762
rect 40383 276570 40449 276571
rect 40383 276506 40384 276570
rect 40448 276506 40449 276570
rect 40383 276505 40449 276506
rect 40770 270651 40830 301073
rect 40959 299658 41025 299659
rect 40959 299594 40960 299658
rect 41024 299594 41025 299658
rect 40959 299593 41025 299594
rect 40767 270650 40833 270651
rect 40767 270586 40768 270650
rect 40832 270586 40833 270650
rect 40767 270585 40833 270586
rect 40962 269171 41022 299593
rect 41151 298770 41217 298771
rect 41151 298706 41152 298770
rect 41216 298706 41217 298770
rect 41151 298705 41217 298706
rect 41154 272279 41214 298705
rect 41535 295514 41601 295515
rect 41535 295450 41536 295514
rect 41600 295450 41601 295514
rect 41535 295449 41601 295450
rect 41343 292406 41409 292407
rect 41343 292342 41344 292406
rect 41408 292342 41409 292406
rect 41343 292341 41409 292342
rect 41151 272278 41217 272279
rect 41151 272214 41152 272278
rect 41216 272214 41217 272278
rect 41151 272213 41217 272214
rect 41346 270059 41406 292341
rect 41538 273019 41598 295449
rect 41730 274943 41790 317797
rect 41922 275535 41982 318685
rect 673986 314903 674046 359977
rect 674178 315791 674238 360717
rect 674370 317271 674430 361383
rect 675330 360191 675390 405265
rect 675519 374546 675585 374547
rect 675519 374482 675520 374546
rect 675584 374482 675585 374546
rect 675519 374481 675585 374482
rect 675327 360190 675393 360191
rect 675327 360126 675328 360190
rect 675392 360126 675393 360190
rect 675327 360125 675393 360126
rect 675522 335179 675582 374481
rect 675711 374102 675777 374103
rect 675711 374038 675712 374102
rect 675776 374038 675777 374102
rect 675711 374037 675777 374038
rect 675519 335178 675585 335179
rect 675519 335114 675520 335178
rect 675584 335114 675585 335178
rect 675519 335113 675585 335114
rect 675714 334029 675774 374037
rect 676479 345538 676545 345539
rect 676479 345474 676480 345538
rect 676544 345474 676545 345538
rect 676479 345473 676545 345474
rect 676287 345390 676353 345391
rect 676287 345326 676288 345390
rect 676352 345326 676353 345390
rect 676287 345325 676353 345326
rect 675330 333969 675774 334029
rect 675330 333847 675390 333969
rect 675327 333846 675393 333847
rect 675327 333782 675328 333846
rect 675392 333782 675393 333846
rect 675327 333781 675393 333782
rect 674367 317270 674433 317271
rect 674367 317206 674368 317270
rect 674432 317206 674433 317270
rect 674367 317205 674433 317206
rect 674943 315938 675009 315939
rect 674943 315874 674944 315938
rect 675008 315874 675009 315938
rect 674943 315873 675009 315874
rect 674175 315790 674241 315791
rect 674175 315726 674176 315790
rect 674240 315726 674241 315790
rect 674175 315725 674241 315726
rect 673983 314902 674049 314903
rect 673983 314838 673984 314902
rect 674048 314838 674049 314902
rect 673983 314837 674049 314838
rect 42303 303210 42369 303211
rect 42303 303146 42304 303210
rect 42368 303146 42369 303210
rect 42303 303145 42369 303146
rect 42111 302322 42177 302323
rect 42111 302258 42112 302322
rect 42176 302258 42177 302322
rect 42111 302257 42177 302258
rect 41919 275534 41985 275535
rect 41919 275470 41920 275534
rect 41984 275470 41985 275534
rect 41919 275469 41985 275470
rect 41727 274942 41793 274943
rect 41727 274878 41728 274942
rect 41792 274878 41793 274942
rect 41727 274877 41793 274878
rect 41535 273018 41601 273019
rect 41535 272954 41536 273018
rect 41600 272954 41601 273018
rect 41535 272953 41601 272954
rect 41730 270503 41790 274877
rect 41727 270502 41793 270503
rect 41727 270438 41728 270502
rect 41792 270438 41793 270502
rect 41727 270437 41793 270438
rect 41343 270058 41409 270059
rect 41343 269994 41344 270058
rect 41408 269994 41409 270058
rect 41343 269993 41409 269994
rect 40959 269170 41025 269171
rect 40959 269106 40960 269170
rect 41024 269106 41025 269170
rect 40959 269105 41025 269106
rect 42114 259551 42174 302257
rect 42306 284745 42366 303145
rect 42306 284685 42558 284745
rect 42303 283378 42369 283379
rect 42303 283314 42304 283378
rect 42368 283314 42369 283378
rect 42303 283313 42369 283314
rect 42306 273759 42366 283313
rect 42303 273758 42369 273759
rect 42303 273694 42304 273758
rect 42368 273694 42369 273758
rect 42303 273693 42369 273694
rect 42498 260439 42558 284685
rect 42687 282490 42753 282491
rect 42687 282426 42688 282490
rect 42752 282426 42753 282490
rect 42687 282425 42753 282426
rect 42690 274203 42750 282425
rect 42879 275534 42945 275535
rect 42879 275470 42880 275534
rect 42944 275470 42945 275534
rect 42879 275469 42945 275470
rect 42687 274202 42753 274203
rect 42687 274138 42688 274202
rect 42752 274138 42753 274202
rect 42687 274137 42753 274138
rect 42495 260438 42561 260439
rect 42495 260374 42496 260438
rect 42560 260374 42561 260438
rect 42495 260373 42561 260374
rect 42111 259550 42177 259551
rect 42111 259486 42112 259550
rect 42176 259486 42177 259550
rect 42111 259485 42177 259486
rect 41535 257922 41601 257923
rect 41535 257858 41536 257922
rect 41600 257858 41601 257922
rect 41535 257857 41601 257858
rect 40383 256294 40449 256295
rect 40383 256230 40384 256294
rect 40448 256230 40449 256294
rect 40383 256229 40449 256230
rect 40386 241939 40446 256229
rect 40959 255702 41025 255703
rect 40959 255638 40960 255702
rect 41024 255638 41025 255702
rect 40959 255637 41025 255638
rect 40767 253482 40833 253483
rect 40767 253418 40768 253482
rect 40832 253418 40833 253482
rect 40767 253417 40833 253418
rect 40383 241938 40449 241939
rect 40383 241874 40384 241938
rect 40448 241874 40449 241938
rect 40383 241873 40449 241874
rect 40770 226695 40830 253417
rect 40962 229063 41022 255637
rect 41151 254814 41217 254815
rect 41151 254750 41152 254814
rect 41216 254750 41217 254814
rect 41151 254749 41217 254750
rect 41154 233355 41214 254749
rect 41343 252742 41409 252743
rect 41343 252678 41344 252742
rect 41408 252678 41409 252742
rect 41343 252677 41409 252678
rect 41151 233354 41217 233355
rect 41151 233290 41152 233354
rect 41216 233290 41217 233354
rect 41151 233289 41217 233290
rect 41346 229803 41406 252677
rect 41343 229802 41409 229803
rect 41343 229738 41344 229802
rect 41408 229738 41409 229802
rect 41343 229737 41409 229738
rect 40959 229062 41025 229063
rect 40959 228998 40960 229062
rect 41024 228998 41025 229062
rect 40959 228997 41025 228998
rect 41538 227287 41598 257857
rect 42111 247118 42177 247119
rect 42111 247054 42112 247118
rect 42176 247054 42177 247118
rect 42111 247053 42177 247054
rect 42114 244899 42174 247053
rect 42882 246823 42942 275469
rect 378495 274942 378561 274943
rect 378495 274878 378496 274942
rect 378560 274878 378561 274942
rect 378495 274877 378561 274878
rect 368511 273610 368577 273611
rect 368511 273546 368512 273610
rect 368576 273546 368577 273610
rect 368511 273545 368577 273546
rect 378111 273610 378177 273611
rect 378111 273546 378112 273610
rect 378176 273546 378177 273610
rect 378111 273545 378177 273546
rect 197439 272722 197505 272723
rect 197439 272658 197440 272722
rect 197504 272658 197505 272722
rect 197439 272657 197505 272658
rect 197442 271425 197502 272657
rect 324159 271686 324225 271687
rect 324159 271622 324160 271686
rect 324224 271622 324225 271686
rect 324159 271621 324225 271622
rect 197058 271365 197502 271425
rect 197058 271095 197118 271365
rect 197055 271094 197121 271095
rect 197055 271030 197056 271094
rect 197120 271030 197121 271094
rect 197055 271029 197121 271030
rect 324162 270847 324222 271621
rect 356991 271538 357057 271539
rect 356991 271474 356992 271538
rect 357056 271474 357057 271538
rect 356991 271473 357057 271474
rect 331071 271242 331137 271243
rect 331071 271178 331072 271242
rect 331136 271178 331137 271242
rect 331071 271177 331137 271178
rect 331074 270847 331134 271177
rect 138111 269910 138177 269911
rect 138111 269846 138112 269910
rect 138176 269846 138177 269910
rect 138111 269845 138177 269846
rect 138114 269615 138174 269845
rect 323010 269763 323070 269945
rect 342594 269763 342654 269945
rect 323007 269762 323073 269763
rect 323007 269698 323008 269762
rect 323072 269698 323073 269762
rect 323007 269697 323073 269698
rect 342591 269762 342657 269763
rect 342591 269698 342592 269762
rect 342656 269698 342657 269762
rect 342591 269697 342657 269698
rect 138111 269614 138177 269615
rect 138111 269550 138112 269614
rect 138176 269550 138177 269614
rect 138111 269549 138177 269550
rect 106431 269466 106497 269467
rect 106431 269402 106432 269466
rect 106496 269427 106497 269466
rect 106623 269466 106689 269467
rect 106623 269427 106624 269466
rect 106496 269402 106624 269427
rect 106688 269402 106689 269466
rect 106431 269401 106689 269402
rect 106434 269367 106686 269401
rect 328575 267838 328641 267839
rect 328575 267774 328576 267838
rect 328640 267774 328641 267838
rect 328575 267773 328641 267774
rect 267519 267690 267585 267691
rect 267519 267626 267520 267690
rect 267584 267626 267585 267690
rect 267519 267625 267585 267626
rect 267522 267429 267582 267625
rect 328578 267429 328638 267773
rect 267522 267395 267774 267429
rect 267522 267394 267777 267395
rect 267522 267369 267712 267394
rect 267711 267330 267712 267369
rect 267776 267330 267777 267394
rect 267711 267329 267777 267330
rect 328386 267369 328638 267429
rect 328386 267099 328446 267369
rect 328383 267098 328449 267099
rect 328383 267034 328384 267098
rect 328448 267034 328449 267098
rect 328383 267033 328449 267034
rect 328575 267098 328641 267099
rect 328575 267034 328576 267098
rect 328640 267034 328641 267098
rect 328575 267033 328641 267034
rect 328383 266802 328449 266803
rect 328383 266738 328384 266802
rect 328448 266763 328449 266802
rect 328578 266763 328638 267033
rect 356994 266851 357054 271473
rect 368514 270847 368574 273545
rect 378114 273315 378174 273545
rect 378111 273314 378177 273315
rect 378111 273250 378112 273314
rect 378176 273250 378177 273314
rect 378111 273249 378177 273250
rect 378498 272720 378558 274877
rect 384639 273166 384705 273167
rect 384639 273102 384640 273166
rect 384704 273102 384705 273166
rect 384639 273101 384705 273102
rect 379647 273018 379713 273019
rect 379647 272954 379648 273018
rect 379712 272954 379713 273018
rect 379647 272953 379713 272954
rect 378498 272660 379518 272720
rect 379458 272279 379518 272660
rect 379455 272278 379521 272279
rect 379455 272214 379456 272278
rect 379520 272214 379521 272278
rect 379455 272213 379521 272214
rect 379650 272091 379710 272953
rect 379074 272031 379710 272091
rect 379074 271687 379134 272031
rect 379071 271686 379137 271687
rect 379071 271622 379072 271686
rect 379136 271622 379137 271686
rect 379071 271621 379137 271622
rect 384642 270181 384702 273101
rect 405375 272426 405441 272427
rect 405375 272362 405376 272426
rect 405440 272362 405441 272426
rect 405375 272361 405441 272362
rect 404223 271834 404289 271835
rect 404223 271770 404224 271834
rect 404288 271770 404289 271834
rect 404223 271769 404289 271770
rect 403839 271686 403905 271687
rect 403839 271622 403840 271686
rect 403904 271622 403905 271686
rect 403839 271621 403905 271622
rect 387135 270946 387201 270947
rect 387135 270882 387136 270946
rect 387200 270882 387201 270946
rect 387135 270881 387201 270882
rect 371010 268579 371070 269945
rect 371007 268578 371073 268579
rect 371007 268514 371008 268578
rect 371072 268514 371073 268578
rect 371007 268513 371073 268514
rect 377154 267987 377214 268613
rect 372927 267986 372993 267987
rect 368514 267099 368574 267947
rect 372927 267922 372928 267986
rect 372992 267922 372993 267986
rect 372927 267921 372993 267922
rect 377151 267986 377217 267987
rect 377151 267922 377152 267986
rect 377216 267922 377217 267986
rect 377151 267921 377217 267922
rect 372930 267517 372990 267921
rect 379074 267543 379134 267947
rect 378687 267542 378753 267543
rect 378687 267478 378688 267542
rect 378752 267478 378753 267542
rect 378687 267477 378753 267478
rect 379071 267542 379137 267543
rect 379071 267478 379072 267542
rect 379136 267478 379137 267542
rect 379071 267477 379137 267478
rect 374463 267246 374529 267247
rect 374463 267182 374464 267246
rect 374528 267182 374529 267246
rect 374463 267181 374529 267182
rect 368511 267098 368577 267099
rect 368511 267034 368512 267098
rect 368576 267034 368577 267098
rect 368511 267033 368577 267034
rect 374466 266851 374526 267181
rect 328448 266738 328638 266763
rect 328383 266737 328638 266738
rect 328767 266802 328833 266803
rect 328767 266738 328768 266802
rect 328832 266738 328833 266802
rect 328767 266737 328833 266738
rect 328386 266703 328638 266737
rect 328770 265519 328830 266737
rect 368511 266590 368512 266615
rect 368576 266590 368577 266615
rect 368511 266589 368577 266590
rect 378690 265519 378750 267477
rect 387138 266851 387198 270881
rect 399039 269762 399105 269763
rect 399039 269698 399040 269762
rect 399104 269698 399105 269762
rect 399039 269697 399105 269698
rect 399042 269427 399102 269697
rect 398658 269367 399102 269427
rect 389247 268430 389313 268431
rect 389247 268366 389248 268430
rect 389312 268366 389313 268430
rect 389247 268365 389313 268366
rect 389250 268135 389310 268365
rect 389247 268134 389313 268135
rect 389247 268070 389248 268134
rect 389312 268070 389313 268134
rect 389247 268069 389313 268070
rect 389247 267838 389313 267839
rect 389247 267774 389248 267838
rect 389312 267774 389313 267838
rect 389247 267773 389313 267774
rect 389055 267542 389121 267543
rect 389055 267478 389056 267542
rect 389120 267478 389121 267542
rect 389055 267477 389121 267478
rect 388290 267099 388350 267281
rect 388095 267098 388161 267099
rect 388095 267034 388096 267098
rect 388160 267096 388161 267098
rect 388287 267098 388353 267099
rect 388160 267034 388206 267096
rect 388095 267033 388206 267034
rect 388287 267034 388288 267098
rect 388352 267034 388353 267098
rect 388287 267033 388353 267034
rect 388146 266948 388206 267033
rect 388146 266888 388542 266948
rect 388482 266504 388542 266888
rect 389058 266803 389118 267477
rect 389055 266802 389121 266803
rect 389055 266738 389056 266802
rect 389120 266738 389121 266802
rect 389055 266737 389121 266738
rect 389250 266652 389310 267773
rect 389442 266951 389502 268613
rect 398658 268579 398718 269367
rect 398655 268578 398721 268579
rect 398655 268514 398656 268578
rect 398720 268514 398721 268578
rect 398655 268513 398721 268514
rect 401151 268430 401217 268431
rect 401151 268366 401152 268430
rect 401216 268366 401217 268430
rect 401151 268365 401217 268366
rect 396735 267986 396801 267987
rect 396735 267922 396736 267986
rect 396800 267922 396801 267986
rect 396735 267921 396801 267922
rect 400383 267986 400449 267987
rect 400383 267922 400384 267986
rect 400448 267922 400449 267986
rect 400383 267921 400449 267922
rect 396738 267395 396798 267921
rect 396735 267394 396801 267395
rect 396735 267330 396736 267394
rect 396800 267330 396801 267394
rect 396735 267329 396801 267330
rect 389439 266950 389505 266951
rect 389439 266886 389440 266950
rect 389504 266886 389505 266950
rect 389439 266885 389505 266886
rect 389631 266802 389697 266803
rect 389631 266738 389632 266802
rect 389696 266738 389697 266802
rect 389631 266737 389697 266738
rect 389439 266654 389505 266655
rect 389439 266652 389440 266654
rect 389250 266592 389440 266652
rect 389439 266590 389440 266592
rect 389504 266590 389505 266654
rect 389439 266589 389505 266590
rect 389634 266504 389694 266737
rect 399999 266654 400065 266655
rect 399999 266590 400000 266654
rect 400064 266590 400065 266654
rect 399999 266589 400065 266590
rect 400191 266654 400257 266655
rect 400191 266590 400192 266654
rect 400256 266590 400257 266654
rect 400191 266589 400257 266590
rect 388482 266444 389694 266504
rect 325506 264990 325566 265283
rect 365058 264990 365118 265283
rect 325503 264989 325569 264990
rect 325503 264925 325504 264989
rect 325568 264925 325569 264989
rect 325503 264924 325569 264925
rect 365055 264989 365121 264990
rect 365055 264925 365056 264989
rect 365120 264925 365121 264989
rect 365055 264924 365121 264925
rect 42879 246822 42945 246823
rect 42879 246758 42880 246822
rect 42944 246758 42945 246822
rect 42879 246757 42945 246758
rect 247551 246822 247617 246823
rect 247551 246758 247552 246822
rect 247616 246758 247617 246822
rect 247551 246757 247617 246758
rect 360063 246822 360129 246823
rect 360063 246758 360064 246822
rect 360128 246783 360129 246822
rect 360447 246822 360513 246823
rect 360447 246783 360448 246822
rect 360128 246758 360448 246783
rect 360512 246758 360513 246822
rect 360063 246757 360513 246758
rect 367743 246822 367809 246823
rect 367743 246758 367744 246822
rect 367808 246758 367809 246822
rect 367743 246757 367809 246758
rect 368511 246822 368577 246823
rect 368511 246758 368512 246822
rect 368576 246758 368577 246822
rect 368511 246757 368577 246758
rect 369279 246822 369345 246823
rect 369279 246758 369280 246822
rect 369344 246758 369345 246822
rect 369279 246757 369345 246758
rect 42111 244898 42177 244899
rect 42111 244834 42112 244898
rect 42176 244834 42177 244898
rect 42111 244833 42177 244834
rect 41919 242678 41985 242679
rect 41919 242614 41920 242678
rect 41984 242614 41985 242678
rect 41919 242613 41985 242614
rect 41727 242086 41793 242087
rect 41727 242022 41728 242086
rect 41792 242022 41793 242086
rect 41727 242021 41793 242022
rect 41730 230395 41790 242021
rect 41922 231727 41982 242613
rect 41919 231726 41985 231727
rect 41919 231662 41920 231726
rect 41984 231662 41985 231726
rect 41919 231661 41985 231662
rect 41727 230394 41793 230395
rect 41727 230330 41728 230394
rect 41792 230330 41793 230394
rect 41727 230329 41793 230330
rect 41727 230246 41793 230247
rect 41727 230182 41728 230246
rect 41792 230182 41793 230246
rect 41727 230181 41793 230182
rect 41535 227286 41601 227287
rect 41535 227222 41536 227286
rect 41600 227222 41601 227286
rect 41535 227221 41601 227222
rect 40767 226694 40833 226695
rect 40767 226630 40768 226694
rect 40832 226630 40833 226694
rect 40767 226629 40833 226630
rect 40383 214706 40449 214707
rect 40383 214642 40384 214706
rect 40448 214642 40449 214706
rect 40383 214641 40449 214642
rect 40386 184219 40446 214641
rect 40575 213226 40641 213227
rect 40575 213162 40576 213226
rect 40640 213162 40641 213226
rect 40575 213161 40641 213162
rect 40383 184218 40449 184219
rect 40383 184154 40384 184218
rect 40448 184154 40449 184218
rect 40383 184153 40449 184154
rect 40578 182887 40638 213161
rect 40959 212486 41025 212487
rect 40959 212422 40960 212486
rect 41024 212422 41025 212486
rect 40959 212421 41025 212422
rect 40767 210414 40833 210415
rect 40767 210350 40768 210414
rect 40832 210350 40833 210414
rect 40767 210349 40833 210350
rect 40770 183627 40830 210349
rect 40962 185995 41022 212421
rect 41151 211598 41217 211599
rect 41151 211534 41152 211598
rect 41216 211534 41217 211598
rect 41151 211533 41217 211534
rect 41154 190139 41214 211533
rect 41343 198722 41409 198723
rect 41343 198658 41344 198722
rect 41408 198658 41409 198722
rect 41343 198657 41409 198658
rect 41346 191027 41406 198657
rect 41343 191026 41409 191027
rect 41343 190962 41344 191026
rect 41408 190962 41409 191026
rect 41343 190961 41409 190962
rect 41151 190138 41217 190139
rect 41151 190074 41152 190138
rect 41216 190074 41217 190138
rect 41151 190073 41217 190074
rect 41730 188363 41790 230181
rect 41922 189103 41982 231661
rect 42114 230987 42174 244833
rect 42882 242679 42942 246757
rect 247554 245451 247614 246757
rect 360066 246723 360510 246757
rect 247362 245391 247614 245451
rect 210303 245194 210369 245195
rect 210303 245130 210304 245194
rect 210368 245130 210369 245194
rect 210303 245129 210369 245130
rect 42879 242678 42945 242679
rect 42879 242614 42880 242678
rect 42944 242614 42945 242678
rect 42879 242613 42945 242614
rect 42303 241938 42369 241939
rect 42303 241874 42304 241938
rect 42368 241874 42369 241938
rect 42303 241873 42369 241874
rect 42111 230986 42177 230987
rect 42111 230922 42112 230986
rect 42176 230922 42177 230986
rect 42111 230921 42177 230922
rect 42306 226251 42366 241873
rect 145407 239866 145473 239867
rect 145407 239802 145408 239866
rect 145472 239802 145473 239866
rect 145407 239801 145473 239802
rect 42303 226250 42369 226251
rect 42303 226186 42304 226250
rect 42368 226186 42369 226250
rect 42303 226185 42369 226186
rect 42303 197538 42369 197539
rect 42303 197474 42304 197538
rect 42368 197474 42369 197538
rect 42303 197473 42369 197474
rect 42306 195171 42366 197473
rect 42303 195170 42369 195171
rect 42303 195106 42304 195170
rect 42368 195106 42369 195170
rect 42303 195105 42369 195106
rect 41919 189102 41985 189103
rect 41919 189038 41920 189102
rect 41984 189038 41985 189102
rect 41919 189037 41985 189038
rect 41727 188362 41793 188363
rect 41727 188298 41728 188362
rect 41792 188298 41793 188362
rect 41727 188297 41793 188298
rect 40959 185994 41025 185995
rect 40959 185930 40960 185994
rect 41024 185930 41025 185994
rect 40959 185929 41025 185930
rect 40767 183626 40833 183627
rect 40767 183562 40768 183626
rect 40832 183562 40833 183626
rect 40767 183561 40833 183562
rect 40575 182886 40641 182887
rect 40575 182822 40576 182886
rect 40640 182822 40641 182886
rect 40575 182821 40641 182822
rect 144447 106518 144513 106519
rect 144447 106454 144448 106518
rect 144512 106454 144513 106518
rect 144447 106453 144513 106454
rect 144450 103707 144510 106453
rect 144447 103706 144513 103707
rect 144447 103642 144448 103706
rect 144512 103642 144513 103706
rect 144447 103641 144513 103642
rect 144831 66262 144897 66263
rect 144831 66198 144832 66262
rect 144896 66198 144897 66262
rect 144831 66197 144897 66198
rect 144834 64635 144894 66197
rect 144831 64634 144897 64635
rect 144831 64570 144832 64634
rect 144896 64570 144897 64634
rect 144831 64569 144897 64570
rect 145410 51463 145470 239801
rect 210306 236315 210366 245129
rect 247362 244751 247422 245391
rect 247359 244750 247425 244751
rect 247359 244686 247360 244750
rect 247424 244686 247425 244750
rect 247359 244685 247425 244686
rect 328383 244602 328449 244603
rect 328383 244538 328384 244602
rect 328448 244538 328449 244602
rect 328383 244537 328449 244538
rect 328386 244119 328446 244537
rect 367746 244307 367806 246757
rect 368514 245451 368574 246757
rect 368514 245391 368766 245451
rect 368706 244455 368766 245391
rect 369282 244603 369342 246757
rect 388863 245046 388929 245047
rect 388863 244982 388864 245046
rect 388928 244982 388929 245046
rect 388863 244981 388929 244982
rect 369279 244602 369345 244603
rect 369279 244538 369280 244602
rect 369344 244538 369345 244602
rect 369279 244537 369345 244538
rect 368703 244454 368769 244455
rect 368703 244390 368704 244454
rect 368768 244390 368769 244454
rect 368703 244389 368769 244390
rect 367743 244306 367809 244307
rect 367743 244242 367744 244306
rect 367808 244242 367809 244306
rect 367743 244241 367809 244242
rect 328386 244059 328638 244119
rect 328578 243567 328638 244059
rect 388866 244011 388926 244981
rect 400002 244603 400062 266589
rect 399999 244602 400065 244603
rect 399999 244538 400000 244602
rect 400064 244538 400065 244602
rect 399999 244537 400065 244538
rect 400194 244455 400254 266589
rect 400191 244454 400257 244455
rect 400191 244390 400192 244454
rect 400256 244390 400257 244454
rect 400191 244389 400257 244390
rect 400386 244159 400446 267921
rect 400575 266654 400641 266655
rect 400575 266590 400576 266654
rect 400640 266652 400641 266654
rect 400640 266592 401022 266652
rect 400640 266590 400641 266592
rect 400575 266589 400641 266590
rect 400767 264989 400833 264990
rect 400767 264925 400768 264989
rect 400832 264925 400833 264989
rect 400767 264924 400833 264925
rect 400770 245451 400830 264924
rect 400578 245391 400830 245451
rect 400578 244307 400638 245391
rect 400767 244750 400833 244751
rect 400767 244686 400768 244750
rect 400832 244748 400833 244750
rect 400962 244748 401022 266592
rect 401154 244751 401214 268365
rect 401343 266654 401409 266655
rect 401343 266590 401344 266654
rect 401408 266590 401409 266654
rect 401343 266589 401409 266590
rect 401535 266654 401601 266655
rect 401535 266590 401536 266654
rect 401600 266590 401601 266654
rect 401535 266589 401601 266590
rect 403263 266654 403329 266655
rect 403263 266590 403264 266654
rect 403328 266590 403329 266654
rect 403263 266589 403329 266590
rect 401346 247119 401406 266589
rect 401538 247449 401598 266589
rect 401538 247389 401982 247449
rect 401343 247118 401409 247119
rect 401343 247054 401344 247118
rect 401408 247054 401409 247118
rect 401343 247053 401409 247054
rect 401535 247118 401601 247119
rect 401535 247054 401536 247118
rect 401600 247054 401601 247118
rect 401535 247053 401601 247054
rect 401343 245046 401409 245047
rect 401343 244982 401344 245046
rect 401408 245044 401409 245046
rect 401538 245044 401598 247053
rect 401922 245047 401982 247389
rect 401408 244984 401598 245044
rect 401919 245046 401985 245047
rect 401408 244982 401409 244984
rect 401343 244981 401409 244982
rect 401919 244982 401920 245046
rect 401984 244982 401985 245046
rect 401919 244981 401985 244982
rect 400832 244688 401022 244748
rect 401151 244750 401217 244751
rect 400832 244686 400833 244688
rect 400767 244685 400833 244686
rect 401151 244686 401152 244750
rect 401216 244686 401217 244750
rect 401151 244685 401217 244686
rect 400575 244306 400641 244307
rect 400575 244242 400576 244306
rect 400640 244242 400641 244306
rect 400575 244241 400641 244242
rect 400383 244158 400449 244159
rect 400383 244094 400384 244158
rect 400448 244094 400449 244158
rect 400383 244093 400449 244094
rect 403266 244011 403326 266589
rect 403842 244603 403902 271621
rect 404031 270798 404097 270799
rect 404031 270734 404032 270798
rect 404096 270734 404097 270798
rect 404031 270733 404097 270734
rect 404034 244751 404094 270733
rect 404226 245047 404286 271769
rect 404418 267369 405246 267429
rect 404418 246971 404478 267369
rect 405186 266655 405246 267369
rect 404607 266654 404673 266655
rect 404607 266590 404608 266654
rect 404672 266590 404673 266654
rect 404607 266589 404673 266590
rect 404799 266654 404865 266655
rect 404799 266590 404800 266654
rect 404864 266590 404865 266654
rect 404799 266589 404865 266590
rect 405183 266654 405249 266655
rect 405183 266590 405184 266654
rect 405248 266590 405249 266654
rect 405183 266589 405249 266590
rect 404415 246970 404481 246971
rect 404415 246906 404416 246970
rect 404480 246906 404481 246970
rect 404415 246905 404481 246906
rect 404223 245046 404289 245047
rect 404223 244982 404224 245046
rect 404288 244982 404289 245046
rect 404223 244981 404289 244982
rect 404610 244751 404670 266589
rect 404802 247563 404862 266589
rect 405378 248781 405438 272361
rect 673983 270946 674049 270947
rect 673983 270882 673984 270946
rect 674048 270882 674049 270946
rect 673983 270881 674049 270882
rect 406143 266654 406209 266655
rect 406143 266590 406144 266654
rect 406208 266590 406209 266654
rect 406143 266589 406209 266590
rect 406527 266654 406593 266655
rect 406527 266590 406528 266654
rect 406592 266590 406593 266654
rect 406527 266589 406593 266590
rect 406911 266654 406977 266655
rect 406911 266590 406912 266654
rect 406976 266590 406977 266654
rect 406911 266589 406977 266590
rect 407103 266654 407169 266655
rect 407103 266590 407104 266654
rect 407168 266590 407169 266654
rect 407103 266589 407169 266590
rect 409023 266654 409089 266655
rect 409023 266590 409024 266654
rect 409088 266590 409089 266654
rect 409023 266589 409089 266590
rect 409407 266654 409473 266655
rect 409407 266590 409408 266654
rect 409472 266590 409473 266654
rect 409407 266589 409473 266590
rect 404994 248721 405438 248781
rect 404799 247562 404865 247563
rect 404799 247498 404800 247562
rect 404864 247498 404865 247562
rect 404799 247497 404865 247498
rect 404994 245047 405054 248721
rect 406146 247119 406206 266589
rect 406530 248115 406590 266589
rect 406338 248055 406590 248115
rect 406338 247415 406398 248055
rect 406335 247414 406401 247415
rect 406335 247350 406336 247414
rect 406400 247350 406401 247414
rect 406335 247349 406401 247350
rect 406143 247118 406209 247119
rect 406143 247054 406144 247118
rect 406208 247054 406209 247118
rect 406143 247053 406209 247054
rect 406914 245047 406974 266589
rect 407106 247267 407166 266589
rect 407103 247266 407169 247267
rect 407103 247202 407104 247266
rect 407168 247202 407169 247266
rect 407103 247201 407169 247202
rect 409026 245047 409086 266589
rect 409410 245047 409470 266589
rect 404991 245046 405057 245047
rect 404991 244982 404992 245046
rect 405056 244982 405057 245046
rect 404991 244981 405057 244982
rect 406911 245046 406977 245047
rect 406911 244982 406912 245046
rect 406976 244982 406977 245046
rect 406911 244981 406977 244982
rect 409023 245046 409089 245047
rect 409023 244982 409024 245046
rect 409088 244982 409089 245046
rect 409023 244981 409089 244982
rect 409407 245046 409473 245047
rect 409407 244982 409408 245046
rect 409472 244982 409473 245046
rect 409407 244981 409473 244982
rect 404031 244750 404097 244751
rect 404031 244686 404032 244750
rect 404096 244686 404097 244750
rect 404031 244685 404097 244686
rect 404607 244750 404673 244751
rect 404607 244686 404608 244750
rect 404672 244686 404673 244750
rect 404607 244685 404673 244686
rect 403839 244602 403905 244603
rect 403839 244538 403840 244602
rect 403904 244538 403905 244602
rect 403839 244537 403905 244538
rect 388863 244010 388929 244011
rect 388863 243946 388864 244010
rect 388928 243946 388929 244010
rect 388863 243945 388929 243946
rect 403263 244010 403329 244011
rect 403263 243946 403264 244010
rect 403328 243946 403329 244010
rect 403263 243945 403329 243946
rect 328575 243566 328641 243567
rect 328575 243502 328576 243566
rect 328640 243502 328641 243566
rect 328575 243501 328641 243502
rect 383103 241790 383169 241791
rect 383103 241726 383104 241790
rect 383168 241726 383169 241790
rect 383103 241725 383169 241726
rect 383106 239127 383166 241725
rect 383103 239126 383169 239127
rect 383103 239062 383104 239126
rect 383168 239062 383169 239126
rect 383103 239061 383169 239062
rect 212991 237646 213057 237647
rect 212991 237582 212992 237646
rect 213056 237582 213057 237646
rect 212991 237581 213057 237582
rect 212994 236611 213054 237581
rect 212991 236610 213057 236611
rect 212991 236546 212992 236610
rect 213056 236546 213057 236610
rect 212991 236545 213057 236546
rect 210303 236314 210369 236315
rect 210303 236250 210304 236314
rect 210368 236250 210369 236314
rect 210303 236249 210369 236250
rect 211455 234686 211521 234687
rect 211455 234622 211456 234686
rect 211520 234622 211521 234686
rect 211455 234621 211521 234622
rect 211071 233650 211137 233651
rect 211071 233586 211072 233650
rect 211136 233586 211137 233650
rect 211071 233585 211137 233586
rect 210879 233354 210945 233355
rect 210879 233290 210880 233354
rect 210944 233290 210945 233354
rect 210879 233289 210945 233290
rect 210303 232910 210369 232911
rect 210303 232846 210304 232910
rect 210368 232846 210369 232910
rect 210303 232845 210369 232846
rect 145599 221810 145665 221811
rect 145599 221746 145600 221810
rect 145664 221746 145665 221810
rect 145599 221745 145665 221746
rect 145407 51462 145473 51463
rect 145407 51398 145408 51462
rect 145472 51398 145473 51462
rect 145407 51397 145473 51398
rect 145602 51315 145662 221745
rect 207231 210266 207297 210267
rect 207231 210202 207232 210266
rect 207296 210202 207297 210266
rect 207231 210201 207297 210202
rect 207234 190139 207294 210201
rect 210306 200647 210366 232845
rect 210495 223142 210561 223143
rect 210495 223078 210496 223142
rect 210560 223078 210561 223142
rect 210495 223077 210561 223078
rect 210303 200646 210369 200647
rect 210303 200582 210304 200646
rect 210368 200582 210369 200646
rect 210303 200581 210369 200582
rect 210498 199019 210558 223077
rect 210882 200163 210942 233289
rect 211074 223143 211134 233585
rect 211071 223142 211137 223143
rect 211071 223078 211072 223142
rect 211136 223078 211137 223142
rect 211071 223077 211137 223078
rect 211458 218811 211518 234621
rect 212031 233798 212097 233799
rect 212031 233734 212032 233798
rect 212096 233734 212097 233798
rect 212031 233733 212097 233734
rect 211647 233650 211713 233651
rect 211647 233586 211648 233650
rect 211712 233586 211713 233650
rect 211647 233585 211713 233586
rect 211650 222141 211710 233585
rect 211650 222081 211758 222141
rect 211698 221475 211758 222081
rect 211266 218751 211518 218811
rect 211650 221415 211758 221475
rect 211266 207489 211326 218751
rect 211650 208821 211710 221415
rect 211650 208761 211902 208821
rect 211266 207429 211710 207489
rect 211071 200646 211137 200647
rect 211071 200582 211072 200646
rect 211136 200582 211137 200646
rect 211071 200581 211137 200582
rect 210690 200103 210942 200163
rect 211074 200163 211134 200581
rect 211074 200103 211326 200163
rect 210495 199018 210561 199019
rect 210495 198954 210496 199018
rect 210560 198954 210561 199018
rect 210495 198953 210561 198954
rect 210690 198831 210750 200103
rect 211071 198870 211137 198871
rect 210690 198771 210942 198831
rect 211071 198806 211072 198870
rect 211136 198806 211137 198870
rect 211071 198805 211137 198806
rect 207231 190138 207297 190139
rect 207231 190074 207232 190138
rect 207296 190074 207297 190138
rect 207231 190073 207297 190074
rect 210882 172675 210942 198771
rect 211074 172823 211134 198805
rect 211071 172822 211137 172823
rect 211071 172758 211072 172822
rect 211136 172758 211137 172822
rect 211071 172757 211137 172758
rect 210879 172674 210945 172675
rect 210879 172610 210880 172674
rect 210944 172610 210945 172674
rect 210879 172609 210945 172610
rect 210303 172526 210369 172527
rect 210303 172462 210304 172526
rect 210368 172462 210369 172526
rect 211266 172524 211326 200103
rect 211650 177519 211710 207429
rect 210303 172461 210369 172462
rect 210690 172464 211326 172524
rect 211458 177459 211710 177519
rect 210306 162867 210366 172461
rect 210306 162807 210558 162867
rect 210303 151658 210369 151659
rect 210303 151594 210304 151658
rect 210368 151594 210369 151658
rect 210303 151593 210369 151594
rect 146751 134490 146817 134491
rect 146751 134426 146752 134490
rect 146816 134426 146817 134490
rect 146751 134425 146817 134426
rect 146754 132567 146814 134425
rect 146751 132566 146817 132567
rect 146751 132502 146752 132566
rect 146816 132502 146817 132566
rect 146751 132501 146817 132502
rect 146559 126794 146625 126795
rect 146559 126730 146560 126794
rect 146624 126730 146625 126794
rect 146559 126729 146625 126730
rect 146562 115251 146622 126729
rect 209727 123834 209793 123835
rect 209727 123770 209728 123834
rect 209792 123770 209793 123834
rect 209727 123769 209793 123770
rect 146559 115250 146625 115251
rect 146559 115186 146560 115250
rect 146624 115186 146625 115250
rect 146559 115185 146625 115186
rect 209730 77807 209790 123769
rect 210306 122503 210366 151593
rect 210498 132715 210558 162807
rect 210690 152843 210750 172464
rect 211458 163533 211518 177459
rect 211842 169527 211902 208761
rect 211650 169467 211902 169527
rect 211650 164199 211710 169467
rect 212034 168861 212094 233733
rect 212994 233651 213054 236545
rect 637311 233798 637377 233799
rect 637311 233734 637312 233798
rect 637376 233734 637377 233798
rect 637311 233733 637377 233734
rect 212223 233650 212289 233651
rect 212223 233586 212224 233650
rect 212288 233586 212289 233650
rect 212223 233585 212289 233586
rect 212415 233650 212481 233651
rect 212415 233586 212416 233650
rect 212480 233586 212481 233650
rect 212415 233585 212481 233586
rect 212991 233650 213057 233651
rect 212991 233586 212992 233650
rect 213056 233586 213057 233650
rect 212991 233585 213057 233586
rect 636927 233650 636993 233651
rect 636927 233586 636928 233650
rect 636992 233586 636993 233650
rect 636927 233585 636993 233586
rect 212226 169527 212286 233585
rect 212418 232911 212478 233585
rect 212991 233502 213057 233503
rect 212991 233438 212992 233502
rect 213056 233438 213057 233502
rect 212991 233437 213057 233438
rect 212415 232910 212481 232911
rect 212415 232846 212416 232910
rect 212480 232846 212481 232910
rect 212415 232845 212481 232846
rect 212994 196167 213054 233437
rect 212418 196107 213054 196167
rect 212418 185511 212478 196107
rect 212418 185451 213054 185511
rect 212226 169467 212670 169527
rect 212034 168801 212478 168861
rect 211650 164139 211902 164199
rect 210882 163473 211518 163533
rect 210687 152842 210753 152843
rect 210687 152778 210688 152842
rect 210752 152778 210753 152842
rect 210687 152777 210753 152778
rect 210687 152694 210753 152695
rect 210687 152630 210688 152694
rect 210752 152630 210753 152694
rect 210687 152629 210753 152630
rect 210690 142036 210750 152629
rect 210882 142887 210942 163473
rect 211071 152694 211137 152695
rect 211071 152630 211072 152694
rect 211136 152692 211137 152694
rect 211136 152632 211710 152692
rect 211136 152630 211137 152632
rect 211071 152629 211137 152630
rect 211071 151658 211137 151659
rect 211071 151594 211072 151658
rect 211136 151656 211137 151658
rect 211650 151656 211710 152632
rect 211136 151596 211710 151656
rect 211136 151594 211137 151596
rect 211071 151593 211137 151594
rect 211842 149547 211902 164139
rect 212418 162867 212478 168801
rect 211650 149487 211902 149547
rect 212034 162807 212478 162867
rect 211650 143553 211710 149487
rect 211650 143493 211902 143553
rect 210882 142827 211134 142887
rect 210690 141976 210942 142036
rect 210495 132714 210561 132715
rect 210495 132650 210496 132714
rect 210560 132650 210561 132714
rect 210495 132649 210561 132650
rect 210495 123982 210561 123983
rect 210495 123918 210496 123982
rect 210560 123918 210561 123982
rect 210495 123917 210561 123918
rect 210303 122502 210369 122503
rect 210303 122438 210304 122502
rect 210368 122438 210369 122502
rect 210303 122437 210369 122438
rect 209919 118506 209985 118507
rect 209919 118442 209920 118506
rect 209984 118442 209985 118506
rect 209919 118441 209985 118442
rect 209922 82247 209982 118441
rect 210111 106814 210177 106815
rect 210111 106750 210112 106814
rect 210176 106750 210177 106814
rect 210111 106749 210177 106750
rect 210114 93199 210174 106749
rect 210303 95862 210369 95863
rect 210303 95798 210304 95862
rect 210368 95798 210369 95862
rect 210303 95797 210369 95798
rect 210111 93198 210177 93199
rect 210111 93134 210112 93198
rect 210176 93134 210177 93198
rect 210111 93133 210177 93134
rect 210306 93051 210366 95797
rect 210303 93050 210369 93051
rect 210303 92986 210304 93050
rect 210368 92986 210369 93050
rect 210303 92985 210369 92986
rect 209919 82246 209985 82247
rect 209919 82182 209920 82246
rect 209984 82182 209985 82246
rect 209919 82181 209985 82182
rect 210498 81211 210558 123917
rect 210882 123835 210942 141976
rect 211074 133563 211134 142827
rect 211074 133503 211710 133563
rect 211071 132714 211137 132715
rect 211071 132650 211072 132714
rect 211136 132650 211137 132714
rect 211071 132649 211137 132650
rect 211074 123983 211134 132649
rect 211071 123982 211137 123983
rect 211071 123918 211072 123982
rect 211136 123918 211137 123982
rect 211071 123917 211137 123918
rect 210879 123834 210945 123835
rect 210879 123770 210880 123834
rect 210944 123770 210945 123834
rect 210879 123769 210945 123770
rect 211650 123573 211710 133503
rect 211074 123513 211710 123573
rect 210879 122502 210945 122503
rect 210879 122438 210880 122502
rect 210944 122438 210945 122502
rect 210879 122437 210945 122438
rect 210882 106815 210942 122437
rect 211074 119099 211134 123513
rect 211842 123240 211902 143493
rect 212034 123832 212094 162807
rect 212610 162201 212670 169467
rect 212226 162141 212670 162201
rect 212226 148881 212286 162141
rect 212226 148821 212478 148881
rect 212418 124239 212478 148821
rect 212994 142887 213054 185451
rect 212802 142827 213054 142887
rect 212418 124179 212670 124239
rect 212034 123772 212478 123832
rect 211650 123180 211902 123240
rect 211071 119098 211137 119099
rect 211071 119034 211072 119098
rect 211136 119034 211137 119098
rect 211071 119033 211137 119034
rect 211650 118911 211710 123180
rect 211074 118851 211710 118911
rect 211074 118507 211134 118851
rect 211071 118506 211137 118507
rect 211071 118442 211072 118506
rect 211136 118442 211137 118506
rect 211071 118441 211137 118442
rect 212418 118245 212478 123772
rect 211074 118185 212478 118245
rect 210879 106814 210945 106815
rect 210879 106750 210880 106814
rect 210944 106750 210945 106814
rect 210879 106749 210945 106750
rect 211074 106257 211134 118185
rect 212610 117579 212670 124179
rect 210690 106197 211134 106257
rect 212226 117519 212670 117579
rect 210690 99597 210750 106197
rect 210690 99537 212094 99597
rect 212034 97599 212094 99537
rect 210882 97539 212094 97599
rect 210687 96898 210753 96899
rect 210687 96834 210688 96898
rect 210752 96834 210753 96898
rect 210687 96833 210753 96834
rect 210495 81210 210561 81211
rect 210495 81146 210496 81210
rect 210560 81146 210561 81210
rect 210495 81145 210561 81146
rect 209727 77806 209793 77807
rect 209727 77742 209728 77806
rect 209792 77742 209793 77806
rect 209727 77741 209793 77742
rect 210690 53831 210750 96833
rect 210882 82947 210942 97539
rect 212226 96933 212286 117519
rect 212802 116913 212862 142827
rect 211074 96899 212286 96933
rect 211071 96898 212286 96899
rect 211071 96834 211072 96898
rect 211136 96873 212286 96898
rect 212418 116853 212862 116913
rect 211136 96834 211137 96873
rect 211071 96833 211137 96834
rect 212418 96267 212478 116853
rect 211074 96207 212478 96267
rect 211074 95863 211134 96207
rect 211071 95862 211137 95863
rect 211071 95798 211072 95862
rect 211136 95798 211137 95862
rect 211071 95797 211137 95798
rect 211071 94234 211137 94235
rect 211071 94170 211072 94234
rect 211136 94232 211137 94234
rect 211136 94172 211902 94232
rect 211136 94170 211137 94172
rect 211071 94169 211137 94170
rect 211071 93198 211137 93199
rect 211071 93134 211072 93198
rect 211136 93196 211137 93198
rect 211136 93136 211326 93196
rect 211136 93134 211137 93136
rect 211071 93133 211137 93134
rect 211071 93050 211137 93051
rect 211071 92986 211072 93050
rect 211136 92986 211137 93050
rect 211071 92985 211137 92986
rect 211074 90273 211134 92985
rect 211266 91605 211326 93136
rect 211842 92271 211902 94172
rect 211842 92211 213054 92271
rect 211266 91545 212862 91605
rect 211074 90213 211518 90273
rect 211458 84279 211518 90213
rect 211458 84219 212286 84279
rect 212226 83613 212286 84219
rect 212226 83553 212478 83613
rect 210882 82887 211134 82947
rect 211074 82281 211134 82887
rect 210879 82246 210945 82247
rect 210879 82182 210880 82246
rect 210944 82182 210945 82246
rect 211074 82221 212286 82281
rect 210879 82181 210945 82182
rect 210882 81615 210942 82181
rect 210882 81555 211326 81615
rect 211071 81210 211137 81211
rect 211071 81146 211072 81210
rect 211136 81146 211137 81210
rect 211071 81145 211137 81146
rect 210879 77806 210945 77807
rect 210879 77742 210880 77806
rect 210944 77742 210945 77806
rect 210879 77741 210945 77742
rect 210882 54275 210942 77741
rect 211074 59637 211134 81145
rect 211266 68961 211326 81555
rect 211266 68901 211710 68961
rect 211074 59577 211326 59637
rect 211071 58270 211137 58271
rect 211071 58206 211072 58270
rect 211136 58206 211137 58270
rect 211071 58205 211137 58206
rect 210879 54274 210945 54275
rect 210879 54210 210880 54274
rect 210944 54210 210945 54274
rect 210879 54209 210945 54210
rect 210687 53830 210753 53831
rect 210687 53766 210688 53830
rect 210752 53766 210753 53830
rect 210687 53765 210753 53766
rect 211074 53091 211134 58205
rect 211266 54127 211326 59577
rect 211650 57639 211710 68901
rect 211650 57579 211902 57639
rect 211263 54126 211329 54127
rect 211263 54062 211264 54126
rect 211328 54062 211329 54126
rect 211263 54061 211329 54062
rect 211842 53683 211902 57579
rect 212226 53979 212286 82221
rect 212223 53978 212289 53979
rect 212223 53914 212224 53978
rect 212288 53914 212289 53978
rect 212223 53913 212289 53914
rect 211839 53682 211905 53683
rect 211839 53618 211840 53682
rect 211904 53618 211905 53682
rect 211839 53617 211905 53618
rect 212418 53387 212478 83553
rect 212802 60303 212862 91545
rect 212610 60243 212862 60303
rect 212610 54275 212670 60243
rect 212994 56307 213054 92211
rect 212994 56247 213102 56307
rect 213042 54975 213102 56247
rect 212994 54915 213102 54975
rect 212607 54274 212673 54275
rect 212607 54210 212608 54274
rect 212672 54210 212673 54274
rect 212607 54209 212673 54210
rect 212994 53535 213054 54915
rect 212991 53534 213057 53535
rect 212991 53470 212992 53534
rect 213056 53470 213057 53534
rect 212991 53469 213057 53470
rect 212415 53386 212481 53387
rect 212415 53322 212416 53386
rect 212480 53322 212481 53386
rect 212415 53321 212481 53322
rect 211071 53090 211137 53091
rect 211071 53026 211072 53090
rect 211136 53026 211137 53090
rect 211071 53025 211137 53026
rect 145599 51314 145665 51315
rect 145599 51250 145600 51314
rect 145664 51250 145665 51314
rect 145599 51249 145665 51250
rect 636930 50427 636990 233585
rect 637119 233502 637185 233503
rect 637119 233438 637120 233502
rect 637184 233438 637185 233502
rect 637119 233437 637185 233438
rect 637122 51611 637182 233437
rect 637314 51759 637374 233733
rect 637503 233650 637569 233651
rect 637503 233586 637504 233650
rect 637568 233586 637569 233650
rect 637503 233585 637569 233586
rect 637506 52055 637566 233585
rect 637887 233502 637953 233503
rect 637887 233438 637888 233502
rect 637952 233438 637953 233502
rect 637887 233437 637953 233438
rect 637695 233354 637761 233355
rect 637695 233290 637696 233354
rect 637760 233290 637761 233354
rect 637695 233289 637761 233290
rect 637503 52054 637569 52055
rect 637503 51990 637504 52054
rect 637568 51990 637569 52054
rect 637503 51989 637569 51990
rect 637698 51907 637758 233289
rect 637890 52203 637950 233437
rect 673986 227435 674046 270881
rect 674178 270207 674238 315725
rect 674559 314310 674625 314311
rect 674559 314246 674560 314310
rect 674624 314246 674625 314310
rect 674559 314245 674625 314246
rect 674367 313274 674433 313275
rect 674367 313210 674368 313274
rect 674432 313210 674433 313274
rect 674367 313209 674433 313210
rect 674370 283675 674430 313209
rect 674367 283674 674433 283675
rect 674367 283610 674368 283674
rect 674432 283610 674433 283674
rect 674367 283609 674433 283610
rect 674175 270206 674241 270207
rect 674175 270142 674176 270206
rect 674240 270142 674241 270206
rect 674175 270141 674241 270142
rect 674178 244751 674238 270141
rect 674562 269763 674622 314245
rect 674751 285006 674817 285007
rect 674751 284942 674752 285006
rect 674816 284942 674817 285006
rect 674751 284941 674817 284942
rect 674559 269762 674625 269763
rect 674559 269698 674560 269762
rect 674624 269698 674625 269762
rect 674559 269697 674625 269698
rect 674559 265470 674625 265471
rect 674559 265406 674560 265470
rect 674624 265406 674625 265470
rect 674559 265405 674625 265406
rect 674175 244750 674241 244751
rect 674175 244686 674176 244750
rect 674240 244686 674241 244750
rect 674175 244685 674241 244686
rect 674562 243567 674622 265405
rect 674754 246823 674814 284941
rect 674946 272871 675006 315873
rect 675330 289595 675390 333781
rect 676290 333551 676350 345325
rect 676287 333550 676353 333551
rect 676287 333486 676288 333550
rect 676352 333486 676353 333550
rect 676287 333485 676353 333486
rect 675519 329554 675585 329555
rect 675519 329490 675520 329554
rect 675584 329490 675585 329554
rect 675519 329489 675585 329490
rect 675522 289743 675582 329489
rect 676482 328075 676542 345473
rect 676671 345242 676737 345243
rect 676671 345178 676672 345242
rect 676736 345178 676737 345242
rect 676671 345177 676737 345178
rect 676479 328074 676545 328075
rect 676479 328010 676480 328074
rect 676544 328010 676545 328074
rect 676479 328009 676545 328010
rect 676674 326891 676734 345177
rect 676671 326890 676737 326891
rect 676671 326826 676672 326890
rect 676736 326826 676737 326890
rect 676671 326825 676737 326826
rect 675903 299510 675969 299511
rect 675903 299446 675904 299510
rect 675968 299446 675969 299510
rect 675903 299445 675969 299446
rect 675519 289742 675585 289743
rect 675519 289678 675520 289742
rect 675584 289678 675585 289742
rect 675519 289677 675585 289678
rect 675327 289594 675393 289595
rect 675327 289530 675328 289594
rect 675392 289530 675393 289594
rect 675327 289529 675393 289530
rect 674943 272870 675009 272871
rect 674943 272806 674944 272870
rect 675008 272806 675009 272870
rect 674943 272805 675009 272806
rect 675135 269762 675201 269763
rect 675135 269698 675136 269762
rect 675200 269698 675201 269762
rect 675135 269697 675201 269698
rect 674943 267986 675009 267987
rect 674943 267922 674944 267986
rect 675008 267922 675009 267986
rect 674943 267921 675009 267922
rect 674751 246822 674817 246823
rect 674751 246758 674752 246822
rect 674816 246758 674817 246822
rect 674751 246757 674817 246758
rect 674754 245935 674814 246757
rect 674751 245934 674817 245935
rect 674751 245870 674752 245934
rect 674816 245870 674817 245934
rect 674751 245869 674817 245870
rect 674559 243566 674625 243567
rect 674559 243502 674560 243566
rect 674624 243502 674625 243566
rect 674559 243501 674625 243502
rect 674946 238683 675006 267921
rect 675138 244603 675198 269697
rect 675522 245195 675582 289677
rect 675906 284859 675966 299445
rect 676671 299362 676737 299363
rect 676671 299298 676672 299362
rect 676736 299298 676737 299362
rect 676671 299297 676737 299298
rect 675903 284858 675969 284859
rect 675903 284794 675904 284858
rect 675968 284794 675969 284858
rect 675903 284793 675969 284794
rect 676674 281899 676734 299297
rect 676671 281898 676737 281899
rect 676671 281834 676672 281898
rect 676736 281834 676737 281898
rect 676671 281833 676737 281834
rect 675711 253482 675777 253483
rect 675711 253418 675712 253482
rect 675776 253418 675777 253482
rect 675711 253417 675777 253418
rect 675519 245194 675585 245195
rect 675519 245130 675520 245194
rect 675584 245130 675585 245194
rect 675519 245129 675585 245130
rect 675135 244602 675201 244603
rect 675135 244538 675136 244602
rect 675200 244538 675201 244602
rect 675135 244537 675201 244538
rect 675327 241938 675393 241939
rect 675327 241874 675328 241938
rect 675392 241874 675393 241938
rect 675327 241873 675393 241874
rect 674943 238682 675009 238683
rect 674943 238618 674944 238682
rect 675008 238618 675009 238682
rect 674943 238617 675009 238618
rect 673983 227434 674049 227435
rect 673983 227370 673984 227434
rect 674048 227370 674049 227434
rect 673983 227369 674049 227370
rect 673983 226250 674049 226251
rect 673983 226186 673984 226250
rect 674048 226186 674049 226250
rect 673983 226185 674049 226186
rect 673986 182591 674046 226185
rect 674367 223142 674433 223143
rect 674367 223078 674368 223142
rect 674432 223078 674433 223142
rect 674367 223077 674433 223078
rect 674370 193543 674430 223077
rect 675330 199315 675390 241873
rect 675519 238978 675585 238979
rect 675519 238914 675520 238978
rect 675584 238914 675585 238978
rect 675519 238913 675585 238914
rect 675327 199314 675393 199315
rect 675327 199250 675328 199314
rect 675392 199250 675393 199314
rect 675327 199249 675393 199250
rect 674367 193542 674433 193543
rect 674367 193478 674368 193542
rect 674432 193478 674433 193542
rect 674367 193477 674433 193478
rect 673983 182590 674049 182591
rect 673983 182526 673984 182590
rect 674048 182526 674049 182590
rect 673983 182525 674049 182526
rect 673983 181258 674049 181259
rect 673983 181194 673984 181258
rect 674048 181194 674049 181258
rect 673983 181193 674049 181194
rect 673986 136859 674046 181193
rect 674751 178594 674817 178595
rect 674751 178530 674752 178594
rect 674816 178530 674817 178594
rect 674751 178529 674817 178530
rect 674175 178150 674241 178151
rect 674175 178086 674176 178150
rect 674240 178086 674241 178150
rect 674175 178085 674241 178086
rect 674178 148551 674238 178085
rect 674559 166458 674625 166459
rect 674559 166394 674560 166458
rect 674624 166394 674625 166458
rect 674559 166393 674625 166394
rect 674367 165570 674433 165571
rect 674367 165506 674368 165570
rect 674432 165506 674433 165570
rect 674367 165505 674433 165506
rect 674175 148550 674241 148551
rect 674175 148486 674176 148550
rect 674240 148486 674241 148550
rect 674175 148485 674241 148486
rect 673983 136858 674049 136859
rect 673983 136794 673984 136858
rect 674048 136794 674049 136858
rect 673983 136793 674049 136794
rect 674370 134565 674430 165505
rect 674562 135527 674622 166393
rect 674754 159355 674814 178529
rect 674751 159354 674817 159355
rect 674751 159290 674752 159354
rect 674816 159290 674817 159354
rect 674751 159289 674817 159290
rect 675330 154619 675390 199249
rect 675522 198723 675582 238913
rect 675714 236907 675774 253417
rect 675711 236906 675777 236907
rect 675711 236842 675712 236906
rect 675776 236842 675777 236906
rect 675711 236841 675777 236842
rect 676479 210266 676545 210267
rect 676479 210202 676480 210266
rect 676544 210202 676545 210266
rect 676479 210201 676545 210202
rect 675903 207750 675969 207751
rect 675903 207686 675904 207750
rect 675968 207686 675969 207750
rect 675903 207685 675969 207686
rect 675519 198722 675585 198723
rect 675519 198658 675520 198722
rect 675584 198658 675585 198722
rect 675519 198657 675585 198658
rect 675327 154618 675393 154619
rect 675327 154554 675328 154618
rect 675392 154554 675393 154618
rect 675327 154553 675393 154554
rect 674751 148402 674817 148403
rect 674751 148338 674752 148402
rect 674816 148338 674817 148402
rect 674751 148337 674817 148338
rect 674559 135526 674625 135527
rect 674559 135462 674560 135526
rect 674624 135462 674625 135526
rect 674559 135461 674625 135462
rect 674559 134934 674625 134935
rect 674559 134870 674560 134934
rect 674624 134895 674625 134934
rect 674754 134895 674814 148337
rect 674624 134870 674814 134895
rect 674559 134869 674814 134870
rect 674562 134835 674814 134869
rect 674367 134564 674433 134565
rect 674367 134500 674368 134564
rect 674432 134500 674433 134564
rect 674367 134499 674433 134500
rect 674175 133750 674241 133751
rect 674175 133686 674176 133750
rect 674240 133686 674241 133750
rect 674175 133685 674241 133686
rect 674178 114215 674238 133685
rect 674175 114214 674241 114215
rect 674175 114150 674176 114214
rect 674240 114150 674241 114214
rect 674175 114149 674241 114150
rect 674754 109331 674814 134835
rect 674943 132566 675009 132567
rect 674943 132502 674944 132566
rect 675008 132502 675009 132566
rect 674943 132501 675009 132502
rect 674751 109330 674817 109331
rect 674751 109266 674752 109330
rect 674816 109266 674817 109330
rect 674751 109265 674817 109266
rect 674946 103263 675006 132501
rect 675330 110071 675390 154553
rect 675522 154323 675582 198657
rect 675906 198427 675966 207685
rect 676287 207602 676353 207603
rect 676287 207538 676288 207602
rect 676352 207538 676353 207602
rect 676287 207537 676353 207538
rect 676095 207454 676161 207455
rect 676095 207390 676096 207454
rect 676160 207390 676161 207454
rect 676095 207389 676161 207390
rect 675903 198426 675969 198427
rect 675903 198362 675904 198426
rect 675968 198362 675969 198426
rect 675903 198361 675969 198362
rect 676098 195319 676158 207389
rect 676095 195318 676161 195319
rect 676095 195254 676096 195318
rect 676160 195254 676161 195318
rect 676095 195253 676161 195254
rect 676290 191619 676350 207537
rect 676287 191618 676353 191619
rect 676287 191554 676288 191618
rect 676352 191554 676353 191618
rect 676287 191553 676353 191554
rect 676482 180963 676542 210201
rect 676671 210118 676737 210119
rect 676671 210054 676672 210118
rect 676736 210054 676737 210118
rect 676671 210053 676737 210054
rect 676479 180962 676545 180963
rect 676479 180898 676480 180962
rect 676544 180898 676545 180962
rect 676479 180897 676545 180898
rect 676674 179483 676734 210053
rect 676671 179482 676737 179483
rect 676671 179418 676672 179482
rect 676736 179418 676737 179482
rect 676671 179417 676737 179418
rect 676671 164090 676737 164091
rect 676671 164026 676672 164090
rect 676736 164026 676737 164090
rect 676671 164025 676737 164026
rect 676479 162906 676545 162907
rect 676479 162842 676480 162906
rect 676544 162842 676545 162906
rect 676479 162841 676545 162842
rect 675903 161426 675969 161427
rect 675903 161362 675904 161426
rect 675968 161362 675969 161426
rect 675903 161361 675969 161362
rect 675906 157727 675966 161361
rect 675903 157726 675969 157727
rect 675903 157662 675904 157726
rect 675968 157662 675969 157726
rect 675903 157661 675969 157662
rect 675519 154322 675585 154323
rect 675519 154258 675520 154322
rect 675584 154258 675585 154322
rect 675519 154257 675585 154258
rect 676482 153435 676542 162841
rect 676479 153434 676545 153435
rect 676479 153370 676480 153434
rect 676544 153370 676545 153434
rect 676479 153369 676545 153370
rect 676674 146627 676734 164025
rect 676671 146626 676737 146627
rect 676671 146562 676672 146626
rect 676736 146562 676737 146626
rect 676671 146561 676737 146562
rect 675903 120430 675969 120431
rect 675903 120366 675904 120430
rect 675968 120366 675969 120430
rect 675903 120365 675969 120366
rect 675327 110070 675393 110071
rect 675327 110006 675328 110070
rect 675392 110006 675393 110070
rect 675327 110005 675393 110006
rect 675906 108147 675966 120365
rect 676671 118062 676737 118063
rect 676671 117998 676672 118062
rect 676736 117998 676737 118062
rect 676671 117997 676737 117998
rect 675903 108146 675969 108147
rect 675903 108082 675904 108146
rect 675968 108082 675969 108146
rect 675903 108081 675969 108082
rect 674943 103262 675009 103263
rect 674943 103198 674944 103262
rect 675008 103198 675009 103262
rect 674943 103197 675009 103198
rect 676674 101487 676734 117997
rect 676671 101486 676737 101487
rect 676671 101422 676672 101486
rect 676736 101422 676737 101486
rect 676671 101421 676737 101422
rect 637887 52202 637953 52203
rect 637887 52138 637888 52202
rect 637952 52138 637953 52202
rect 637887 52137 637953 52138
rect 637695 51906 637761 51907
rect 637695 51842 637696 51906
rect 637760 51842 637761 51906
rect 637695 51841 637761 51842
rect 637311 51758 637377 51759
rect 637311 51694 637312 51758
rect 637376 51694 637377 51758
rect 637311 51693 637377 51694
rect 637119 51610 637185 51611
rect 637119 51546 637120 51610
rect 637184 51546 637185 51610
rect 637119 51545 637185 51546
rect 636927 50426 636993 50427
rect 636927 50362 636928 50426
rect 636992 50362 636993 50426
rect 636927 50361 636993 50362
rect 471039 46134 471105 46135
rect 471039 46070 471040 46134
rect 471104 46070 471105 46134
rect 471039 46069 471105 46070
rect 302463 45098 302529 45099
rect 302463 45034 302464 45098
rect 302528 45034 302529 45098
rect 302463 45033 302529 45034
rect 302466 43323 302526 45033
rect 414783 44950 414849 44951
rect 414783 44886 414784 44950
rect 414848 44886 414849 44950
rect 414783 44885 414849 44886
rect 414786 43323 414846 44885
rect 302463 43322 302529 43323
rect 302463 43258 302464 43322
rect 302528 43258 302529 43322
rect 302463 43257 302529 43258
rect 414783 43322 414849 43323
rect 414783 43258 414784 43322
rect 414848 43258 414849 43322
rect 414783 43257 414849 43258
rect 471042 42139 471102 46069
rect 471039 42138 471105 42139
rect 471039 42074 471040 42138
rect 471104 42074 471105 42138
rect 471039 42073 471105 42074
rect 189951 41842 190017 41843
rect 189951 41778 189952 41842
rect 190016 41778 190017 41842
rect 189951 41777 190017 41778
rect 194943 41842 195009 41843
rect 194943 41778 194944 41842
rect 195008 41778 195009 41842
rect 194943 41777 195009 41778
rect 360063 41842 360129 41843
rect 360063 41778 360064 41842
rect 360128 41778 360129 41842
rect 360063 41777 360129 41778
rect 362943 41842 363009 41843
rect 362943 41778 362944 41842
rect 363008 41778 363009 41842
rect 362943 41777 363009 41778
rect 459327 41842 459393 41843
rect 459327 41778 459328 41842
rect 459392 41778 459393 41842
rect 459327 41777 459393 41778
rect 189954 40807 190014 41777
rect 189951 40806 190017 40807
rect 189951 40742 189952 40806
rect 190016 40742 190017 40806
rect 189951 40741 190017 40742
rect 194946 40659 195006 41777
rect 360066 40955 360126 41777
rect 360063 40954 360129 40955
rect 360063 40890 360064 40954
rect 360128 40890 360129 40954
rect 360063 40889 360129 40890
rect 362946 40807 363006 41777
rect 362943 40806 363009 40807
rect 362943 40742 362944 40806
rect 363008 40742 363009 40806
rect 362943 40741 363009 40742
rect 194943 40658 195009 40659
rect 194943 40594 194944 40658
rect 195008 40594 195009 40658
rect 194943 40593 195009 40594
rect 459330 40411 459390 41777
<< via4 >>
rect 324074 270611 324310 270847
rect 330986 270611 331222 270847
rect 322922 269945 323158 270181
rect 342506 269945 342742 270181
rect 368426 270611 368662 270847
rect 383978 270798 384214 270847
rect 383978 270734 384064 270798
rect 384064 270734 384128 270798
rect 384128 270734 384214 270798
rect 383978 270611 384214 270734
rect 370922 269945 371158 270181
rect 384554 269945 384790 270181
rect 377066 268613 377302 268849
rect 368426 267947 368662 268183
rect 378986 267947 379222 268183
rect 372842 267281 373078 267517
rect 356906 266615 357142 266851
rect 368426 266654 368662 266851
rect 368426 266615 368512 266654
rect 368512 266615 368576 266654
rect 368576 266615 368662 266654
rect 374378 266615 374614 266851
rect 389354 268613 389590 268849
rect 388202 267281 388438 267517
rect 387050 266615 387286 266851
rect 325418 265283 325654 265519
rect 328682 265283 328918 265519
rect 364970 265283 365206 265519
rect 378602 265283 378838 265519
rect 455018 40362 455254 40411
rect 455018 40298 455104 40362
rect 455104 40298 455168 40362
rect 455168 40298 455254 40362
rect 455018 40175 455254 40298
rect 459242 40175 459478 40411
<< metal5 >>
rect 324032 270847 331264 270889
rect 324032 270611 324074 270847
rect 324310 270611 330986 270847
rect 331222 270611 331264 270847
rect 324032 270569 331264 270611
rect 368384 270847 384256 270889
rect 368384 270611 368426 270847
rect 368662 270611 383978 270847
rect 384214 270611 384256 270847
rect 368384 270569 384256 270611
rect 322880 270181 342784 270223
rect 322880 269945 322922 270181
rect 323158 269945 342506 270181
rect 342742 269945 342784 270181
rect 322880 269903 342784 269945
rect 370880 270181 384832 270223
rect 370880 269945 370922 270181
rect 371158 269945 384554 270181
rect 384790 269945 384832 270181
rect 370880 269903 384832 269945
rect 377024 268849 389632 268891
rect 377024 268613 377066 268849
rect 377302 268613 389354 268849
rect 389590 268613 389632 268849
rect 377024 268571 389632 268613
rect 368384 268183 379264 268225
rect 368384 267947 368426 268183
rect 368662 267947 378986 268183
rect 379222 267947 379264 268183
rect 368384 267905 379264 267947
rect 372800 267517 388480 267559
rect 372800 267281 372842 267517
rect 373078 267281 388202 267517
rect 388438 267281 388480 267517
rect 372800 267239 388480 267281
rect 356864 266851 368704 266893
rect 356864 266615 356906 266851
rect 357142 266615 368426 266851
rect 368662 266615 368704 266851
rect 356864 266573 368704 266615
rect 374336 266851 387328 266893
rect 374336 266615 374378 266851
rect 374614 266615 387050 266851
rect 387286 266615 387328 266851
rect 374336 266573 387328 266615
rect 325376 265519 328960 265561
rect 325376 265283 325418 265519
rect 325654 265283 328682 265519
rect 328918 265283 328960 265519
rect 325376 265241 328960 265283
rect 364928 265519 378880 265561
rect 364928 265283 364970 265519
rect 365206 265283 378602 265519
rect 378838 265283 378880 265519
rect 364928 265241 378880 265283
rect 454976 40411 459520 40453
rect 454976 40175 455018 40411
rect 455254 40175 459242 40411
rect 459478 40175 459520 40411
rect 454976 40133 459520 40175
use user_id_programming  user_id_value ../mag
timestamp 1608153117
transform 1 0 656624 0 1 80926
box 0 0 7109 7077
use storage  storage ../mag
timestamp 1608153117
transform 1 0 52032 0 1 53156
box 0 0 88934 189234
use mgmt_core  soc ../mag
timestamp 1608153117
transform 1 0 210422 0 1 53602
box 0 0 430000 180000
use sky130_fd_sc_hvl__lsbufhv2lv_1_wrapped  rstb_level ../mag
timestamp 1608153117
transform -1 0 137896 0 -1 51956
box -66 -83 5058 5000
use simple_por  por ../mag
timestamp 1608153117
transform 1 0 654176 0 -1 112880
box 25 11 11344 8338
use mgmt_protect  mgmt_buffers ../mag
timestamp 1608153117
transform 1 0 212180 0 1 246848
box -1586 -1605 201502 19557
use gpio_control_block  gpio_control_bidir\[1\] ../mag
timestamp 1608153117
transform -1 0 708537 0 1 166200
box 0 0 33934 18344
use gpio_control_block  gpio_control_bidir\[0\]
timestamp 1608153117
transform -1 0 708537 0 1 121000
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[36\]
timestamp 1608153117
transform 1 0 8567 0 1 245800
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[37\]
timestamp 1608153117
transform 1 0 8567 0 1 202600
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[2\]
timestamp 1608153117
transform -1 0 708537 0 1 211200
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[3\]
timestamp 1608153117
transform -1 0 708537 0 1 256400
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[33\]
timestamp 1608153117
transform 1 0 8567 0 1 375400
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[34\]
timestamp 1608153117
transform 1 0 8567 0 1 332200
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[35\]
timestamp 1608153117
transform 1 0 8567 0 1 289000
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[4\]
timestamp 1608153117
transform -1 0 708537 0 1 301400
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[5\]
timestamp 1608153117
transform -1 0 708537 0 1 346400
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[7\]
timestamp 1608153117
transform -1 0 708537 0 1 479800
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[6\]
timestamp 1608153117
transform -1 0 708537 0 1 391600
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[32\]
timestamp 1608153117
transform 1 0 8567 0 1 418600
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[31\]
timestamp 1608153117
transform 1 0 8567 0 1 546200
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[30\]
timestamp 1608153117
transform 1 0 8567 0 1 589400
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[29\]
timestamp 1608153117
transform 1 0 8567 0 1 632600
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[9\]
timestamp 1608153117
transform -1 0 708537 0 1 568800
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[8\]
timestamp 1608153117
transform -1 0 708537 0 1 523800
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[10\]
timestamp 1608153117
transform -1 0 708537 0 1 614000
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[28\]
timestamp 1608153117
transform 1 0 8567 0 1 675800
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[27\]
timestamp 1608153117
transform 1 0 8567 0 1 719000
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[26\]
timestamp 1608153117
transform 1 0 8567 0 1 762200
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[13\]
timestamp 1608153117
transform -1 0 708537 0 1 749200
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[12\]
timestamp 1608153117
transform -1 0 708537 0 1 704200
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[11\]
timestamp 1608153117
transform -1 0 708537 0 1 659000
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[25\]
timestamp 1608153117
transform 1 0 8567 0 1 805400
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[24\]
timestamp 1608153117
transform 1 0 8567 0 1 931224
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[23\]
timestamp 1608153117
transform 0 1 97200 -1 0 1029747
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[22\]
timestamp 1608153117
transform 0 1 148600 -1 0 1029747
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[21\]
timestamp 1608153117
transform 0 1 200000 -1 0 1029747
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[20\]
timestamp 1608153117
transform 0 1 251400 -1 0 1029747
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[19\]
timestamp 1608153117
transform 0 1 303000 -1 0 1029747
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[18\]
timestamp 1608153117
transform 0 1 353400 -1 0 1029747
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[17\]
timestamp 1608153117
transform 0 1 420800 -1 0 1029747
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[16\]
timestamp 1608153117
transform 0 1 497800 -1 0 1029747
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[15\]
timestamp 1608153117
transform 0 1 549200 -1 0 1029747
box 0 0 33934 18344
use gpio_control_block  gpio_control_in\[14\]
timestamp 1608153117
transform -1 0 708537 0 1 927600
box 0 0 33934 18344
use user_project_wrapper  mprj ../mag
timestamp 1608153117
transform 1 0 65308 0 1 278716
box -960 -7504 592500 711440
use chip_io  padframe ../mag
timestamp 1608153117
transform 1 0 0 0 1 0
box 0 0 717600 1037600
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
